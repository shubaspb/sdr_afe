  (* BSCAN_SLAVE_INDEX = 0 *)output update_0,
  (* BSCAN_SLAVE_INDEX = 0 *)output capture_0,
  (* BSCAN_SLAVE_INDEX = 0 *)output reset_0,
  (* BSCAN_SLAVE_INDEX = 0 *)output runtest_0,
  (* BSCAN_SLAVE_INDEX = 0 *)output tms_0,
  (* BSCAN_SLAVE_INDEX = 0 *)output tck_0,
  (* BSCAN_SLAVE_INDEX = 0 *)output tdi_0,
  (* BSCAN_SLAVE_INDEX = 0 *)output sel_0,
  (* BSCAN_SLAVE_INDEX = 0 *)output shift_0,
  (* BSCAN_SLAVE_INDEX = 0 *)output drck_0,
  (* BSCAN_SLAVE_INDEX = 0 *)input tdo_0,
  (* BSCAN_SLAVE_INDEX = 1 *)output update_1,
  (* BSCAN_SLAVE_INDEX = 1 *)output capture_1,
  (* BSCAN_SLAVE_INDEX = 1 *)output reset_1,
  (* BSCAN_SLAVE_INDEX = 1 *)output runtest_1,
  (* BSCAN_SLAVE_INDEX = 1 *)output tms_1,
  (* BSCAN_SLAVE_INDEX = 1 *)output tck_1,
  (* BSCAN_SLAVE_INDEX = 1 *)output tdi_1,
  (* BSCAN_SLAVE_INDEX = 1 *)output sel_1,
  (* BSCAN_SLAVE_INDEX = 1 *)output shift_1,
  (* BSCAN_SLAVE_INDEX = 1 *)output drck_1,
  (* BSCAN_SLAVE_INDEX = 1 *)input tdo_1,
  (* BSCAN_SLAVE_INDEX = 2 *)output update_2,
  (* BSCAN_SLAVE_INDEX = 2 *)output capture_2,
  (* BSCAN_SLAVE_INDEX = 2 *)output reset_2,
  (* BSCAN_SLAVE_INDEX = 2 *)output runtest_2,
  (* BSCAN_SLAVE_INDEX = 2 *)output tms_2,
  (* BSCAN_SLAVE_INDEX = 2 *)output tck_2,
  (* BSCAN_SLAVE_INDEX = 2 *)output tdi_2,
  (* BSCAN_SLAVE_INDEX = 2 *)output sel_2,
  (* BSCAN_SLAVE_INDEX = 2 *)output shift_2,
  (* BSCAN_SLAVE_INDEX = 2 *)output drck_2,
  (* BSCAN_SLAVE_INDEX = 2 *)input tdo_2,
  (* BSCAN_SLAVE_INDEX = 3 *)output update_3,
  (* BSCAN_SLAVE_INDEX = 3 *)output capture_3,
  (* BSCAN_SLAVE_INDEX = 3 *)output reset_3,
  (* BSCAN_SLAVE_INDEX = 3 *)output runtest_3,
  (* BSCAN_SLAVE_INDEX = 3 *)output tms_3,
  (* BSCAN_SLAVE_INDEX = 3 *)output tck_3,
  (* BSCAN_SLAVE_INDEX = 3 *)output tdi_3,
  (* BSCAN_SLAVE_INDEX = 3 *)output sel_3,
  (* BSCAN_SLAVE_INDEX = 3 *)output shift_3,
  (* BSCAN_SLAVE_INDEX = 3 *)output drck_3,
  (* BSCAN_SLAVE_INDEX = 3 *)input tdo_3,
  (* BSCAN_SLAVE_INDEX = 4 *)output update_4,
  (* BSCAN_SLAVE_INDEX = 4 *)output capture_4,
  (* BSCAN_SLAVE_INDEX = 4 *)output reset_4,
  (* BSCAN_SLAVE_INDEX = 4 *)output runtest_4,
  (* BSCAN_SLAVE_INDEX = 4 *)output tms_4,
  (* BSCAN_SLAVE_INDEX = 4 *)output tck_4,
  (* BSCAN_SLAVE_INDEX = 4 *)output tdi_4,
  (* BSCAN_SLAVE_INDEX = 4 *)output sel_4,
  (* BSCAN_SLAVE_INDEX = 4 *)output shift_4,
  (* BSCAN_SLAVE_INDEX = 4 *)output drck_4,
  (* BSCAN_SLAVE_INDEX = 4 *)input tdo_4,
  (* BSCAN_SLAVE_INDEX = 5 *)output update_5,
  (* BSCAN_SLAVE_INDEX = 5 *)output capture_5,
  (* BSCAN_SLAVE_INDEX = 5 *)output reset_5,
  (* BSCAN_SLAVE_INDEX = 5 *)output runtest_5,
  (* BSCAN_SLAVE_INDEX = 5 *)output tms_5,
  (* BSCAN_SLAVE_INDEX = 5 *)output tck_5,
  (* BSCAN_SLAVE_INDEX = 5 *)output tdi_5,
  (* BSCAN_SLAVE_INDEX = 5 *)output sel_5,
  (* BSCAN_SLAVE_INDEX = 5 *)output shift_5,
  (* BSCAN_SLAVE_INDEX = 5 *)output drck_5,
  (* BSCAN_SLAVE_INDEX = 5 *)input tdo_5,
  (* BSCAN_SLAVE_INDEX = 6 *)output update_6,
  (* BSCAN_SLAVE_INDEX = 6 *)output capture_6,
  (* BSCAN_SLAVE_INDEX = 6 *)output reset_6,
  (* BSCAN_SLAVE_INDEX = 6 *)output runtest_6,
  (* BSCAN_SLAVE_INDEX = 6 *)output tms_6,
  (* BSCAN_SLAVE_INDEX = 6 *)output tck_6,
  (* BSCAN_SLAVE_INDEX = 6 *)output tdi_6,
  (* BSCAN_SLAVE_INDEX = 6 *)output sel_6,
  (* BSCAN_SLAVE_INDEX = 6 *)output shift_6,
  (* BSCAN_SLAVE_INDEX = 6 *)output drck_6,
  (* BSCAN_SLAVE_INDEX = 6 *)input tdo_6,
  (* BSCAN_SLAVE_INDEX = 7 *)output update_7,
  (* BSCAN_SLAVE_INDEX = 7 *)output capture_7,
  (* BSCAN_SLAVE_INDEX = 7 *)output reset_7,
  (* BSCAN_SLAVE_INDEX = 7 *)output runtest_7,
  (* BSCAN_SLAVE_INDEX = 7 *)output tms_7,
  (* BSCAN_SLAVE_INDEX = 7 *)output tck_7,
  (* BSCAN_SLAVE_INDEX = 7 *)output tdi_7,
  (* BSCAN_SLAVE_INDEX = 7 *)output sel_7,
  (* BSCAN_SLAVE_INDEX = 7 *)output shift_7,
  (* BSCAN_SLAVE_INDEX = 7 *)output drck_7,
  (* BSCAN_SLAVE_INDEX = 7 *)input tdo_7,
  (* BSCAN_SLAVE_INDEX = 8 *)output update_8,
  (* BSCAN_SLAVE_INDEX = 8 *)output capture_8,
  (* BSCAN_SLAVE_INDEX = 8 *)output reset_8,
  (* BSCAN_SLAVE_INDEX = 8 *)output runtest_8,
  (* BSCAN_SLAVE_INDEX = 8 *)output tms_8,
  (* BSCAN_SLAVE_INDEX = 8 *)output tck_8,
  (* BSCAN_SLAVE_INDEX = 8 *)output tdi_8,
  (* BSCAN_SLAVE_INDEX = 8 *)output sel_8,
  (* BSCAN_SLAVE_INDEX = 8 *)output shift_8,
  (* BSCAN_SLAVE_INDEX = 8 *)output drck_8,
  (* BSCAN_SLAVE_INDEX = 8 *)input tdo_8,
  (* BSCAN_SLAVE_INDEX = 9 *)output update_9,
  (* BSCAN_SLAVE_INDEX = 9 *)output capture_9,
  (* BSCAN_SLAVE_INDEX = 9 *)output reset_9,
  (* BSCAN_SLAVE_INDEX = 9 *)output runtest_9,
  (* BSCAN_SLAVE_INDEX = 9 *)output tms_9,
  (* BSCAN_SLAVE_INDEX = 9 *)output tck_9,
  (* BSCAN_SLAVE_INDEX = 9 *)output tdi_9,
  (* BSCAN_SLAVE_INDEX = 9 *)output sel_9,
  (* BSCAN_SLAVE_INDEX = 9 *)output shift_9,
  (* BSCAN_SLAVE_INDEX = 9 *)output drck_9,
  (* BSCAN_SLAVE_INDEX = 9 *)input tdo_9,
  (* BSCAN_SLAVE_INDEX = 10 *)output update_10,
  (* BSCAN_SLAVE_INDEX = 10 *)output capture_10,
  (* BSCAN_SLAVE_INDEX = 10 *)output reset_10,
  (* BSCAN_SLAVE_INDEX = 10 *)output runtest_10,
  (* BSCAN_SLAVE_INDEX = 10 *)output tms_10,
  (* BSCAN_SLAVE_INDEX = 10 *)output tck_10,
  (* BSCAN_SLAVE_INDEX = 10 *)output tdi_10,
  (* BSCAN_SLAVE_INDEX = 10 *)output sel_10,
  (* BSCAN_SLAVE_INDEX = 10 *)output shift_10,
  (* BSCAN_SLAVE_INDEX = 10 *)output drck_10,
  (* BSCAN_SLAVE_INDEX = 10 *)input tdo_10,
  (* BSCAN_SLAVE_INDEX = 11 *)output update_11,
  (* BSCAN_SLAVE_INDEX = 11 *)output capture_11,
  (* BSCAN_SLAVE_INDEX = 11 *)output reset_11,
  (* BSCAN_SLAVE_INDEX = 11 *)output runtest_11,
  (* BSCAN_SLAVE_INDEX = 11 *)output tms_11,
  (* BSCAN_SLAVE_INDEX = 11 *)output tck_11,
  (* BSCAN_SLAVE_INDEX = 11 *)output tdi_11,
  (* BSCAN_SLAVE_INDEX = 11 *)output sel_11,
  (* BSCAN_SLAVE_INDEX = 11 *)output shift_11,
  (* BSCAN_SLAVE_INDEX = 11 *)output drck_11,
  (* BSCAN_SLAVE_INDEX = 11 *)input tdo_11,
  (* BSCAN_SLAVE_INDEX = 12 *)output update_12,
  (* BSCAN_SLAVE_INDEX = 12 *)output capture_12,
  (* BSCAN_SLAVE_INDEX = 12 *)output reset_12,
  (* BSCAN_SLAVE_INDEX = 12 *)output runtest_12,
  (* BSCAN_SLAVE_INDEX = 12 *)output tms_12,
  (* BSCAN_SLAVE_INDEX = 12 *)output tck_12,
  (* BSCAN_SLAVE_INDEX = 12 *)output tdi_12,
  (* BSCAN_SLAVE_INDEX = 12 *)output sel_12,
  (* BSCAN_SLAVE_INDEX = 12 *)output shift_12,
  (* BSCAN_SLAVE_INDEX = 12 *)output drck_12,
  (* BSCAN_SLAVE_INDEX = 12 *)input tdo_12,
  (* BSCAN_SLAVE_INDEX = 13 *)output update_13,
  (* BSCAN_SLAVE_INDEX = 13 *)output capture_13,
  (* BSCAN_SLAVE_INDEX = 13 *)output reset_13,
  (* BSCAN_SLAVE_INDEX = 13 *)output runtest_13,
  (* BSCAN_SLAVE_INDEX = 13 *)output tms_13,
  (* BSCAN_SLAVE_INDEX = 13 *)output tck_13,
  (* BSCAN_SLAVE_INDEX = 13 *)output tdi_13,
  (* BSCAN_SLAVE_INDEX = 13 *)output sel_13,
  (* BSCAN_SLAVE_INDEX = 13 *)output shift_13,
  (* BSCAN_SLAVE_INDEX = 13 *)output drck_13,
  (* BSCAN_SLAVE_INDEX = 13 *)input tdo_13,
  (* BSCAN_SLAVE_INDEX = 14 *)output update_14,
  (* BSCAN_SLAVE_INDEX = 14 *)output capture_14,
  (* BSCAN_SLAVE_INDEX = 14 *)output reset_14,
  (* BSCAN_SLAVE_INDEX = 14 *)output runtest_14,
  (* BSCAN_SLAVE_INDEX = 14 *)output tms_14,
  (* BSCAN_SLAVE_INDEX = 14 *)output tck_14,
  (* BSCAN_SLAVE_INDEX = 14 *)output tdi_14,
  (* BSCAN_SLAVE_INDEX = 14 *)output sel_14,
  (* BSCAN_SLAVE_INDEX = 14 *)output shift_14,
  (* BSCAN_SLAVE_INDEX = 14 *)output drck_14,
  (* BSCAN_SLAVE_INDEX = 14 *)input tdo_14,
  (* BSCAN_SLAVE_INDEX = 15 *)output update_15,
  (* BSCAN_SLAVE_INDEX = 15 *)output capture_15,
  (* BSCAN_SLAVE_INDEX = 15 *)output reset_15,
  (* BSCAN_SLAVE_INDEX = 15 *)output runtest_15,
  (* BSCAN_SLAVE_INDEX = 15 *)output tms_15,
  (* BSCAN_SLAVE_INDEX = 15 *)output tck_15,
  (* BSCAN_SLAVE_INDEX = 15 *)output tdi_15,
  (* BSCAN_SLAVE_INDEX = 15 *)output sel_15,
  (* BSCAN_SLAVE_INDEX = 15 *)output shift_15,
  (* BSCAN_SLAVE_INDEX = 15 *)output drck_15,
  (* BSCAN_SLAVE_INDEX = 15 *)input tdo_15,
