  (* BSCAN_SLAVE_INDEX = 0 *)input [31:0] bscanid_0,
  (* BSCAN_SLAVE_INDEX = 1 *)input [31:0] bscanid_1,
  (* BSCAN_SLAVE_INDEX = 2 *)input [31:0] bscanid_2,
  (* BSCAN_SLAVE_INDEX = 3 *)input [31:0] bscanid_3,
  (* BSCAN_SLAVE_INDEX = 4 *)input [31:0] bscanid_4,
  (* BSCAN_SLAVE_INDEX = 5 *)input [31:0] bscanid_5,
  (* BSCAN_SLAVE_INDEX = 6 *)input [31:0] bscanid_6,
  (* BSCAN_SLAVE_INDEX = 7 *)input [31:0] bscanid_7,
  (* BSCAN_SLAVE_INDEX = 8 *)input [31:0] bscanid_8,
  (* BSCAN_SLAVE_INDEX = 9 *)input [31:0] bscanid_9,
  (* BSCAN_SLAVE_INDEX = 10 *)input [31:0] bscanid_10,
  (* BSCAN_SLAVE_INDEX = 11 *)input [31:0] bscanid_11,
  (* BSCAN_SLAVE_INDEX = 12 *)input [31:0] bscanid_12,
  (* BSCAN_SLAVE_INDEX = 13 *)input [31:0] bscanid_13,
  (* BSCAN_SLAVE_INDEX = 14 *)input [31:0] bscanid_14,
  (* BSCAN_SLAVE_INDEX = 15 *)input [31:0] bscanid_15,
