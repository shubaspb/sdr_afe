`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
W3QYENMyB4OIfVo0wlON0s7Z4KbziP2GAj5Jk6g2nY67XnPU9cq5R0Ru7hecNqzDzTsFlXb5U4Qj
qQMKNe8+uw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
AJpl9/ZLfl2K7X7Ffb3xvHvdWeWxH4YUxmX8RY0i4M6gGSwhBkH1mCxRIm1xcgWZdyzqDkt1cnpa
WwBxuBauHP9Rl+PsMOxLWL1pbK5Hl8ViwkdcONjZ+kXZ6xCXgXMgh/N9l6g4D2cxe6HhGjN++ZXz
wsrr904iaXupmBEnJoE=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
uOjmCY/kmmiuhkEdB0KlL1XvJlmtXEwCLrjeR0fmFXMMVlQ79b50qikIAGc9zm74RUPNqDMtfVDz
5/VBy1QEJFMQ82v10G0YeDjPo7tUA0gMy4IuY4KROdhEM4NJq6P8E76abW+NhXctVwxd4heMHXZF
k1Ne3eKXfrAPvluaaMOX7Ioku5FWJYaDeBvKt6JK9CcTK+CsO5UbAmGEEz/j8T0a2TMr5H+QHbNU
VSn3xDp0tLK63NmNMbDSMhHkytpYrFQztzvYtPGuxks1yqgOLTeI1j10bwcRhpnlHflbQ2ucp1iV
ONbgz9wOXXNFYLcsYzGzm5lrnSlE6Ka4ZmxSuA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lME5n30WjvWwWXzKRcQiy9NG+x2U59/EMqzhpBqDfGL5r+KFCSMvBxO/8hmSwhDD3+yz8gEdvZdR
Rl+gmiPo+Ps/p9NdcRm7mthzjnKnU3k3FdRQp+S2lhYHSeYzKQPl4HkPHcSBy99/a0shpw+syyPr
lVZsH17exhw+SZZS5Lkjod9Jo04D5B8Noh0SanKpkhGzSQ9sOY7CW2PODFoAJl/RchWmu+88xGrO
nmtE+DjC9776/jDJN6KlfWRb4Hyw45iwk8+Yuhp/xNDZNNauEW/eZM4psojITFA0BbNYNjXK3k0d
33NfAR+mIXalnQQbdtmKLKkO/TtSEduRIPUkkQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VVMXGhEfK6FFfvlcSwxIiFqJ9oQ2yHdR67AaGM/TEZK2Y2CYUMrhuZw2fOVG6SFlN1gjck2L60eY
glmcSVaaKSKc3n5fK7a32FFMKPj6RSiwfXaDCHQ3hiknyc2x2400dh6B9ZLQQMyiNYg1CM1ckBZ8
1JqneMnQC08ECmBMN7rdYPQy5KeVeHTPFmrlu8cCuoA2uYLVaW/UdokXozDxDJPvSukiezAjCxMP
cieoCVxD4WiCNnlNUCDCQn8hkuloTORYODgEgRdkVFgMVzk3MmEXao1Oo9Ku5qWw2+ZbKiwOAU/X
IrZaKB6I+UP3d4iZaX819FQlZ6FL7hNc38VAiQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GoGoxy/t9RLFZqe8/xU96F64dZCv79e2ce++JMkCgNPUR4SLCLaVzCxJQuUGAvOplw9S4oEFkDMU
BVxa6RmEBALqGa6BXOv+b9HCaDD8kV+4WG/P6OgKjYky8ydq/ng0xEWBliazG9uJe7DmcOLyUb/u
dFKAzcT01NrFtQVIA5o=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TLhvJbErY/BJqXkbfGxUtHlOl55qvwYmyZyGAPhu1DPk+URY+ZmnocQeS+6XeimpeJVlIiPg/aRE
8NNGcq/cmaXuYI87EH78V7FVe+LYvod0voL4SM+cE7Bc1F0FYhNm8eHS+S1hisSbwgDJVuGmvRCB
F6rkV+PCe0pkRdz5Xw2d12KvALMOkxjcmzqhP8rsa8P/XfrS/86JPUNm8Y761cweShPOi3Gz1VnC
B9cUgV0viAO1agJTVZnVAvfnBiYCywt3KqiQhSqBg4IMncGDuPxgEeC6nQ7lD4X2UiwCnogJlXZ3
IbW9lbWN3UPGIjkJ40WO4DFAUtb7fvRZz8ZpcA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1798864)
`protect data_block
F4wt8TTLfBO+bKCbOEigyBFnNyGVFFpuxKzYNvBudw0qo7vtC1hprOuR+3c1Njig8isZigvh/oJ4
nY8F78GSrtOyx20CMnXYxQMxLdKa/MGx93K7utn+dluZCP0u/BpzWUEVf9Xl5TMaxGi0aQwtITxE
sAdmdD00U8Il589hXxgIGbBVuhg6u3fIJzVBjtfIOsnrsJWiddY8+3ILteJ141JsnUtMd2G3KCpL
zD9MWuLYaMukqypgSuEr/hQIxAJ0yqFKf+LSptEbZce3mgPt3SvWlZCCeIv5LKwDCNSPNug9Dd0C
LtoaKD9e6zSADj6P5Q5N37wLE1aCMSbpT3cvoqkka5x0YYbutj/lF0vQYruFr5HfwalCGsPuQ5qu
5ElfghowFw/97KTHB+KFqP2+mkcqeUPB5pBXdYJVqwAkJ//c5zC5q8rZsUOTaPY9+Z6LU2XIWXXO
Xnosf25F4i0ZaIS85KYegdTSJseDJqztlqJD6fgMDUqpbVlEamIp2/TySNHTmWNNB9SLmlnKTA8a
/i137Y9bGpZKHN0dH5t6tIj8wRjFlnxyKIa+ER6RsHYCyfBLT0PyOA43pICOkEXbxJFjf+MgHhve
zSb6MK5uiVIBgdLag0SYBk173Lk4KfMTBVr8AmPEM/jBWDEGHL7TudKuAonjRqFXqTax40s4MYho
VK+4H8UtdzoQCu5EwCYNgKN4qjDRhG8lOtk+342RpP4zqeaOnrenRHlYvzpbweYo8UwxA7og7K9C
WlD+Mm4CRaAxvb0lZr9FO5oDXqTZv+CS+80GytLI4PSny//NG6Bq+KYOjvXHtWW8eJRT5ydYnsPZ
TSShKVnO1juVGKY2d+vx3THrG1PJzPleDDCrJavfIqzdyHVlz4zb3UEpeG0lHkBnJMlUz7RZEQNq
6Cn+yHRfFkTyBAsVGmKwKHq60qB2MkzAn0yqrSD5RHZRKF+Lj709uvHfo1+EMC9YpdsP1wuH/lWa
Iy9KfkoFssGLkw39+hiWKULSTjf1O06MHbMxlVody2Su0dGbALKy2+LRfNAs6cePUeprd0vfWI8t
jZFS8cxaU/sAWw3j2dRfp3PCweIC9C/IUJg+lPKbWnyv1lso0Vo1jRtwtZbOfMD29oAZioWZ/1vL
WYJvVnCvLBw0RZ6zzkl8NEGe7gxVoYoA1R0xuOvhNm6+ptKriU8e/vh44QPgVWWBH9OqqYkTaNoU
/7IrcKKb11Qp3k73OXRGIV9Id0MMW+B2PsoJAWqILTzkAHcPOA2S3CloxMfqnJYXwAGIs9q+y/0S
eF84YUU4v7PZan8u7Z1scmezwZYeZATw1Cy/sqAWMJ0XxyldokeoboiM8ZHAIJrLkKZ14kZ5oKuS
cyPl6PtXcqIKue6SndGN04rAlavEuec6SNNHyZARxSi+TmyeUh9QtnGTs4gK1DJwywc+gayTO6gX
SX+KiVpQqdPSyTw/XR461D6O/Gh5JHXNv4zBrpQz4DEDunsSf9TwYnpGMrQwmskHKYoCBXl2Cg9r
yKRD2W/4xB6/QXjSqrvWn1T88U6QmNylcJpfeeyFNPIBY9TZBEOCfrgHZCrWdtLD0RgUdQoj0qvK
r69cnmweVgq5zqC3bwwcGO1SpJBt+YQ4C0qjMG4RxmugmheeAothcNKv4aCfPA3rBkSCpHOjt2If
GxPx5549QS3FEZkuQwBkM29dXzqGJxU3zen+3uepfVI+ZTV6TfEtKnMNDwFbISj1QRERxz/eT3oa
ssK18L3Y99ILWi86HNP+0K9QGNurrJmv53DIIvjD5/degjnWMWdyYkd7a0CQ71zHRbWAeIqsdrMx
sptE/YfnJnG4ZUtKRIytwwzBi0SqMk+jIrM1gAKv4UESJPyQUUHDmUcDdJgoz7YjyFddrx1wZqOl
Q5zsoXM+7qVSH3FKxymr0ItBdT1FzjyuBlu8hKtbfQNsH9sCuUg6DvjB855nqH7pqiHCcHS+BL/c
G/O42HH4eLnhdcl0vZrXQPF/CnoQqwaSr5dPejA6jgP8wOCsP1tQ0SWXP6zIi7MAMmB4B2xsgfmL
RpH+x49WFiDAMoXgbHGkaR68zaOjoin0VbttFxQddkacSd4IVAqBo0Vr4FmSIv947SHAfgoJ8je2
lbKMjMKA85gvH98/1t1F7zkrDaAzcmtjIwmAFBl1vRgohVbRCZYW+iNTeqnSZ1BlLCTf7rgpGggg
jQv3tYNKtCJZy3uHe2Lg3mow1E5JkFgqgJPG1tWrU1dVXogeWDG28bCygycLa6i700QZQRdhV7AV
xvOsAId/oS47jE6RRe/+Q5LkyOOAm3BdNVx662pAF6XiJUQpj4dP7DBhZgqIFIi2bQKgtKRbD6qQ
Bp4xXC46MOO3+W618vZfC30tlxrFr4QfnmZOcjr/X/udsyyhV65GssEDQQb5satSKzvk3qA62uug
kff2tkMQ2cn0xqpyORX2ybbr3BIP7iXRkDtFshgl3u/r4FCNPOi492brqtm1P+YmlbqFnDivBNNR
P9L6WmroFoaUsMgbLSbmqyFLkblwpti9/WUyPBJM6OgCXTh8kuRBjFcfEdgRmHD2TAFWM4F9aW/n
nBnvgKuXGCTHdPnAfyw/uEA9ZvTnXEw44n58UM6LIfRw6Svz89TOz+ShuuoGsefjrVtlol/yFA6X
MCWqTZufiWOF2twkA1od+vL68XiPmnP3zbTDjliaUunGCCsE3usrRAn7tUqHJWVRkZ0Mzh6nTyUw
unhN9m0wAseyLdsnZlLoLSxDuh9hIP5xJdSMjLrKQgIA0G8h2mO5KooBGU0fp4fBzTAnIx32a1bk
4mRe9Sb0RrIyn7rLTJCrmoNtrm5Tm0JZAQTWvd0b9BwMcsldmWfpnidTDL4mVIG8zND2R1yVZ/yD
qSwve7tbTWreM9YzYqg6wlds11BtD3B7v9sqmPxdWky3itWW2P+f9OVzlv2RgSwkhy/Dlfw7E3M8
rQHxOi7H6KPhT+5BUgqhYfnxMX0PITY9eoKjAgvmzfMB/26FgWzflmnA54xeO1PkIbTEMMw/MlD6
jjIR6fC0N8Ph1e9dS3cHmwAYWa3+YrsG3nf6jOrI7Ao7l5us9sI3EfXTNJiw4Ld8b4IIdP/F5ya5
6MgZkxGldcp6o6Ey8QH02JUhn8p/n4Jg7tI8rDF2ERaPtFSC2LcLXBIFwg+6KVXwj+fOE802ksgb
iaXYJJ6x7IS42r6GJf9pMYYnJdC630VGpgqqomjAHHN63sBLWppVXorDY0EwLe5+Y2M0l+1bW5Go
IRC9rO7UNvw/gVRdNySAvRH5g1pkEfk5seUev8JbCyMNXd3Jw4wjC2p12f+4mLaCyGYLV6cO0w24
1cRE+nei4X76Fx0WxX2yJPGG25BdJ6suPddm/xsyf4Ok1nz1A8c9aioZqtxxSuD+iIrD3glIcUKw
zv6AehJQIZ39bt6noSxmpbKzY1dxGJlga8WGvJqt2VfXy9hFf0jSdV+2uR7NAZar1w6j/nuk9pGk
kfTmRquk2kfXHh5bPkafTJEpFTwbZe3wRcpUMqbMfeekzFerD4phrUULDVfuILlheDtoQsFsgYiL
b+BKIM8WqDU9eSKo9TfF84I5HeoO8E1Lb6d2Ol275cpW1lrD9k+lj7RgBPtUsY2qWLPVKLxhYZ8B
sBHYb/hhFzVB+WIpctctilYojw03F9tK6PRVeS96mK93u/M8905QhJ2LBbinrw6Uv6D45Zbra385
QpjND5M7DG7Lmn92xGT38aiAZusLEsVXIxvpknRNQf5179ECVD0zsDOnn7IZ/zosmDpK5PrgIQHj
xZoevVbOkG8XtQaG6Jb0wsV65GVB4/CisMDUqepwvxV571pZa86B/dBpjjPYuaan3YxJzqnkMMJC
EgIpjG1k4dvmgBe2fQhXiVEficM0eJQ1JYGuk5kowHUpXTenknHi38k8BEsB7roO8KwPhlWm601n
3qp8qKXV8KL+TCQT/JIjB5axg8HzdQrhtbvdaz8xd2531bIfiIJIht+8xOL+2SiG+R2tU5KY4ojb
XXD653JkS6juUMvY3lURz9mj1yLmAFXfF2lC3dRXlMzIBDMzjdgu15f09bSpBm5/cDXnIFMCk1el
kAzofBGs0ye99YO1DzuLHqPvpKAY+brlrOFPggkpV+7HoEFaQbGA5xjh0GQ6Vu34mGLOfVlT9Mkg
6zckL5VXWgNi1dgKS8MP1Gu+5+7p3w9qqgxPXWUceWCfdmt8nXoCwMVHCgDwvSXhhnNXLWACNBjD
JeKiSAFGGEUVT2PyBRkiCrNqm9UDKYd90vTN4yVnSDGn/VgiPVBw2y0kJT1yyUV6rEoGVzZTYRLZ
ZN19aJJCHOKSsRyFlUPH1e9qaeOqxUlOynSDPvgALCbS5gFLavfo/+v/7YGMW6SyZIa49pNJsvQP
JIZYGBrGNyGt8VhisSu8qmys5eaOcPOzX6S1grQ4UIsRgPhOCFY8myoRJ0s4FzFZJRkqRhBuDHLY
XNwvmyAOnEsYXAhcFa/Z1cNUkGknUyllNeapa5F+4Sy6Vz5lmwcdHzzxhTPRF1Tl2sMm2BLowM8B
4/zE5jgg2D/OWsNzDikd60kvijYN4cJPqEDmd12zjKP+ytG8cxPdb5JOcM+m3fHCC2Wx2Qj+odUP
lfwfQ3O5xc15LjaLG/j5d+lZYl3zxtj0lrraq62mhTyGifkD8Q7AMUlQ8V67vQDWjhV//8OcvnsW
RJAkAIbY/UBnyAbx1VXsULzztH7XXEXAEtYuhuPO146IWYZRj0OizGzQFSlrIiKp9NRQFaeiWwvx
ftzXi/SC3j6Jhdy2KsMmFsfnlALSlNE3rlnWt4PSOp+Cvb34yR+sitz3y6tXCvFKFMSuHwpMDVTy
Akjga2Iu/NrDGHkN+xGrovdic2sr0VZEMNSpKQY5b0YO4NjFEYBd7pKnu2+4P4jESLcRw3qIuBOR
uNG7VU1dM7CJdsKX0Tay9IN7U7XGkkZoTfqWDKAPhNDUrH+f6c12x+KRMWz1AT6Kk4m8aANxk9nf
Eood9LwGP9vdfydDOWZuRIpU3/UB2waPagio6Su8iNjys5SaZvoh1G7qJqdoLigCpO5AkKGh21pX
vXiVHbJ3/fYeGe3z6DlJpFqHZN6m+NKwrHcfrtG982Qgp9TLPDLm6UOiQJ2jahMGqLFNMqJtWP55
PYq3j0ZkMVXFcgm4yaaqwGXlTnhN9OqDiYB7aREtkFV8tSeDW9cP1/06L4eHHGfuvAfJ52sSI9Vw
4aJT2OkmE7dOQ3MaUH+AvwrwT+wFG0d7twFzca5oaKRGitbhrDnI7eAJZiswS7oZ8uiCyJy+ffgc
DzxCop3jTQFctuJwGDj6hs2Edg4orKQFWIp7PoKyqFcovFXMMxWQRTAueHfBeQnwFWusrS50nGt0
DqzWSZ5AsnYh3UddUArFl82uBAd5snBAQjLIR36f0g7wlrHyMomVGNVECldRxLp2mE0VPqrlJWDq
ytbLOZHZ/vgrv1GthgvtS531LAc7KT+4TSh/pKm3ggfzjHrVu9Y464qOyjdej7x+22XBpVGKAr7O
0tMqJOQY2tFXJme84i+XSloTB4zFwZ0NB5/4cPNU+5uf29KNdJVqpAJtNL7HcoZqAIg6iD2Mdrez
I4Hj6UH/AiMN3qp9w6TccnEtz7/kmVCqfwLnMJtGRHKjMYeL8OWDed1F8d/Rhoo3HJs7XCL6tBpn
jtZi8EHz4q8lLjEkuIqug6PO2GfK6haNt/FW4gxSti8EcxYhTSHGR0kjNCM513YnigXEkfVv6S6N
rxfJ55sgZXdok6zI86JWCac3typsuQtyfaOFhXqiPvj8zqKh1IZlbdiNuuCoLDfrTAMruhGcCdLX
nOG2yiqtHqGJ2K0Jk8iYAnlDh7t0CmMvrjfNs+VrXr60SkMU2msy00awIJuAfbrOICyRhD/SwBsY
N9tUZfPwlzWZ7Mg8x2f6NGNTjtxKsNnKHvHBXEyICe8No/iYXZTUMA36CA0wkIfuKuB4w8oEo6ik
6Wb56CB9KH4NZGRxOXP/H9CE18X+bUbIqA+OgcrWX4fFr9KafBJwk+gK7Ke2xaIYiv5Bc5dqLk3U
1oYXkENG2jW9IBqsTN35vQU7sRIqz1KH2jXDsWVUVBmNz2LGKe8QUFBDhfGr65dDoD7ueYRKhOZ0
/Dg4MKTVu6TXJR1IvN+tSJbC0sFpKGgOhy78Mi/dJo8vhIybFY6gdBW5a9AyoOURXK4Bxb3+J+6J
37h9z/vkF/4bVpu1sVAp0h1aTwDR+OWFrFPkK0wovUCxYqext63Tw8DSvvxjCDga19ByAz5+PDRE
Jp4vmvsrs7KJv3cRT6jIXCSOa8L2tC45khzo57vlYcLMhw2GqWPdDK9n/GdPnHPX7WwO+GCHnejP
ZcLM50UB1bDRlIvbEmfrbRUrPxYsNuEt1NHL5GJ1+T+WE78HLVz8vGqvsCOJ7Rvw9Yd0K9v3cjXC
gNeLv91LfofKNfBOfjoLEt0WndWTm9ATJClx3EQfxhkU7C/uqADQqhcjFEsPcHOjb+2JgFiBMmBJ
9qyjBZMCU3M26XZVwXyojX8eJ6/UST6sDO2dWgao1/Nz1fBDaTdFnbw8T4R5Q685/IcgeRiEaipG
rh8kpe1ZS2ThEOU0/pvvWmONRIpKOvqvsla4p083/PxNjb0pOn9iavcV3mpSyCaYcEso5RjHovO4
7TZUQavGSwAZeN9TIkZYgNSWg6B3KVx0sg8woTQ6RSaXI2KosvSFQzwGDf6Hn0FD5ec5nQW4+Au8
2XTUD3spzdLUhLh9KZtlKEunzPpkInw8ePwoRu03GmSs7ByxMUnK2HNNSXXAUt56307p2tR547zF
+b1YAFtZfSgiB/lOO5JgAzuOntQXLPg8X6TGk73Tfgu0gzGbjmAW7dkvLX7lp5OJFpvtyzXFLhSL
9i0QJNQDMHo5/JapeMX5Gdr03o/+u7ADPgtqEYNnj2QJAyF2HU9BRLsHOmd54bJmWw1cS6RaaZoT
1bNGIVF4mkXdqTeHi00j8aHOs2oGNdesujyrzhUVtwg2qUfPocrwm4+d5EKdI6NMOkpoWa11VDV9
bO5FUn49x6OMR87R/BMVYLxgKiasGMwcxtxDnwpGh1/IQwAdL5w3/1YNv8VTld54GjbGXBgyoOmY
gZOUmCluPBQ6AAXUs5M2aJH52zG0ub4f5P6phkM98cU872GiBJkLMYgdSj++/W0vCYeWCwihhcbY
Y/jI0eSl7YdCUATzRv/0OtYTPs/k2VRkiyExvPRdwrP/K9tFamY3wDQIyvIzr3SvUJGVDjaAZHVQ
mTBOuzX/8AuTcvppViDStZR+gtqV9uF8qG/qEpfEISl7Wxy/eAKYou59TIMv3/n8fSzmEkMnpjM+
MQOGfkgpqHO9FN5NKLlCajI3jhZDNPzCELOvtR8X4r5D894IlRKZxj3LXOqLwrVwe4e0OyZUhNho
QMKqLEl6ZFEcLwj5J9o1FaJAr8amTK5nE1ZP3X7nCuC+JvD5ph114guHcsilTbgfVVwbQMMLTFTs
BbfLXO5XvKN28mJl0mQYzJkAgNwHXrXWvsrR7VAALeIzJNa3lhv1Ft7RcWUzIl1MJZrF6D0EHjGC
PsIEJLgGqD7OP04Sha1XyAiQnf6Ac4uDHsVZEgb47lf/GTuqBEuesg2o3YNIekW7IPKwY/bfsUSl
P/fYXn7+tOqkKBnJForcyuKA86q5rOBBeaQ0YFoX5C1Gb+hMOcnrBkiTbT40LMXU47myVe3rnv2q
2ULyZEyDzbNzPodckKK+mjkdqEdZc2t+dsP90VUU6LWKpbmXE7D49s8uEvozvFVrQsU8bStRHi56
zHQVrnyBWKwvie+QcnmQvuf/thixNV1mLMLdqXNuET+0qByaIfT6AkzVFU1RdMQ/trEvObdwoYMZ
/9aP/9foOC+qTWV9hLNzPefjXV26Naesim7NR+N6ZIVk+fxFRH5q18KQpRP+9GCyafeUxyRJvn5r
lHZ74rU7FBB8scvCgWsBugTIvNlwW7fsOK94e7jcGgG5h7xvQuXnbmSycCrYq3jkeriUlyrZSmgY
FLMWppA1tFfY9P4zza4vyG+j54ZqyydS7B/fAPCfbydpNweoyNZzZJi3VXrt1Aq0AzfsdxIKPFM6
s8EAlCdtgRMb1GczSmwRTF8u8s3yOu1d/+TSqhI6kpTSvDFExe4LX7rEuJ2yujxnRM7GSQR0WQTT
tfqCu+gsrgdoCaF6dxzNXtxYnbuBKNtrVq7rbIPwQfO4L9d9DSCQrAlArucMUavCMxw1M7uv+GOX
ZTKYljRsKG+MmUiX28v0Vz1SolTEwykwsY4VMMSh2ebI8i8DdeplrM3e5XYbHOUckNmetZ6pNsD7
RLRFOe/Xl/WrAo2OJLruKaDsLWEEOOw5VyB4uez5HKcaJWMmLB+Nw3PU68iJMs20zwGspK+R8zv/
E4mYR+SU5QwB/94ej26/hBlg8aAFc+I020ihNx8Z3D5gGBr4JccGrFveEUuSPOtR4IW8qXH2vumu
W49YdLjOeETwa/A4H3vK+gBGsNSKH1RCYyuQ2DBh/ms/fJbTeo2UBpHXui3MaXgr61mbQps3yJPG
XfYX2yv1b/yI39sYOrf0yHk4yaJ0OBSpc487/BkGXlHaMFCJvHzGZEiyBGw801YtNJrSlCLzAFMh
hzyiLOazV1EFDnXP0+drexK1ltwZNDflv8rXIokc3D9xWe9wEih+lcyG4IykzrQ44CDX5xazzT6P
thW57tbJubRwBlGPQMEnC75IGaOcKmcF0OA9E8P3sCXpfsV+m5bo77WdQuAgSSnWZiscopOmwxJd
OUoO9EwxZIjWp6C54QIvXfAMfWMt88dLpLkdnvCYIE+QOKrmeIZtKco4vDXHYb5VLf7oHJiynDKw
BfBz1IvQCqsWjk3AQKgqVhgmhd6tzJsLp4eWiegjORsmBavIce0MGpn2V4kRBTZKUqULLu7h3kod
xu86ZEF3aV2q6+2t4RTIh7CqAArEjuSnDGaSPZJw9v59UawkEcfxQHQ+7DhG0pG7+N8Qixkw2bs5
EPYEvIKCHZ5s3bj4JYSyIiIF2m0IU2b0hg0dJr2TgVx5pTIG+XI0Ks+ChPwdtAoYwRv1g+J44InG
2nuXrMvf1dycQ4NyPDEUyWNWnODQvJtZLPqg1Ln4/gicVieDFs0FMRMHOn8/dQmuH/L6uemTYcV1
LZn6xuh7bawSyb16zZgLViR24tPeo15qRYM7733rrSIlq9bRIgVaYYF0Ypsuc6AYDZpR8R7wcyZg
fWGw7BMY6fILebfGsgw/dK7BdeYBOzplIcGFZIB9A+v4ljZQacD1A7DAop2bx1kYHchXiWsU+6pN
EvMef8u3aIWfS4Mit3fxPGKBWM6sCUW3O+zk1ZqdML7mlq1uhqY4oYU0YRknJPQoRfpA7UrYPS8X
Ouszris1qB1ImOxwMOXiui6+NBUfJz7hhTvILkDTwkhmA+POyYQhMj+2eG682jr2bSdCrdcRt/Z+
m+IRijKnkP/XMgkXeL+yfFjUO9j0o2GylM0NOhN9tniBLljtrNhCp7tyRCRalHvRq5xUgoAKgQcO
7alNsYlkLEx+Q1qyfuMzSD0PVrpOZ7iybZ96Zqv5oN5tSAlVHWFthZ3s78UPdml15YJnZaEV2kgT
uMYvQu6y9RpKAQnYXY/ZHPGp2mg38YAZpj1sxkx5vIsbDX7COQTmq1asSMWRsy1JY1pvVePFSdAY
Jj+bDNcjLXR46RgFy1+W8yyGm9ab7i4EoaS+A9xMlbFLMpjzVJiTxfI2MXka39+9QHsNSUcVMon5
IoXpOrlkczYvHNnnXGyDiZ/wowRme5rRFTmOQZgYPbaJ+rTkaBAQEhaKFOCTdsvZc29Nu/xOK2RW
YDbhLdiF8Z8iIjKqWOzN6FP2hClZ9DMjgjbKLuvFXeCqMpDG10Ge5cksaPDBwghTyRAmOHBr9Mgn
oSWPnHEZoQM7coSxrpVue45APnLG/G0dI3widIJVRGgX4P0uBfTBzT4TRDd454kEs0b2SXCLT5ZX
Re/YplYkRQUc+NQOWoCd02I0ijkkOqsI8T5gZFlbdDIbPGtvosnzaK+0uSGt2SsTbHcRHLLJ/7VL
5VBb2GSHRg4YasEZARn5nBpepw17TsryZvS8KEeUgEoVv7qbqkoLAs1qc4d2y4UPbhcuLz2ISFDR
XkeO1ONDM1uNvtt7E3KzCZYvaPo8H9wAuQliGuYbXaheF5hfaLDFMDqqcqZP+3iUdDz6zQYi9R2Q
ELJ4mh9Qu9fPkquRMlE+/iPXVJQdcYcKFdXY3C2dTzH1swZBgYVSI+kxi3TRPkGVuCacKttBApNy
Uz3ZlVz36a6F1wZ5YF4QihYKMOzDtljscxEVrkHl8CiJRBZkHRoTW7ojCfeJRON4OIpvX+jhSJdl
hyOdQHJeXmaneT/m6ND1dUBUap2uuWVKftOZVDhYWsgyELKhExdMPTqDvJysJitpZuPTejnJwEIv
H+GM3D6IAGwoN/178wMUgTUiQVU2Pm+dZuCvchuec4Ol92nYMjf9vzIPTKyfIn+hskM2nmlr7ePb
qxoyCeJWqEjzOxXt5rWF1jrRLsbenEaw2Sv1Igan2ZyugeosYGsgvZH6NBTt2gvXiqIHCaYs6ld4
XHZzTbSlscHMS/xbjZKcNdiEQW2OiG/C1vOACyn6vjp1E40z4ElY76dxv0CtwN8juLdX2QxGOS7o
jxS44kOkxWj+7QgxdgnzVkNgOsVaD5BiScJRHsJOXrpL5ycnxDh5QqybG8aat0hwlWGBaEZHkGMj
e4Y7n4owH6EZm8nZvZ8jyJkbt9qoYGF5IjxlvVvTn1DsdXG/RQzKYhd0THB9zAQ8BMJkbe6cCO6h
TTnDpccTPQtjBHf4b088/HeCyW+3ZiIK/A14XeEbkWnLT4nJcXc90jw5tF/Inm/ocgNiiPwIvFMz
7NhA34L3E7wSKTeQTnSRsTRfoED45WurJYdUT/+FJp5MO/MRhO2jBtTaK2H8d/BZGTFVO3dthQVa
MHeG8+xaKv1Xsiyglv8v9Ql80i9+aCWzSXtKVDcSco53KtU2KfCxJ+ykFlfmLk5UyTEatxnVMfs/
ZbHN+gJMjFet/cDd4GQDd5M5btkzOBsTdccuBAzqRJsEK5Hniz/pFcVQmNpv7aBsmCnIk5VlPDyu
djDGZiHOfmhaYgNmxb38flQjKgTxr82jbBzQ2b0vY+UNd7nfvi75iomB9W3btBhnrszbEt9RIhTE
hjVzrkGpU6Z8jhA+BLZXxS6aGmZx/4uGOMz0aEwARPbU7gjwjHv0hK76RzyCWYXdLIGbeFqZsyEq
UBBrwMXLqM73DTpbw8NVlDw5nP3xzAxh0d28F793PBYlBcHIOfF0kH4Vxgj3z/bEcqRRfFOBFlAQ
VokeyEigdKuPkpayN19Rwo/EoR0nZpA/gXYIFn1v8DGmpdXgLCbwN3NNvb7rcHpRmD50hn5DS1GF
TxmcM4gQUSVGZha6l95R2EQSO7geEQMErsxyo31/Zy0Yfs8GKodnNh5IA+pmrMZ+Sl/kaDTCugxU
5K8PVcaZnn1mLDIkc7hZyaF+ybdAKiYcnH/HUvPR0MtxzaBBV81x6JEoDAROeWzakoUkZCWv2HJu
9FdPD+J/IrvoGZc0LP9k+OLEsMpyI757SmgVzMzPvv9c3GbZff2epSlClFMk1iH1e0r1Az93mNAo
bsXxLghnmkkMLgCA+Y5mim08sQi9QU6853ulirKXDZQegftDACeJBu8RK+sCRhJC1fN8ZJfjhRgP
KXY0l0Pj4cuoq56N5l7AUlqTbEcr+UK7c3wMGzteN7/jqCzobCWh2LNI31g4krsYQPa1hyjDtOzz
O8QMe3ezL8jSoFgHboPuWYVokfEgsWXho8pIVReIonGZvrGy+3Q35PFC/LSaqDZ3qFdiaZ7YmcFm
+gCM3EC32jSo427ZIQQHWBE3rVlSIHEN0VaEF7dIyK1gKozpAaozf3+b3C915PzRAsfFs//KMTZH
hzFjT7Suh1hvYj7W6BTMpvBH/B4YHzmt8B7mN4L0Zr4mEFQ+zidwsGXHqAwi6v+1FTvVnqrzzn7t
ac3igah5tmjiz+I9B8ObuXs4q2dQp4F07crdra3Ckk4Ewvx1zbCOzsuC6nb6t6tT1RBOMBdnSTrV
hWxjE9YQqFeU0IRnoNt8ltJT+h3f+9U5RdMtmcAarQZKBeunO82S4MFb5y1+mSD3IgublN4HIG6Y
jlTX/7F2trfNPKfgVQgg5ZCW7GDlm/VmGkkiq/IDRlvt7v4ZdZHYcxgL0SDXbph7Vwz8wuJlR+DL
zUxPtlPAUWwl00gqyfekOHJLrJEb/2yPDk82dTvMdhrPczEG1B0qj8RAbyuqkYddOq9jhWU489KD
falvP4YyYhnzxO6YIUKY39g9LWKMJi+4gSGFI49BU5wiv6QFt+Dj03g+W1E7cJSK17b5RyyvO7n8
x7hnl7yrgYpBkqgA/vedtqLxqZm/xXa7msbMeuUwkz5ZwR13o4TZx9GORKhQq2FTdhFvG9CDmh03
VMYD1FAJBfwujMmzsQ/ebASXyB71aMeUYN/sSelQaqRsFJOpOcnR/8DhVoVKnRD3ENEiHW/YN0Dw
t6MfnrRUFKOKzqjCiCcpum2d2h1lzqvA5TY6NM/uUCj0hqvyzZtiUfzggsFVEvE6UbHeC+Ac7p7G
XdojwDuymW3zvbySNm+jTEKjl5cDnsQFWPT/xiVbZJXsT/JtMy4CdExanUKaf/nd1/Q8Iar9PZir
Tifk86QVYo0inxd7B5atam/5z55qiywIqNoC4YRMpcUdNLW9nHaCxIB6VZe8dHh8rbBWVrAbMC8X
xrmYMlBrXwnNoNr+VpVR+sWdvMl6LbjedLtZDkjLW30n9PC4h/TiVL5KQa1aMm884lj2dBrcPEJA
FhijR80/oDfMxT8RP+Aj/6PCTIXAm+9bP6FTGwuI+rt97AdSYKl36KTQfLmSWZZ9uKkTCOLwN+C0
jW352VM4t6XM16Ya6C9w7R72wSbcYEditcTl1fssHs68LczM/Rmew8kDSn7xruw/2vw2tHZOMpU8
BRyDPtVwZlhwlqBDda75aievYd4Ji0f66XjBpLAM7JUeX7vc1emvg4odNAgXyt9CK56ePdxfCiP9
ewndMYGaaB3cztTn6ikwiNGq8yLfDNGEkTVgpz1X6vame72hvNFYr5RSBA6UfrJ4QiLdTK1GrBYH
fnInMNDax3SSNaVfyTqHD7nqBxeGnpN2i6iw0IsY0Z6T+qvZ4vME/YsbgRmpWs2ppxZwt3+Hqnpw
GsIMNXlUS4lSItwTzMM66oW0d7ODUQuFGKzA3QprzEisOn8gL5fL+5yHpiCRl49Mp9oLX73GTJNw
7EatZ70rt+M1dSozF5I5u3SMAYQZJW7N35BoZvaIB+xughqhvC339vVuQlr6b29QBwfLfTD+a3sb
TNYs0mZY/lj0PyjQ0jIjLCiy0wXIQjgnRoVlNRUvxYPDv/M6Qt6/KXtdO76ook1kRK3p9GHFAutJ
ki69YIBQaVoUq1wAyn1nUAxqumb9M0zEW+XEYcrVgY66RKCkm9gq6Z1yMJKdNUlSPiCxsvTtUM1Z
wntfDrrPV6xQLXMWo75xKgUIK4BnhaRjQemSNCadV0FycerdT8vUojnHUZn+6M0KJhZT/NoQQenr
AAbJmwvB8YRwNFAUXB8m820s688kuBZQ01p/a/GQuFY6071kJHNrLcvnD7Y+mb9G8fC+Yc+PzBfg
4QLnxs4xfkxvxfBlVDyjWpz2Eb/WnDI8SNa0z4NKOV+0PHoPIKhe3DZ2YkJOwLnfe/3k1nHUk/I2
Bxz200UAgALRdV/xhtZzVRdV2RXRwEcAUgP6huWWZtwiPK4kvdNoIoq3MDib78YryEnNjwGN1mFU
X5ctmHVeWXYmrB7OR9PEXezC9iwF+QLUMaiZJqw/qQ/9hy+MPVjXWhDgrSIKHNC1yO+Zq74VYX4V
QXw578sCIgOdv+wBOCh0lRXr9fr0qw9+RvmYWNuKIbttx4P1PEoZ6pyyiNJClnCZZ/hZy7GRr6sa
qBCZJpkEsWT8B/qmdT2fJvbGV7/gq8dYUK/Psmb49YJsQYf4qk+0z1WmiePVK/nABljfvIriltVm
aaz+PiWlulVpJKQneKQqwAwGPK5N5Ig6mNA+TD9+SoIywIIh7DFlwJJzIE9ndBgs9V47lUTkbZ/D
0lj5zO7yU3buTVzu29mllfmT4GeqWn8hiffRu9BO5Ifqbgmjshty0AHgiCSVR3qZCiiO/u5TOliy
u+rop9+l9dGhpC6G+KZCQjIUCl9/eUHhCDVd0ZMiRUCLn/Y4NFzjFgxilfW/QnL2/zGUq/+E41aC
6XXrsuanDwQx32ypxbEvY2YML4B7jIapjC85kw9ChiU8f1vbMPZL9gmhjiWEcy89+aAYnTOxrgjN
hXYFPtgdF6PsZGkKUoaxwz6p6QLAAGE68VAu86/q/XeV9oVN43VYNecUdzaKRyPxPzALoX531CnP
+B/UB2o4ByHZaS2HJwSU+ZiFWrD59xILfTbpHCJj6bxHrnh0gYZtf6Wg78m0OkOh+mFFPbR6lBut
9fgEknzlKalFqSvioM+wueSfXeYiG8dXCZlNnigdpARRUzYSLA0BVCZJcwWXDPhoPaXEW/Ai7akI
WiPDwD9X4/FJ/YmrMS++f6y3+P2tknOnhQ4MbwDQacP3pGVjtPVcQulHyWzp0rym/UYAkctZjvAT
QJGhmvCvyj12+OhAkXCk48n1sUEu8c7go3sOcM51sMc1W5kt+1M5Q18VNoGykJLkmJYdWe3numOQ
xsl2MT0igH8oXZj2qSwFQyeDtbPM97QXBf3LTSGYBCG0c9yLJ7VIxV6daZKoCK+wmJ+uMOWeXvqO
I2FL+xOJlfzBFBlKhxGBgADxBBRrvRgh+wp5NOHpGAX2cUCdBs+Pd9hdxrRyGOJOXbNtzTDfGqgD
/LL9hu+03HhbEbJPmmQX8P3Au8rFKg4MMgeGIsoOwooyljO2zC23oSNIj7LKsy0l5ss/qydo/KBf
4AdxUvrHzw1IvV8Ho4hv/0F9o8IzYoHWzDEXoms50Jj4nun1ziHUERb6UJZeQPo4spL6R7i/m0VA
e0sQkH1NrzTQkvxsTzU1xYN2x9S9G4sBRZY1Ei5zFPBTk7iHoQs5XZ/zfLsQkZ3xvTaFuB8Iv6XI
YkikSv4d0qhkQwzxdD5oshtnsFgRxAmZo7tgGAL4S6n0AjFNjzzpaN4y5JmpLKJ5Ex4D2ehFkWuW
B+ZRCn60KHPQgq4Ui32ixEGfTF3ZR0BNX9H2qLjz73D17RFavlk6TcgUrVuFANeHF7LF+YK8cg56
JhD0E3X+o+BspS+BlnUuUzRy5O1pSrBH8A5LeEgzKMIJX4R47JjHgx1o2YgP2/e/RE9P3QCsWED1
Cn0Nvc22y2em/5EbWCF+JVi6LFslLk74V4gNy7zbA6VTLPAqXYvuTl2YH8jRp1iKDxOpUtxDLkTC
UoJf3eA9iuoxN4rqwiv41cBfWlPm6XsYb0lI7/l6Id+HjsgGWbnS7DTpxowl/42xNCRB0AR6Cpc4
xvHFtmzODC7OjpM2XLfK+r2us3jfaXczVwoa0l6IekUWsl6TWR0KpKgITNFIr/mm5oEkdEK4Yywq
xcUP8qPHZoBACx2gcaRKM8mE//wuhdnBuRHLEGHC2KBgClRpnvcQX8j0gH6pWZsYbBBXgEyx9whs
E7cdIC3nQzlUNZUd26t8hmnlSjRt7QFf4AMggiCFFylvbwczM3HonrnMjaLRJYXLJ15G38BGOVbi
LitiDM56k9tHxTGyQQdQLhyt6PEaUS3B85EbKxCgD+PMRhtzphJk05ZQJEPbohV62AGuGkZoI9Oh
8/PgTFmx5/0xhhg3VqXLhZphSBSr6qJItdT8Re9QT4p6KzL01W4lfOzf9w85q/iPcSZHyD1Yp4Nw
qwdH5dEqjD8Hmwd3nrlOk0a2uomvItRFCYagNh+7laP30VpBnr8htX0zX1T3bL2x1htZuutfL+C/
o0TeYEc09jDvXZgUj2dNdQ79ar005m+UPl9374HjnH48Sf7wAOKVtdcYODbvrWYW1QBi/e2Cbzbu
CbPcrMgGZlS2MV63AjDfDX1hcHJE5ZaBfqaJ/48cfWc7s4OzZu7vmQcC87SXWzliyTmQLV2Qu64n
g0Zcu53MUi+rr91oAt5k6Z25tVQdeSREaG3bfE8VCTYdcfhN8VTaKlEiOzylmtYAI/fPfgwRKlcM
tI1u0iGVSagGGhTbAJ3LucFYF1vmA2jN9y4zAKa5eWXSgu82XXQNOy+bZpbq/7mXeoTcZDrN+rTY
IIrPhc54jBn0eXw6a3Y07YQ3eVZomU6ROMMw9TgvbgrCthhIpxZVEVi+fHWsWLb/BPFsZ0MYekbl
A1xTg9p3zrNwkyfcgAnGozjG0Bq/+fKwXHVCTyAWl4rhACO1lujpj3Nv0DabrddeQ5vxlp5Mevlr
KCW0yd3+Pbgs90t0HOGgr5ntNajfmcpPzjCUeBjZ0H1f0Xx+EDRVyndbP+1Bo0sQH92NdU060wTd
vSX28Vv58+5DoOaZ0axqeFrfvzAxBEXHr5+t1b1R3V9VrteIuZ6qZMertfoLgch6hAne9q1yA+rU
8cGqnTi4XybIMaySujpzCGcPmeK0sK3S6ZWMI9QlZ+UDHOCu2nyvzZ1HpjCfGV4ziXYrMjHahnxK
MKl1iFKfvcKa9DhYIcUxXvC8J8jKkToKKI4CSPfESb/l1DM2nBvxpTIPWxcIoU4dvcfF4Iv2pRYG
rHaWB497APfkLN2615J0LSKmUGaY9QHurcQn1FP4i/dyNgbP4aL+kIYhNlJcDAQqM8u4ewTxfrrd
fjJor/dOhGZ/tZn1mYNl/knfXBmkm8HL5dNJh0nH6nIrwB9YY1xOrPy4YaVfn1XMwTc4o8yDyVMt
mg4nXxmI/p8pA2ATmk65E8FLE/5lyR/36xlrkh1ZV+RApU1PNLQBmZ4lZrrTFjY3Mw69nUADXCoV
7kpiVE7PH+/uq66hWqDS3G9IAshMBL7yoYB8yP3uSJVEsD1nusAL6PCN1cFJCs0Xr0NTVy3P6HuM
oS2eg1OExbeN7p8PxNeOglpAnvfJ1AJLClndm0TOWLR9uId1XzlinsLUkyINyAw1y9asLoT0172T
1olGYqHY92H4lKh0iLEzlnr941SJWdNjO2boAQlkafszhm4BHePLRVT6FcZwAhMdc1iMOvRs67M9
u4NEABFDVgyGdqhItwoHMWnFZD1OR4H8G1wwe8Dg2TPRtJFooPCqmKY9+teScwxJ2TiteYSyugmr
c2IXtAIIbucN4tK1ZCHdHPQ/YEuERgWFQTA1/IgxLCspnmHTXN64zNkNcuy4dGdqMa4aQIxCrj2l
BZCZgxT384Ig3mLleycppNFG6AkE0pJNejhtp3UM2B6nk4YUtZSAgq2Ep3zX+9g6bjSDyFzcgB15
zthR0zBLwePdOzlMEIDsH/Wk3qCUJCD3GUqh9t9PzQ5dmpQkOf7D9tu7CDZ8gxHeXlepnTFcmdYe
sjubZdvOSsvx3Tv3R7/5uORldhimcFeAZ6WA8snuP1G2HaAae/FAi4Jrf6CLJdljcj5h3pSEi+xZ
NpKbuyr1uOUHpXTYuhECw/SUfrpd4AbU36gVObFzYzVNRiWSnnJpVAnszGMNerNbUR3Lxd3nb32X
J8RsqSFs9WbZ1L3ULQkXyEXo/jjd9jTLczEfcOagugyu8ecdvCXrVE1vXV2ilULIWunXqgTLNk/C
NYLdsB6R6KUkBp6hiY5iob4ah+mbp2F1o+vA7i45rtm/pTr78dWfLScmebu4Zaa5e7YQOl8cFCOj
PBzo6nJybOeTxhZryhXM2OnC8dHJ/rPQjftLUvrF67Gst+OU56A0I9hSVW8QDqJM1V3I+iMIEgUm
e58kwM2IN3YdMXwnmrU2PC1gEZ0pQZLeKj6VLoOhq9BPA0/xHy410R7Cq971/yd3+kPB2nZlowHQ
VKRf02qzrPUInWEPrPGJ4gIRTzfW7omLBGwx1YPfgv5540k5kRxqlGEXy6/KhnSy0KA0y+LvIIXX
ucHWje+eyojcCQQTuO7Uzx0Z76rNeLU500CNM8SVv+ZShQQRvQpfLFwqJYwYeoCDBh8Z3Cq2Umcr
Edb7DqvSgV6T6awsodx/MQX5H1Wvv/wYkOinriutGm915zB/ahX4ZaWhLA/BJqouVDY2LmjcQa0+
5YvD/HvnWmvYmU3VxNDYkK676fbEqA44UP8Btlfd673s5oY04jalIVCZvScUcP7ffRAf3FbYS0zj
o/IsXphAxp2bwTSRHiMLrXMv7Plice0wtZy7JcPIbZooV462//iVnnnQC/AadXHsM/MQ5lVaGgtq
u9dIUhInJ3/pyJLbHy1DWImqoR6xoXlg4uK8JK/NMsSZsl78vdgdvxlN7K+XE+a0VHbwnPB69QnU
BNr+Zt6OF+EHBTakZV82Qz5kF9sf80pLeylollKmaLdr9VDsorVpmkAxAKamvEAFIeurFLLfg3pM
D6MBFRyFCTJGPkp5zqnm7HxXXqIt0Zle467xzCMcx2G1mdGnqyR+ttFW9fgsjmX0jYjDaKnwYWHC
mAkIvGdu2GSrf9LjA+EbWw+HIenRVhaXsPOWXMB/UofDE3G74NT1B5U1oglDRfuxmaAKcAZff3HC
jWQUr27LMwZ+CyP+2Cn/ColVN0CtzaD5Sjf/Vv1OnKNY3ouYG8xflpE9uzEBPvETu81vjbIDgAue
G2DxkaBiL7iCKfD58UFTkgJM5eT0vxCyqwhdvo6QGDbEzao3aq24cVPCujZU0oyhiEmCmMp7Q7FO
RBgfZuxlI/k5zavW8w7Gf9CQvdAIn7ld4wmBTj445pN3eVWCugd8LlzDUcMTrDIofluMYhwlmEPa
Vs04OIEl7fV+unPDyKRnb2KJnZBgyrfVox4dK7lHB3dwNwNvmvF/XO7tK4fBCYCIwE3gCt03CqzH
q6frxUZ58u8lvWZpC9lwuftU42BBe3D8BU+c8e+kYprpAbWcSZAosZB54AlDmRo7imp01L8hL/Te
l7v0YDKZUBNFCdMYftodrrp1MTsyboDqKIZ7P2Il2+XVRz0XxEvBWsnpV70EgFbI+6HQxUeIK9Eb
rN4wln1db9p7sgK6Gxwqai8ubhmQUgjoaZbPuObeqyKclfK4iQzO+hAwfaLLLUI+AjMZpfbag+tV
ujHNg2/FhcRmZtVV9+ohQXoP+ohTfIcsE4ghNGV8xuFOtsATPEwLrblDGMEYuwf45FoM8GhxzR2D
Eg+OwfAhFhGaUpz4TEwzB3N6G6X9hHb8+Qg+7PBrek8qtBee8FiqWTX5RQwLEuDAUsFB3+Cdnn7+
XKGv+Cp+ITeY8ma7MEPcCiIYBpLoFhMsU8VXh9aHxxYV89CD/h6R4xAmMcOUxTY2jwSSar0KXE4o
qGv6bzv23Iqp96940KJXBkb5P2DYnR2Sr/oSXU847CXOoBfCntFDOGFz5OWBqw4kH7uNKFr0ffDK
oY+EazyTyyR5Vatqv3v+ONt3QUsC7PK5a5hpgATq9WQK0pQ80aHhDNJ37yWzjlrLxtRZ3VVzJ1Zi
yBM2OqAvPn0TtQL7yKRPhb6RC71pSOEz6D+71x5mryElO0mQzWgjm+JvExcw9nHr1iiRKkiC8992
Pv6skWXwupq7qJ/8Lk0ay7F1a0/qZAerajGfo1zSvGG71BtX5+fvbHDH2fsc9ydY1tcHySyLfAGW
EfgcemlPIl9L4BsBChYrbZmeRppfSDSIiOOmDtS4AafMPcBPzMVTUC2Vyf6jEfR2dQppbaeh8VCb
hP1SkkEj4LuOlXO351YQu3Ys7ZTKdFgwcQefF2t4WE2Y7A3JXBtqI3nzhqqZOmPJsNl7sYUaND3P
W7Pxty40R1sZ5QRdMKqBELnMb8evLEn8QvhIutJkv9bSyzQgVmEcGz06Y/LnqP2hFFt3AqEOlSzz
lcFHRTG90RDHdqazaIQ4QXjXBLKDROPedvPrfJee2W+gt5ms1rIoC/+tDu6djwBJtGZvqkFY05Fb
/JtQBEUC1nW/SwBtKwV6pkhRHntdn5L73+X+6XF5BVbrBju9HxeAJXG/XefOx/XljuW7M/TTbT72
Z1lkgx/rFwwffi79IESntkcnTaiOMgHPhd4AFJojBxwKJoCCCTMdnMv7tZpW2LXwyYFBaHr520yq
0mydrc9Tmn8stSfKtDZjxQA4QEDulpQUFkyWhddgQJsDwaJ6wQsEvvNtsSaR56+fw5rmIsqud/S3
YSI39QRuU5GPKzXr9z3Kzh1LVDhIpiSM93IIf2zvrBzW02ba/92UYBwOz8NryzRq24498a4O65fm
AC0joC8rImx1YNIT/naeVDEsq57yUGj/cYRwmeePPBZhhEbOUEJPHchs59GhIxsDVGs4BaAqbUnH
cOKAl8FDIHiIq7nYlZ59FAtfVVpEI2z2Rgc874YzWww577fA7Il5fmILeokYDjsBiU90jQLOfnZJ
zXA/SPsQIllrpQLipxBtF/O0nZUQTIGsnfKvpsKJ86536AmivPHMGJXRkiexpTC+zeK/rPXZxgtA
vkAM3LzBdtl19SQQ/CuYF2TOpFcg2BdRecCYhA+LtZn/g92P90nmAbUM15qoCVREnSxZeWU26IEn
CcOjjNHSNIrBz9LLOAaPJfXXylHeuLnCny4kB01ePkuTzVnw5ICaT6Dzy9hqKcNdyvuKhVNI8R/o
ILoeck8qirtRsdx2cKwhQ8m4cLllzARykeNWEnlcG5ErKDy3utupEUsc+u8IzoaqhRxIz95DLFbZ
ISD/Lj9GtzZ6yAhNU2L+CKuKbs2TrltzXt4x16vsCr3cazXFAHXFWuSTXVVXqKxeLpJKw0OtNyI5
qz/ktoqcgZMINcBwD/F3+2+IQgd/KijoYCKk5S9ZLCG2v2vjL3pFL73SfptsEVMYiREkPjXWJwN6
Tp9dQM/7O5K7U0I1Idi95sgmbkJu/0LNt0sLstKJs5iKUduPlyx0olMPdksDxN2yBtMQKU6jsIWx
r2u3XIManua6VJut6zM21GTfJv2PkEnftP7SX0DuHNHKIU41jUZLwHeRbt1LVgQ84KQdDtn3yH6u
nYa9GarYvFV+Qu0wkN8ru5n0C31jYU2SDT31t6U06uh6jMMDmPY6VomTuidO+Bt2tP41IP0xwSAs
2C0Weiysil9cLEUDZrJd/X2Q95c3blJ2QWhF07nbqgio04UxdIEyfmw33o3hTO2YjJais8X7jUR9
813xGsVb9SI2/7B9rvIWBm9XBG/bCmDSsOGNI31s/RSH80oporLaKC9fhmFY3bS9cjdIj6zLcqhB
C0hzjRrmnlbnhb8KAyCYDwoxcaBO4EfuFil6O1RuPM9YGH5ojOFkHq4iJQ7146PYNnq/aIgNaStD
F08dF3B02ivtmEazQ+86ZPfmJl5oGYIAjziOEf+xC6Bu8HJdmbiFZL18vWyINukrOcMfWCz4r0EN
Ttnm5K8yjRZGZlGTbRULAKMVJb3J+yfOYbiZ5k+/JOVOv+ZLhDpId8c/H2oWwrABcljk6LYcz+Sh
H3bnHeSTgOAWvSpSN99vZ62ftmfCg+6NrXzfc2ibktXIZ+RKvt+9DVGdpyV5ycRYOIZYPaHbhpUA
eKQYf5vIMe8GXssE/nUgrfLqJSL8aNR59nAX8WqEL3WmaIWWKQfAIBlz2Dxl4E2dcB8eLq1hxZxS
53leE0wdefYI7tIYtgC2N3pp1E8tMacr6iXJPpX32Yf2gyOnVnDQsBHFpDWYUFdIGaaF1JRId+hF
9Y19NhZ5vE4FUNXjfX5fSC+SZorzdBJ19xYkCNP6YVQdtyxVXtHsgEg3KZ6DjFqAJ0Et8WPzu1ry
V+sqKQ2SBmrMk/v/ySeAqd4ZpT5Og70sf8yY3Yw1e6NqJck3O0tCKs3wMEyd/bOT+ULP51kd8I+n
iGHjGGsKXanB1eHfWXpI12RcmxmA4wVXD8exk2tRnbvW2hPMUAj8lX5g6CykQpsBH9iRugMaTObN
ZjfzJG1msOK1WnysZKSPFgsmFddFeQX0g/yBUpx407G30aDbSKHCP0ZPpAN2qlvAoC5tgcLftyPm
zwmFjPIt3ig1MsWPdKbOck/AEmTEx0+GK5R1GekF+sNexQl5q05MDxezzx6hRSGAscMNKnyLaSus
Gdk3EqQh61G58A9zobb0AGjlmHzrjlV/i08/6nLzGRatpm+PmvwIbhl7KGLj+CWLsJUwVV0PE2Ad
WnntSGpVmltvCFMvV1hBXv0aK7s4o4IyABHbzJYX4quf9lnsLeKPGYwzVht12Sy1FhxVKoRcjhV6
IJuOj0K5gkhtho2bCLNsu8uRvhmjsWAI08AWg4/FuGcpw8b05o8OhnYmlRDrmLSfFl4pcG42YKQi
/LpJBI7wRaZXj/QFKlhgPth8yKnAcAcgCwUqH2TR0sA6cz/FLE3k1gA1o1DAROI/eT4fMkKtp03p
6cjB4LlQ/zIAqqzDrqs9BjH0Z93TphmeBq0drZmvvvGuoZl0Wyki8UVLmxasOM+weSpWNHGtveK+
GOF0WlT+phPeWm9E2Y2nlk47bM1HAO3CW+K3QQWaQ3590BISf8pzWNwqYIWMoB1V2cYCTbYLFFeB
Jn1cE5bBHKNT/LYIQVwvFFfT8TO/WEYkV3aIkxe7p85BKQDi3YiULZ5aussSBFxyas1p4lAyrbNq
sK+RzQAqWzHhOY0GyxTtOYlCoqdjeT5QESZGFgklWUo1hpAGTu4CSSVU+JLHYAHnOrB6Ca27lbzh
GHK9vaBELXpnKYmL4b5XA97XYjBl+Heis6nEazGwjkwMyEFMge6HyoGx+z0RhPd9yHXgkZEYnfk5
HwOdhLjlX3s2Ut84zkpyGI168hc/oqUCC/DU2w9lCLm+8h4g2gbiwWy3amB4rhp8vmiwePAUBdXh
af7FGxicQGtW1rVwcZTCaJO6w3HRBtgV8ILpNF1FESOdmHSxIHmhGi5UqOSPwZ4l/gFB0Ev/uwkH
XBopPM2brNve8vwloSO1G65V0cMb23lK+ngTVuzz9Rz5iPZyFJl2GIIoimCGTcjWcmDc6wHWIdSr
iB7pB48DeX4R8eFk5j3XA7X5UE1nb/UNEuGoa3552TGQYYjWF25LDm1/NGzcZemveVqfHGyhCPO5
WKTbJ68RXVLcZL3CtxfNQCdNvr5UV63XgTyljvcbufmgnrSORDzN0rWGEc90ifCeYmsOB7xPuzgo
00A8eoab/XCrp3/Kxb+M6zHT70MUxmqGpbJ9KUmBNUj6gKUPfFzVz50hu07a0S7C6bP7qumtV+Vq
QRWTPJR0/+00oKvTk9PfL+ZSrFzNdN53v8u1xD5CEzrGLo66H3e4IA1rY2pYzK9ooO3q7ixFhDRX
eukPiwEowMhiaD5/zXo5aUCCGJsNjq+41LNXa0Ya5aab7N7KvhVbkfEMbXHvTZ/QpjgpUexYWgPS
DNe1Tsp9XP+safGPI6MGnv5Pkk+C7tao8sQKbDTwn9MW3WR0+zliF7ZLlrj4SAc23hKY0/c9r3Z8
V4jSXfeZXIfmTTDurdtGRLPvcHGIpPhV3kfS7Nb36NQjMViuv77IWe9hyh8l7yJ+K21RfwVJKldF
TtuvSnL7AatBy3u0B8ydT6tv3Nj1A4jEPujd/VLGsY2GxdR7M+gHr59bDLF55jmB42XbhUbO2H3V
KGbHYtgPfPlABuyBwU/7EsKir3Ou76vmM600g4dgP/Xk/q49DpR3WhB11vDIxYX9TKk84VdeWCnW
1dBMe1WiXlrazUJloZpCXxibwlm4E7aeJR3/AGWPMYB0I4vPi7FaInM3LCCmMETd1aTXzyx1V8+1
Hmu7e1QKj2hGnCm/fxH7GqLJYiYEMXcKGUMiN8egA+jSOK+hpLU9lrhoeKq9npn15Ror4YoZN2kR
//Lb0Q+uSCtWF06CLrKYUhu+f7IWNIZqZEkBePRsQMw4EP+4VbSNqCpgX4lnuN1DtZCO6U511dVG
a45ySVZOiVFTmABKPu62qVmG2FTigCBOvIcGedtky+owlQj7QylZn+0Qaf6FOjRGWT/DWVuHvWu/
iaxUdjuYC/nXwRqKRnS04oip39VhbhJl9Jhqy2wPylrzL4asTGv/LDU/C2eIDX6KWqRs/T01iHZy
O+7LL5KXhTCPbe/BdUFggBo5Nnd/alkvhxjsq5evnAs/vrksvWlGmt76576v5kxRKqZF4u5ZikWT
xIFXuoNF7Rz+BfUtuKQoEWtUwwMdw7Zl0m3mAuWKTYtiRp+B3tRmqMNm0gLD8pbMpozRxdQZpd1B
3VpkK6sfWlJNOq2ArpG6cgVcFR3K0tF5LunP6z6v5cjDE3HfkGP4RDlXF3OZquzQZLF6NZLmo2r2
abkJv3WhkSUjWBvovDOyCpTbVKGhyE7sAUAH986AO3JQG8qImXaFkf2By3nOxYvXIO2GnORPTqJK
IVtWVXbqjoGNcZ0EyYb1FyCQggzL+i+BIpVxtCmELjT84/lEt8PoT2pO7pEhZ36y1eqk4s1VKExp
jIG5ipT0IrX7SHiORN85G5RU7jJU2yxMEXzuymppbuX/DCSwyuAcVInh1RTrtogciGe2/6GTli6C
QFqggua0i34rvcyGdFvMY7wlKvDvGShjVxEWfworOVxIuOncSGmDGjBLgUfgu7Rosoa16BeyLB5h
eysSP360C310ZzcQ6xtJTzORT9NAZ2HZ9JaHzB6veSE/hwmBw0FRFxBG1nTyZCgwRHbqCLtyJXxh
zyVHMgsPzmlQl1kbGORxunkH75O9uzrVTNQA+ScspNubX3PPwjioMZa+lgyMbHKbngXHhtSV3mrT
Q/Ag15JjsecuY4ajqQJhqKHfyWXtsSkJDDnbagp3Ge1Q+RM6eEgMQbYMyBX8n6gLt721uTGDgpcm
lxmBIqBQShjzoZSAy9bKjJZ1fIZlfMKP8Jux/oA5ywKMJU8l6LI7ndWAiDQigZjEuKFiwi1BNXTD
ARqTx4c1AkBMDc8rHMobf9IuOq+N3ko4uGyohLEak/2uY1lIr/6BbdZ2H6ABW2YmSbaliWkDu6yG
4eBnBqj3B7pl6Aht1W9rM+Ecf1DXcQf95Yhf74pXVbW+c9lbKrWbXRuFanqcOYMjusEYZ4O2vWm8
lOLs10/CVfc0Pxz/n63IxDQtJJkU3oV0psL7dDWG/l7Lchkw6c1sziL5EG2wvSG3c+yMuWm4K4yd
IkeHJApCqNIsoj8wWF8mUlHRbz9/W91LC9FHYwU6AL5cH6F3PtFpt7iVI9xl3XrLTilY2XTGlQvB
AzIxAqVmuGon9nzZQ8M8bKxD5kfLmyQoY+t9HQVxGOuCvcRraG8LdVLBeSsj+96u+9Qj8WYNxXLD
wCCc9B7lbYNHmvtyy0AWsHDsWoalXfLiaXkfdyQQ9WV55sfBU6HaYvygCKGgPVyQUozU506xeQp8
hqJIA5yfWrTDX9MzwhryFWLKjmk/oAQVtERscKNZ7hc922yXvYZqMHleJEr2KIsl/Qdt9J4uVJ9I
n9JxbwzsbwpgDpTi6Il2NbvDhKZuaQ+mG0PkP5vTtrJeVfBfHLQsOkfm6IjKCqRLMMysqnFRgDSn
5ZpOGM3pk+3SfxCrW9l/MRUHph+13c9z/xEuf9YFFN/5MSSO/7Ht7U7PMyM3hfPD/Zyst1Ev0+7U
sU/chaXd3b85yifdFGcBQ0I/Isy3wrHW422uRqCCkgoGdG8Ij2Yh8MkAONIR7xV2EXzJ758rxnh5
twevfo0ufm0mBLImWI5DHaftLgqroK9O/98dgzzy4fvptk6wNDasnUE+b1KeZWZdRVSKcbNoJGAQ
h3UnafsoJQjtu3yZSz6XWp4ZZVqpLLaV5u+tJEiW8KmvMQ9Pp34xRkTN8WYTAkiT5BoOFLCI+FVO
7ej11gd6B4z94VtZyh6v9Ij6yqlR5ZJw2VOHIwqJJ58KzYqFIKgRxflU0G1iY2bVzcqxfIR92fDM
3iKLKJlazt8HvR4eO8Kd5LMM6ZIGGOd+DKIr0P8a0aa9PWT/+guDZWSFb7IYdqV+HYv5h4/w80sW
3ALIY96+l/SeAVEux6KuX+6VsrQcX60dtDXPeMiqdoN7XVXWpi+lALK/4vz5WELA2srR58jJt4kZ
px2X8lK9UJxf17u3he60dJ6yM65H2BxAIMJcH5X6tY0kCs5O5Hg+g5muBfoBtZwd1wrLel64anop
7e/7YHVytRAX6KYm1BekmGWSMyy9WGtgg/wtrn8i/nD8DWjQCJ6bDLPuM5srLWlWK/95dAkwtq/G
l1lPfw58XBpyak/xkvM0ORvF5Z0DrvClIMOsCqs8W1ucxEP1wB66zbaleJ8HlWam6Ed9rhJ32cgk
QnqENFPzLHJ2cOrJx4l10FEPTRGAH9VfJcG9mpbimGqBga2PecXWaPiI3TJlpHNJMs9yH5ukjsyv
wBDU+nVBDMd0f5Tt5+Y+QJuXWBlb6CjSHRxUDFn9FexdYnRPTqvpufdT2wumk30oqM2+nitbfIOM
18Tw80xfG29/21M4Dk1uYbdRlxytnY31aMTASYj2uT6A+4qzaFFiKTxpGN2Kw4Q3RTB2O6VRtKhq
hEwj21vV5BAxuWS780LeiZ2RpaQ8q3R3nKOjNsH1gaHoP6tuCrd42unADjscumab0m5574GzKS9r
Euxi9Ldkg18H7cLLJaexiXJo95LhE6fLrYwtolbpXmnoMq0THO3f7Xzn2f6C2y3qPbBRQZQ/dr9j
EhfL3F8mw7NsO9DnbEdDj3eM7En7uHie2ldz23Y2rxrNl8SA3Wgub5hoL2KkseDDUg2BqCzdNAd3
445a/VnOYesUs7IFGCRbavYnjauFZwBFCsJRc6hMxpSuF4sAsyJrsQRNWLk/qYfV0Hq4weZkTWTH
jSFLx/AH8SKs9vz2lvMb+zJ+3JDCAIbnKYppUDcvyb3WGsMHVgtzRSGTDXoqqFd/1EeqZPdwMSpZ
56oXi40F1+NrQv3pVPcY6lTY8g2tCrSDLJyvjdq8P79gPR8azc2r7ddjfBUKgNUb2nojUhwjhEN3
8vNCye5MRHifgq51CgwwjNzKpc1Bgw3qeOuSS604A1AQrGYA3rvqIpufzWx1euupoFkJ9YKEjB9l
bIOJ0Z9TfhLaoUXNbcRJD8PMOhMh55Wz19c3JspHupU85Je6l8QwLbRtg/qfndW/VnXz2Pe77AI5
jqyuOYTHSUGHzk1vXsiY/2H/hb4wnqGXQf/dhrcP8kqsSs3eBdP459VEtIJHKhXVSBDvGLh9Cm37
LiS8v5lIwV9UkvlfMfutEArHxjmLZsvXhaxJYCUhzIgSEhr8BG/++uDeKX7JSKIvZ1uHKw9e3bqi
0DK8hZIssRoGdaccDsTB9C3QbwG6H4gPrfyr4TPCQZRk7TCl1Kew622Eh/WK16488Wga/f+NrTtA
+j8+THJxoeJXyRPgchhKzZvQt0sjskd0HrbNJrmEKZR6DQMXKBDAqVFNbLAOCmufhcreLCu9GUdh
GJtGHPQkpn+UM6BDNHMpHdrEiLeYXvI1F08hHEXOMuHC7GSDjUxZpKKhtU4BxJXnycKfxpN0bS4b
UyH8qEeD/oDtMEUku/Jj06kRpAp6FOOqfTrMt1HaLCdO1UbDfxYZyp0GtscH4NRmQNa2Mk8FZWzq
O7JptymI6l19Hyozmw3U+aEqVVNthIayX2kFhNiwI1fI49jGtATfYMItHv8GHfr2SbzoBi/SBBVR
yb7nVQhi7cD0yZOHYE9xjU/lkXS+9+DgLDj8zStNbV6NvFQLGeNgDvs8PbkWlsK0kQN9Za9/4dAu
Cym05tU0D1T8vlrOReTs8dv5xveRpvvYc3aikSu8KIm8dxrv/UE2TdzWPKSpzueH8MmmMwWvtwGc
8cIkh9shFHbBodDxDx/cw4zU6lbD5w6ZHa4tASW5vlcdj56RsXeb6kn3UmnTj8++4agF7s2Qyt5S
hAid3GewbtLpuhKNt1OE2LjDMritIyTOZ1V++HSzdz3ipJNpHP2jvTZWKM2MxmtuXcoUHf88AkFb
1Ufi2N0ELWwdr4O5YDtG95owZ0hMiTE5nXymeSlWYGtIobm4/BTlLgx0Mi9aCisNC9C6C4JvFc3y
7K3Ntc4oXsgE45nIxj1HiL72oGr/tiw0pkcYrJGplsBHpiU/ksbTuvpPYCjLN/KhreqDOXCY6pL2
IP1/r9iZAfEF2iGw2RJp87SGrmmBfBa1LvjBWo/h0AlMqqGSaNAn7YzM9ifTYECNn+64N5TvuP2F
s2s4til2sLYlEgfL2bK+U+AXWVnxU2usgW737FI4ktvdTb9lI4haITni8Ykwme7sR1f2mhdEnz42
4DmrMo4VE5mukIw0pPyXW07ag287fpWyoj250jKuxJGw8mnN97O/KQW6aCxaH0OHytp4vsiDSgmY
KAbnBIFVNDO0Iu4wZtLB0buG5VeBthUzPWF8P5QtR78Qs5HCUekpx3xp8VFafQ+dLVF/cacR2BTG
hE7OVZcxdV5M3AfKu0c5X/ylxwIWkFSVk2Qu8/DGgAc3xa7sF/x5KgC4geHRE/oMkjUJYGcHIdi2
hk8gqzD14MOEIPcSH98Lh9pGXKB1JY7FwGOGXBd4F0tXs9lLbpHuperLXxPyR058UKpfEESn6ynf
KdwHjuEgxZEqV1W/gflm5b8uqfoUYthUgzE4UhdX10U+EV3y9bfJRoPZvwMigcWbUbjj7yNlCvoo
IxMHfrbio4Ky1HibnA3m26TIywFMYmpN7CACpHm8tMJAdu0Ah1uUU0mzO00je/kZcltzTS0g+uBo
rhsxClYIFUE1wrWKUPax1qUxKTZCx446pCL/VhDpcyQriNYNNWVT3XaAWd4MMfk8mlMrT5BLoCt4
LLV/taJdKEAJL14vx9IMYumLp2JTbxVBuTPZMTrv/qGIPxgOBBlMLQl6Bw0ysX5CK1aNT6AHwflo
7P6lF29dHdrwEDf0Pv3k7ux/QS6jCOTyNJyV4ZeO0ZM73OagnVRgdJNwSSeNRWMDHm8Z6AQpdkVM
YQJyhgMIst1Fspv6MMxTwTxhbyks3flVclNPOm6lOqFsxua1auhcJCR4jeLTH+WkcW6vs/zN4SmW
WQqkRe8w3J8FU8pv2+nQ1BH1OpyoKeXeYYnPAJRAczm4zrIokBxXJui9x75LYqULsCMb/QFR5pII
eX32rOVoqEgWQD1T0DVMHxJC7598usVQ8uLhOE3QH4aqVhoQbaSG1BTYLpmf8ulYmb5cXAH1BXEc
HejHrg0QspRQGnm2urVJVh8GpoApW/qcXu/Z2aOqQDMF8vJvxibLpsX6d/JwT5uKTHg/XU4glUs4
qVX6a2t+S7+xRToWYYBjNXWAf1GphT67nerh5yjkKCNgwHoTLIX3TXcOg5ODbKouSNvdqqpSWyz4
NGxpDJU/wGJCGpuTyL42+o/eBUh5xD4ZUgRRvt2o5xc3hzQjrIrOnZZUQkjstpWfAE1WoImJ7bHr
6Qn8DAiuBkUdpI0rF4x3YOlymaCQUL1Jk9PXqAEdpH922KsfqVso3lhe0mjPjSdfiKCKBNbVxg5P
rTCfNagRxCMSfHVfq0B3wYZ6ZL5LNJ9u9espqDE5iQZ/ja+pGNJPd5Zz2RUU8Ik6HYDIe7h/AtuQ
2JwNw09WZpYR86S5/V/uK3hXFScJqOuzBL0yLs1XV181X0mIVPeRnsneUdU5WF4jJAEnMXrXHBtd
hkyekGoQwGGDjgYddEkKannwgEGuKZEgsCT3jCSO9e3XzjH8VcjmQ7BntYA23/UkUww+AgXyw2EN
QuPWKYjYb+B3m52x1bXGeuZErNSdAAsMYvyD2D8bmChaFySHVgB6eMBBdFignDvb1bsH/BLWY0oo
rJX+J6WWXhQbLlL15kU9F0y23G63PfbNR1tb5sG+Md7ZjrLALzOsKW7WuD6V6HlnOoYNmIKcd3Ti
/ckGjIG7FQ3kpRBn8juqZ8JwgEb4OQx1jVVCc7VJGCvl0mZBOHpqkvmyskJ3pkIjo+xq2dksjR+Q
TpDptzzPmj3FfXs5teGFJ+UwVyV0Um7DqOZ5keH2f/Ga4fse2jmcvQw6JseEz9a2ItwPxQA+H+hW
BWLIesRp+yFy39FKx4QtpltsHM0699PVaToy7ja4m7SxmN3Qw3EzGXsPojUwXpdidQ2fQlND4Dom
ddSuFubLQkzc3y1IoUvTv39gaoMwKLr1Wg6+JbSvVSb2rdoe88QUYWui9kflpiL/7ATMrXNzSuly
pq9zKcWXndVFx4fHse+fxzc6FBjL/+hCv7zu6j8f/6AKAGWx4JYXNEw688dl1WECH6EZ4+c50ZZ3
+e2eUnkKUd9jCreG5Cpe0YuXYdkoQKc3A5+qBJfk1HMzanqDCSPKKeWVk2fqH1aR5GIw1RuSUxZ4
iOjGXicCs4dXGy3rWytfzhNwr2qIXPzl3AcMKFDnvnZoMi435uVpyMLjBMOOrQ26K9RfrLh2UVG9
k4N12zEL+VNwohlCxOHUyaQA6VJ2TI+ENMHz9QXV4OaGW+Aia5ukY8HPXF17CPgbpBREWG5c9NFd
mkg3lqvoKWNsI41m7rSmbDAjuQ/V+2BjQvpo55gvt/ooDwildd9OsCC1pG/na/bEECZUH4ZGLYvJ
TmrOzvQ9pdFFM/hXpz2SOjdPfrQV7anhxbhk3uzLrfiARywUoiIkYGYLj4c4cTw9lbwTgP/NKhEZ
sljg1eQNDk2SMjMoktMuAtwf3Kd1NJnZUMy1lLaaHuU26cMAibHuaW4h2GQngM0KwYSpyRY2zJjb
n4Bp3AqJS7EkIaU0bGmqh12NVikCpf4QRButbDiCzZjfr7h99evsmv6zpFHp6dmyCUDxZIsCDlKp
wwyCbgqGxxTnEUToXZ7iZlLoIF3rx0W+Rw+myEQYEgi8BF0BP09MAAEKqYWnCfUzJV4u5Lf/XMg7
4SEykRQM6/21oMFpa6w2yvnWHvGg5HOY6igwWpm0hiPdzX6ltw1A5E6DmTmsfjwBoq8+R2XLbK/Z
Fl18xB7Fr9xJj9djB56rKt/AZbjG/foKp9qMU+UdUQ9S77UsoB7N3l0UeVaFH7MP5trNtUiXxA8K
4JTifHsn7yf50RcxisdAXT6bQ3i9mKzgDL0osZojLZPk6b8GiUPxlZBhR7CXHDJhsIos4Wa9wN2s
egwK5ai7T3LUStv24fCjreojh+yzovWkytq1mLmRicZfpEhqu7lcheuTIb3NgIymKkHPeoAfVrbR
Jq/io24hkkU/dp6f1s+ZTFC3Z0A/1+JPMNJofkhzo6VbRX6MFFDiEwE7DHVCLTxSw6YVYFhhaTb5
DcG0ETTvNiQskkNHpNXxO9vAD7oPerajuDE+6sl1DnrlkwSwDPt+CIJOFcWaES4GI7kvx/Q0cysk
3b/ooVV2200j9QNt0uYkLlynz63AlV2jJnwZmP80VrN5Nd8rMQV7latg295+TQzNsBqMx1eisb8i
e7aBkbuQ5cYN1nWCAauWwj+9oQjO4iaSw0fz538kH09SyC81uVizulRrRyz73ll22cvHNrtqBzxY
hfsWGNaMK8iDP5g2Gs91pBl4HFYqLHG/8sB5LnlJbBhtMD/mT7KxePCDM0iRiO6gRt+DYpQBtr1G
3nkAdr0cqoR+J/vVJy0pDT0saR7CUA+JkbM097CiJEOMWBru5Lzefe1EXJXraH4lGY4Am7eLn4U1
+Nz7+MU2TzRXbBnpcODhK0KikzBoZ2vZtvfIpm8bnUiv4Y42bChVDiBvbvsOGQjO3kLQkaB60PSW
TJDveUjHaAEQvT+r4Ol6WK6svD7QY87QbpNrbsUzSCBOtSecARbsPOS0OhF6wc63CwO1Bdmr3vA3
JlXJPqIeAITFoftSKIDfQMsDL995oCt5fBwlykU6Q6UVKQNpIKyEX4ZWLajVgAbXxlHj4ZVOhTE5
7w9ilYqlD90AD94/fGrwME8dhSIcbSnQ64uYtmJPXdL2glae00NHSViC44GS2DNNn6D+0/umjEWj
A9ZFZ+ZVjN//YHgEWUP80rQBJDsVqzQ6kNZomYSEBSgBqarbz4rPGuvEBlAJkirlHjEFt/uPnnfw
dxDt2p+8pTXpzz0+ppC+SSmJDeJvXZKKtOJuhNZG2hyVJV9KQXFZu2cURV/lcZcmWNKzhK5E3t/M
IlD6Q/HVp83IAY21VXu3xsF+bNrLvFZegy5EMHaZNpRpRpACqIdVwob8F2q0vBlEH5XwfloRAGlf
iSpP296UcEAIPBQ15KCcL+L4hsPErLS8Uk+vPTGSmfw7f0Z6Huem32n0d8yXdQPUAxA7yZQVrOjP
KQ6uOG926zP3BXSWq31d4xkUM4qiw6RJIkgrT7nZUUmYX2A1Ekdg9mWh3AN80orhInNS4Gt3iRQH
vEKqj+CNuw0W6mhsnNF3pbnQ18X+zat20j60kSb2blPshrtty5NDvEnI4oTXrnv2tRbTx4AnWmPX
j1pf4igVdHZANber3/Kb0GdqiG1GqdBFnt7JF9P+e+lsjS2rqXsoCSs5oO4gHe8jIRFehyMBVN8U
ZPDWhcSTsS/J1XFF0d67Kg9zpMVnropy/dyRTmAwrss7O4thsMii3p2SshXtdP70xr1vzwqQ5Eh6
OSdgMlXmVcygUi7vj7lAVGFsHKQgOCDNLHOucmxK9cGTjYJxLgezkw3Jedw6q78DeL9tjZfe9DHK
wTlBoDZhbI4tucfQiz1u8+MIk+AF5Tg3acje0wuBbOt3EgKncm5ghamrkebov5ceER7+Zg62X4aK
MpaEY+az0wJ1umxp8NJUQFSw2kEhQ/94BTF2wXIAwKCmn9RZ1ld6gHYnS9+nLlcAx4GTOZ3uiQjL
s5aw3Hp9fQnz4jY6NQM1tj3LgfBsBiPwdwvS3CbT8PWr/TZsfoH4Vz7THfXRxNGo6G4AjKTiBnHJ
70Jd206rX+bItiRETru38LhpXOX5rUNB9Xe+Rn25IN0jzShgTbVZAOBKrTry2cF+GhzmOxYeUTRc
cqYcFLlYQBzzCtNCJktwvh6dgqDnGjKa9D0rysvlaJH5EHK3GHhF6LEfxy0RI+B2z5aPPXLrnJAp
N0fI7Lz4ASvidSWHDpuPBcLo+Yy4MGj/Fvn1MwlOQNHUJtWL5RTMxJjrfR47xRIcS3QBWQ4bha0F
RpomJkIqB5BQk43Iw8osH8t/zpH2PcPhms8475RZeURy9t9qgpBVILskuOoxfofvVlTttYIoq58K
+tIOHWrYMxFcuxmUbHIMbOjIt4Wni96JWQE2XZhIzJ+bz740dhM3+/7QwLlnuqBf186992UgWKzv
4zZDXgIRJk1UkCaOSoN9h1BGdv4s+GJdeSLx3jAfFdFKpjdMMGErnjP3Y4oSFPfTAo5U9pNLHK7t
liP12y5qA4RI1/F35GPg69oWVGOkHI98Quy9UHelaPRw+x2mltgjjFIfT/VKusxS/ezU1y2wbVXk
YCmFplXm/hiKoE0anFQ2aAlBarElCWBQW/ryde+bQUf/HtwUjM1ytkkSUdpOCc0gFj8Cpso3edLc
Zpq+AncxZb3p6h93Oxvo4ykodsw+b1vNJO+u8iDgRdUggLp/O1701KnVWVv28c2DNKqtFAsJ0qvw
8RGM05Jdw1zyb4Qpo8N+qoAjMs/AmdE8vDNpiMwNIq2zxEVIMlN6OCgbhMy534QRTPI5T2XnU9jN
zl8FV6EraByMJvOUbnjBLhhPV4eXvRCJ/2w5CXDfV92G+W1hj7RcErMyDylXU926ojNnvFK9XBOm
F0gIv2JI0h2TJFLwLNqw7SkvwufWfR1oQfU++TDGSp0lj9dCPZMip+r8is5KC7AxvkXmxrL2wMwJ
hwhBaFyN7wjPC87TJB/pdW//potS77gNxQ3mBbk35OOQ9xoZU+x4nTr/iiOqPyr/7C7FS0LBMVXK
pFDvSk98jDU2MVPOrh9gB7iX3Lt8uCsKw8N1wD9U/aOT7YkoL1WyGNm+J6VcFtV6ppTXyOIpTODH
nzHwiBA+JIWoGnGoCJMm3Nm2RWKLFqsuQrgq694E6jPtawqoOvQDVU23N47rlHdrl/e7prPCuwNi
mSx0wSjJNiGGSD+JtW/K+LEkjoCLP4iBYisII1pNILyldCmgLdPzg9bs5o8t+hBASREthq7aD+2z
Ditr7Nq0tSmMutBeDcD4xFGZFXzGaZ8omxg+EomEhmjU/Pamv7NVN7xm+fFsWQdfA7V8AvFsIQYV
5N79W2iC5eAU/t2EaRv5Cpp9dNfAZcPlVWJZ03XS5sX3IKUkyKkJ0wP4P5/dPowGEuWWE+/XCzL/
DfSH1pDUovPv1c4W/Jwk7g5ujYopSYlpShEVELYB+//x5LMdoTtIhxrzmBJCKbHBemWgurXRSzEL
gE/ttf89hElHAr/T1vx0pPVwXkjcaJdt+UxPhp0lcWmXopuTxru3Jlf2nWWDiSXyxxySsoTlzvtY
upzJqLEueYQ7ZyPzYYscNXT+tN6Kq03pG3tBfkTf8oRkNpoQyjVIiU+8V+SeZrO11yFoOpkrTU2i
vz76ksK0WVoiU2nE/sFuna/g4WWQlt7l1xo/a6si223yHgi7GUmCMZKy1mvvOa8fbywC35fi62RT
J5k+p83YzFQB2caVxypmw4x0aMTbKa2jtkL/NM+AifhTDwrfujld2KxuZQHbs3xSZyILIHCAbHuB
3EJ6dBiHwo49oyTUDGBIP5scqtJZvSyFbwDOZHb8nI1rP6A76sJx8Nyw/9694hRe4zfteiafRdtR
BAUcE/wPtZq1f9zrbPTa/gNn5R2nsYDTlzQHyAIal4qC27soR71ZMrgilxnR5cM4epSxkc2M8QVf
Q7k6shoEQmeP6p6fwccwldxInjMqtFbnOQpAWa7TFIVY6CeWoXfkM9he7TjsiO0bBmqhjrctOpBI
/QF++X6BsP3CyWj9KZ/RIiwzKFmBDxhPnAzDEWFa/BmuNry76zpakEYsQxFBUr//8iVciwUnNRW5
mucl/cFYXaNgMERT0LT472CkirfRJqY8N6r7gnyRrxtZzWSQduHNEJMDiWLarho2h4+R5ICGgWxv
wMiQrUTt2xKnU24OucJIyqRCfK2Z1XfolXbztUbGw2v1Urj56zngjFlHmguGBnHrn9Syhcg2LCds
ejQDu9/+sCdKAFaJUEtOTVQ4zD3zTySFJg9SsWqB+4I7BWFlfsDUJbDOUHF42VG5MXuYd+vRtR9x
6NwZrM54Ag0cjfNNqLs1XZMXWP4W79e/tpIod23VMcHC/aA6Vlhu3EyzwuBDzP76gFghuNmZpe65
UCcd/HM2lDVDlY+144csoJyZ+TGkTwBgUIFg+ZDFn5BAki4SiGCtDMxp+Dau+ELDIuXbGz0Lugll
cMad4N97OBj7PLEGV7JwuJO/BN9BUvBYfTixDDy/bg3t0WmGZG2YdmMeGdA+myRnOsOA9AJjRhkQ
gt1/wYm+N+Jln7G8wTjW/q8C8sSWfMyamRTJezZscb4BgRfT6vZfE6l+5Rylk4lMJkemH/x6GRGy
HJPm9cujOAyC6k2b4i/Rh9Qx7YjiNOMq3dHVCB5S+n8RMnD7/LHDNT/NoO8WwBaiPNoKajp6ponK
fPUy8B9rardYZbYOncuKbZPX9TMB9Y1RzKGpfQZs0pTM5cL9dUy7z0RAkged8uhSmxXCxezK2CQp
GH9+yjnRgTzkbqCLXOI3DOVUgMvXlo8ahXi+StthSwXKZAfDhow/crqv7J1UAlrsy7VSvl0i8xMU
9epq11JsIGiL89yo4INMhVTdxrq1/fQaiSpYAOfpRx4ve0fyjI8zxN21a737BHFX6BfjL5v9hzho
/6azOtir+uIP9OFnABF8YDmAdUnoVf8L/piG3Id8cT1VNV1m8pav8Cv03BNb5DYL9kVAOkqxUimS
+omJV2KHyLdwsZdlvtDYu+KPXBElrppiVl04pCzJJ0PlHhWCV//QkbKNDpY26C7iyFvdludKm1+U
ceNGrxn62NzFMdy3mOrICXn2GQE+abunqLVy51A2BRqN5FQuZWQDtsiqsSIVxkpOesgNnsIHRE6q
H8+y0iGwKfomEzXrDE3mZMgsmZa17kwIRyhLwLwfYSWTKa/oFP5JtwwsQQlkF8mF39u4NKAXk2Aa
OdkK4xAGj+y6eLhZU8Cuit50wD3up+7yt4kMpr+5DweL1g8ysheWWUUcSNScgYGSp4RYIFMeIZpo
l+yLei5g4TaNr+8NFYFTKo9zwMUewo2fLL9m0N9+d6ARlzTZ/KuDynBnvqlsoU8pJuyUFL/CrDAP
eo5HkgP4qZAxB8fLNEE0Esc5mzwX7uO4qUn93KRNOQubfXxZwbJZTxLd83giH53XhBL4XRzwWbFT
74GrwRUxWPbcKWgyK5iFnHfknflQ+v756lGPLlI46wSL4vSLTY2FammvNWPCL4MNtPpzFTjfUbrL
dalhOAO5694AhB8NRd0M3FnWeOGAQj7KrhZh/60w4y3RMVbTLfJX2AhIDTL08Y8IibOlkvp9FLSr
MI9Uof/iUbJerA74dQGmHrQ+FN9B02XuCwU3D8awU9y9GDqDy9+TGegueyNOLh7nieUHigIH3QKv
1G8iaTXeWO1MB/W0iR1Gu+jnpSvQTHu4u/g7VycqadgtrqhBJ1IEhIjxkTulFbz12C3l8bbOlIxo
LSG9CYod8pCsnsw1K948rLGDy69DiEzbBY2O/URFIsswNpNNqb+LdDrXO7KaV43lIaodZpWlOsFr
eGS+OWCeWe/LjVLzIhQiekhYQ3PwU2wa9KPwmGLhztBDH2pkhwIsJt0RQ9jy/xIQa//a4ECyOWsZ
7igJ/++JG927uSh7latJjU5/4P54OYgwZPw6dLDUQ7nrm+afoDIRgHvz9OTlB4ov7b1/etnL0VRj
F6YagthG1hFf3ovUZik2nwtEvdSMaywpTufkV2wq5DT6InX4l0KUTvNhyKZxNUmYLxtPGFd/pPC6
RunCi5iB2/fdIIauGGJ9yhDYH90u/V9ONSJGOK7wkY6BdKdKK5TQ0tS0crONsA7TQgWI3+LrtRyp
bAejmHmRxTB3ti8BKBvznqBN9YapTCbB5mZBS/KtM4JR+uI50JfvUvpauLcnXQ5TFGpZbEHpOlcl
OyNuySBvCTv2wzgk3Qk/4H4tset1A7/Mdp5LYqORsf9k55Z5At+4lxgMs1jjSDpKHoWGCOAYK146
VRq/fWaEcaHQbrKqTQ+6908JQbZfhgYWvALuSlDzq0NtYmIn/zZjwreIggNP/mQBfymh8Z8ephml
kq387uK8E51b1GANDUaRoEbhMGYTz1tL0qK/hqL0C4B4J6fsNb5bkkEYmxv6H9fKUxJPxh/nSZ/D
GgBA1v2ySQZxNcTKEsX/7mmUz64+nr6lJ4V0DerZzjs5wXaJjoQ/WNwpQ5sExojsYaZtHZvtHTCf
/h3nsKO+OiRWzZPwcj/WoUkke4RjHuPbCQfqAmfUA7qiAqDNZKTS22EK++b4AbZT5f9Fjv46uzuD
SHZj4Xqy11hMii4PFZeR+0CtyfIhbXNoqQckeswM6tg37oMObV7C6sfJtKTssHeWc2S71TE1gsRT
rq7KLPKsT9xDdFK7DXkYynVI/TPy3fXkTrz8auDS28ZEzTcmHRTI1q/5ErGTgyvLu6v7tL4UctT1
HEFUrCFNF5kRvpwAB1mJHdPiouhXJOjb1IHy6auVR1kAMBF4aceioCRSNN9YdmWyLH+RRn9XHxjT
9VhrcHGSnDlba18GyHEVOHewyRSKBEMVSH6evWfwb4f7zq9UR2pgjgotPwBhPjUr3iOi57rn8THD
+JG55DUQjsodovZ0FZRgZ9x9H5vZu95i/Jxv5bR2gDKxOk3yuUjWu+nw6EWiWSQ/AsooiCUjIXZ7
KI6uMsh3O0VD2ju+vy28GHa475J0bevxcSzi++On5l5HQTsZE7PAd+erpybTFYj9RKXHfdo1zy35
koDfJmVXg+4KZHfyJuhSGBIcHrjESjXOjvBJxVW3v0ovLeaWFyZ0x8/B/WzlYMr86qHFHCAfakJJ
muBECUOA94BtcQxtUdELnMwOByC+1lD1zTvigmiD1d5v6XcJoZT3kdk3QsVYDz2Ih+2eEnePpBk1
dGgAxakmvLYgpcAAhOqEZZwtijpU8zM0xPdAdbhFDD1TeQ+Hqsrku2h7VXQp4QSHHF4lIRFHFFns
f1qTeGFyc3LSMFs7kRDgBX71s1rSoyuTS5hHua1CNeX3Ms6ZkOIjm8y6RhmjgEonno6oBd8hSYPo
6yvHZjnPhHVZXP+iqdouOqDk9ihO62OZgw2qWFM6907xlt2AGdDelfQr79nnljMrokCmwRxASShH
66GsgEYw6PM5CknM572K2D0NVIhdsPZX4HRba0IghdYdgerfjBoLqnxN/M7See12/VHi5aJa3HfB
grIp/xksIeabcP4uH6jVtta5RtuRRlh/e9NxEJUK2qXVgV1D/jEBc8vBQ3Jvp4FFrqZzNT1LTuO+
CyWaZqBnX1vumxHOD10uCdlePv9NqQFOFic951vnB1SBsWuQwBIVJkYktv9dkAVvJzpCaloUngP0
r9cxQYF3Aua5OAwib0yhK7/iQ154IOUF3Rdzid9zM0ts+aOPkjnas4toqZmtOSrUDEXRA31UuFhx
p7vvOTi4U9ouoD07gxEpkFJXLcM2vk5oYeUkrarRqGLmFThApW/uWx/uA3zNAugaenodQ0zcWsCV
eAWGntdxHJGvF+ux4yDxBYAuJlG3gdD0uXImnqH/YL8ddNn7tbYxd4AdUVWcZJmeZUndX8sYQjT1
zzvO3tF5Y7eVKfq/sZZ85CD8yK+m9Eom2TZgr26orua2IkRynhXQ4n8U/vTpK728Pf7BmF5ISFxS
xFRPESve0EsthJFWRQExshKVMEgd36YpXuO5L9aACqFM+2VFMnm1Hov1LshkvVKtVL2MvcThuXnp
AJtyuKxKliN0qbzFp7kEpYrdtPp/RoKi9LKO+euzXTzS8KUTTfpnpqdnByI/EDctYm6FA6oFEDMe
h9tDMe5jg+kpSMfP8sA0BpQtQ9kFT9EE03JLAXu2o8+41eLjjUmUgr6DKMgdrG8o5RNz3+mvCFmQ
D0bHUEXUolxqI12TQLgA/9Ns623dXy3VxkQr5zd9+3Cm9W+YO4jvm38K6NmgjK9uSxFxHg1Qjiae
FuABoVBaeomYJsIIg7d4nbTJgYSEYMMjITk6vinrToYnk4PW7gpfwximpIfdXa5PmgK0NVAb/gY8
TX6HxMb8fsrj+YBVQhmhGRQlKXUgdFi9KKse0rKDkLGr8LwB/TD2VJBmiIhxbdL2P+qg1e4WhVfY
0p/YhpxXEFy6Jhe0xpEcp/N8S5oS4hwripmNW/KTVqnVqSQ8QXoXmHDYFFodEWn63nzsBpmq8Aym
BLPeyfBqH9A9NLCd755dJh16NOx7SvClzM9EfRw02Pw24DqjNOcscnqYsT8n1Gxp5kIpdS8l8K59
TmOMOdo2ctoYWwyWoa2o0A3RmrKyZCoH5WmMk6i2T5mA7kHJe+HJyw8jWC+FMsdaIqRkTJIXaw8v
+bfYUubmVD640m9dXs/0ZnpIXRYIEH82zaHI9odHMEvB6aNmRX+vUp4af5URj8EU6QJKZUJrtACh
U29+tZ+gSGkQh8Qqj78hzmgWeoImxxGrFVD/Sn9xuOZxXmr+lgnyM+86CfpnS1BS3CugpxnT7F/u
/NJsPQUDMTXqNL2ioonet1tCXpzv8WTygBk0HfROlqlEKo58SfiMJU3Z5boKyGN/cpV2uiTNH5RW
p517TNPt4vWAGqHtpHpgucM1vmx3v1NjSzGDWf4F3LuUI4xBnMdEmBpaCxWKn2IjQLtjZBH8GgW1
xtX1WlZ5X2QxXQOvh+0sx1w9elG17Pn3hXUFdgIXmdjINdt66gbs6TW0reJa8nn3qmNZKrvBTA3g
MovoZjysaCxJdAmOT4CilHAG431NF+b3pXNk+X95J7hbv91uErZn1ypuYynCBt2U7FzBSfmZjIhd
IXlghaTlwwno5YA5vQa5FgB4gGHyIzZX1d+z3OwgE3wkkZVJdNgPRPRULWpRp/leCJ9cAquSNTYw
X/KBEcM/O4mozJOMf2/aFKSznbI1TOeTr+oiVJQ8Lv/+Tr2hZKqKZIm3MHcZxCRDgBH2XWJGrjL/
eEKEdJIPM03ot0d9LJxhboxIoQk2XP4w88MIEgijRiBB/qNe7or2ky6NvPSAwjfXy3uXoQMxyzHW
XPA519Hmh5wUxWpJ891qhtVni1ALpaHwQfMRJyo8UkD5je5x7UnLRhf1thBP//i4i94jrwHw3gmO
Mymy5lNI8439JHo3wXcXGm3HzJJKtkg7PfMRJRVSo5+y+1Urk9ufB+ebA4AxxDx4dPCusKtDO0FM
zvQCEXgCmfYkoobxxnzRYd9joylx1VF7F+054i0IZSecVn4IklSmcArM3ILl7Jca5k18Fv2zabBn
/ZDVqKVKl3KPXur4Key/AJTEMHyACZGz4rCt9JXJvtpaLzMc4gguJYhFwc3PdNuxme1fgwOl5+4v
+ZjrgBvcbc35dPvCAyIEWZ6FeS8vA3EnU5UQoceh38j3DAFNFlaKhnsFp0mkOPlzL0j3qG8Pt4ny
LGllM/088zE5JBIfpXcjXz0+ugBXPd7Pd3eOCjXagKklz4+b3bbSztmShLlYNEoRSMLKBX+minx3
SGzyiPn/prpWYuyJgDlmMGdWsvMvv4SRGHaVqhEtFoM2NNtstFv0kdLGSfMOMyG5/lg+xkxx9ozz
GtbRS6NcaXxEQ63El2wRWBEeFi6RZ1Vx36cjxshD9KuNTKnFqfHko6jKNw7lw808Lvl15IVYZTf5
hlxNczh1o7i6ZYHEVim2/c8dbYjXzEontEyY3/4ipAbZr9BdtTomOpDNC/kzddzqF7L4zrBZ4qIE
Tfgmz0aTY99q0iC/gDzC+yS4sKRvbG8TGBTb6GiMyGZsEOnfj6JZUJj8nowwLaK+efalOIO1rwbM
oO1EhKszUyLvTgsJffvK2+ryvbTCUWd4wUWBX9KZ9tyiN0UMZNAPv6++okHG4VN6HJqeW/WkNzDD
drD9fgCY+gCQBnhTObr+XSomjQ6+zvN3RYSUzzrf0A8Blb4WL+xkY7HZYyNTy6aEc9CTclaFZxFA
EV/8N34RISL2aLiwFYVgGZwXlWctIscJdsimi1/Fg0AgGDtW6QOaySWPuQNWtIWdZNHl0qkOf0Q5
r4nsN1YIzQmvNgxDyIf+ic8t9xam6E/elFySe3kWMyWhcjqE4MHx6ox11lcJHfSTH6HPriORVf3U
bZK3TRYYnk40+r5ymKxBE1uaX9AM3b/Nv1/9oD1X43f2QNgyEMFdISTDHFV6Phcugw0l5X2QeKhX
ZKsjBn91gmcpB8RH4FON3GivzK+kIibq0ldWkS7lrFdqDXF7UTJgZ8EfI5vVdqvUBuFO5kbVJ5cX
HJLgsgqKD0mHyUh77xLvUuUfHLRv2+X0qR97/CSqxLLkBWLow/kod+p6jbGxdtG32q1Apdm/lsze
x5+rSe4G6+iySotMJNbJApGlhIr1NcfXSRo440qdtmAn/HPpqL341JY5fVelJ7HOwtT4mGSOFsoy
ReMHeOms3RP5wljoy7rn/cGOjLU8K7Q3+eiSCEL/HQOqlEPUtUvQzH+TwxxWTATkbFwNCNvPozCI
3MoU+aMvXLtsv691moSuJ/8k75jhLfGWbXWSRrdB9imXT79lL0EsK3/4mezP355wMp42WluJ9l3Y
t7cXGl1IT8kaTHa7QX7ZgOxslthe1NSiyt7X2r581zTNzeTDsuas90hUw0sJC3VrN/Zxh/tjoii6
m0ZpBzl9PNwey4konjxdtire972rWC2DX6fQRQHfuf1hrGxNYaSLJVNA0ffcW/q2EGj2K6oOGGFy
v73kCO0pluBnvLeq3txwh+OedgWgg3J2V8Rmhgd+rHeI3ayU9F93zxGiTEmvW5+1C2wLyNtaT96k
MxMVWtmHvkeNREK2RgEqvxJ2USlW4xy7uH5ePXpKfkGECuKNSYf/73mrPpOjkJvqPhywqKyfRNYJ
pQzxeAeeB7R5o/UHMyqcHGM2VCYJi8wnazybjWP0YLdAoAVfwUFEsIi4sjE8KXvEeMk6dnMaa5XL
pwMMXinREAeTuifmagVEXRws0dPP72JX8rBiRjNfk0gj8KEMFSTOb9KlVkRbXS79p6KN/+vFollr
js9Pql+aXhHMwGHVn4qLDxzJ7CCafDznPkUCdWHWZtWClUI+UnEFIftxS+9o2Q8iTgx5yrewOdd+
S7x6d09tgC4Ywi9aeHkiHlrsHlyBmAP8YRNExiXm2KBZWmW0ihYqRBK/mr5F4acBTU+TIkFPj2GO
SPKo08/a1gLJmoKBWRhrMofX7/sk/Wi7fL5k+BDhlaVNhsxeycJZ6/RsnaQjEehjPdd0c92pH5Hd
Si/u1j96yNdjEeAl4w/0ujW0N+nTamF0+U5pFn+JN+UigP4bqMJEXbU8P79Y+qWsZ8As50Mf5Tbi
G5zLNzCnbyo1bfEq3Aloz2ibZMth/xm05oSLM3GvrcfNXJ//SrLA/Q7M1VlSmOiGy4YPVUeuKq0F
Bs+Qp7lwYfkzSKFjmyjS4UOqV0lbbICSVlzjh0COdF9YEISkw5hKtDv3nfJsTksmsScmSpcRe/U7
b3nIkokwIbml5im3r9JNsnJHZPC7cLhPMacxbvJfpUOMlSmHK+fk9w9K3/DKETjziRLqj8diBIRg
Q5cdqS73sJpKRdL+eI0uLkzWjYRcePDRVd/N4pwiamNOh8M2zaKASlyVJUmrm9FZeC9k4BLUP9bp
3BgLSYaqtZTj8vO+12C6ntPXYVwWmnyOFpt/XQ51B7fqWAJi9bmk4WHcMtMamj8Eh1gwIX/dPCzZ
dYzyvm1PShHkWf6cvWT562wALwMUG2QHOec+Kv24jDpEcbr4ffaeMmFCFbPub9cpn09x6+GBuZzt
QjyHCgzsbMeLTCH2woo7fWAW0MBpoZp2KsZYHpi5GbOUJsjPOSaCgfJ3XRhtqwXAsjfmulz3wcXh
OzatPmGdxvRKgY1L7X00v9S8bgdxxFYczNHiIW0nzt+ufw29OrY19hJON4eY7fbq/ElPdtc4w5W+
kYcd9YLFGnzzWAFbIAH4+/Y9eMAnQMCLTl2Eh+jr+YyPxi/osAd8WJG3fGbx5wHUOKgVVnrnMg+M
RGcO6jzpH5/maCCgW5vnJm9iql5tQfs0Yf1OwIGJZsgpic0D+gxPezZjWeEiCgKl/BJU6FCh8Sse
gmI3BXeVUQrmJXU93p2DL6oiOsflHqzhI9UR7hyAeZ8lKPkLmdRSrq3tEtpy3NsV6YSuA1FMwcQI
hJpfQczwQ1PAorttNLvgkG2uNkHIm1MCMeud5Iu+/yP172wkXIjXDHetT54FqL0NqANDd1GWA7Kt
vEPzMl+H2jD5o7Xv8fAbFU6/O4vLtiPuLPh8ypBYJmgkwQjd4lV4X6pFFPuqwgUYEgSfz6uxzIdz
PC5V53qLq0athIc+2K6OMCOnW4/RywSGxeEzoUHCwQH2REY40BiKSUjD13nl1DGut6QTNb8URrWI
zjlExJcTV2JRvmMZb9ZL+rUPimSfeGJrrdiQtCJJasqh0mw+TdeRKGdjZWSdDeiHqaOpKxfkDtei
ntKoAkJPUr++tznwgBfU/+leE/ddEWl6d22nSAEun6ScT7rCS0Mls7FiU/RzuKd74dppWBBGlmvd
kr2JwW3f6+eXxsoZD7okzyRcNxvl56mmU6bE5xvd2zolJj+Zdf5hvP4xWr7X7eyXvFjKDjLi5+9U
3m4cKafSNRmZQFhjbf+cGQYvUHgqEnzYhqvoUS64ALJjtxUO99OM84m61R6/1lVGb4v9FixHa7Zx
QOmFob3mSopFArYtev+WsmTl0bBZOfY+ZoPsd17s1fnmuR7VRiGPmlpp8U82yr67XEzZTDvh/WFh
ZkdfU0SUwjg4e6FiUzWTDKOMGpA/trry/DVYhHn5XR5x5gJ8CZjPWPpTOKp+OVkbCigjfjFGR/FH
4L8cgSbczY/P3ZlZFIOav/If33nKkDUcK22KBgCYz0OO/I5C6AYfBH8ZezDu+7JCF+VDYssrtk2U
+rUQdq3gxURZg+3UDDPA+7NnklraH2PdWrFD7irQjckwdx6DBUkJSAo0roleDDi+GcBaoSYXnbEx
3WI/w4H/2w4C/62Sj28o7is6xw/SVbzekS5kNqYqgC19XFmy2uSpECX74jCDcxlAfL9YyorzlVI1
79b2berh9f/Okan6tdy9k1AQt32Uo204M9yfAqsbR5NRLsVUD0d4jmma/X3umFIAl2StpTh7JfzK
xvWqSLW4WtbD324ZgwEYm9AnagyCPXAttPJtRTC1y6FE+Qze8ugsiWdoZ9fxRSIOo1riu/fbN9dk
KUSMxsihJDI76/9guY9Wti/JM8ai0iJc6fAfyFL+ml3JmpIqQdrDOJF5d43PEktuJgc8j5xriKSq
n5OYuDtmSb4DsvhA7aSOdtC9AmhWUGQ3+iuGwm54BBZJAi/X5sv1Kg0yV5eiAeOG4Cy2ii/asgGV
viXu9ZJzHHpvW4g3QZ8UliiwNevY8dCWVabBJaCCVE6TloG7UaZC2i5M8etIr4UbHibabRNLmNl9
l8zcAecd016xcEt3OpURtWCQJ0jrZfAN/M8uQrjUACfy23I2E4IQChV8sWF+Vzw+ADoZouKc1FWE
82eu1QAqsW+K2Q65AP4SECvWY/1w/kR9iwzNV643x6WV5yyO9+zeijezz1iQ4hHVGGSBahJzin/9
A0UVeplfbhJq/KgG3gX7Dn9ElGgSWEOZTi8MvZQCrnpJVdHV4RvpPNEgb6/hnm45OCoZWNBvkQ4X
yoHjJKiCxy58qhMgQ8qPT+DigT0/gt4v0QfBfKltQNOXEhuJygCIP1T0YQJW5F2DytDMMMvlSyWh
5ZTp7FVXXIkIupQe7uox8bx0zKRprvmRXonNr39Tsu43Fsph2VLHjtKlAUwpykpDyTRay9J7rLm5
XrZ16buUFA26nW6NE9xvRt4v1Mfd+AesC1kXqJVrOMgtQHQJ9yqpETSvfx/8Ml15aePJTOFHi2xq
uzSeSsMy45c4OFl0OpIrqlc9hA2iOHoWor+cg/xRMIy24yngYdpLVTDT1DHOUeHr7rEBZg5VDi/J
pHH8dcbvJiU67lR59RH4LbIV+jRipVUm0wEmj9APHjmc1wOjEBekDB/STtkTZH3nKPrB7Nh7nPS2
htOXipQMbz+zfnVzwzL9GXZCaeI+BqXkWrmOMP4Cd5RCTyMXE5w7u5IbQaZ5oCnhuUGGwiIWG+rn
QXCWcFLUpcNUQd/KSGhGo9WFOOxNh/twwbOwUSjRvDCygeb33U3G7MlXxg+IKpIqZZqYOiJu/LS8
rjchpES0QcEFge56+DwZKUzVLi9642pQPk9yDJL1OENJYkmMoAJNRYzuxN1wWUC/W677ApAKktzS
s185bUfmIehD5nW0aK09v+PQFqi/6jLUOkjhN0QCixmJi///Sl67zbJSPr1QFNViV3oqihATx65G
fx9BcZW0fkBcryg8PehmvbgzPCn4m/jLjCvBtzkrZ62u/EsegOZprmYU07xX8W5cWmW8cDL0iFGr
dp8SqKORn6bV7pDDh994iboKEyBKTutgGvtE+5SspOGSJtOdk2ni7o3dQqmkFOGT8WzsqvIyr2Ou
qPmY+vtVUP7/H8G06xxEPVdCH2d7n48w+KOo1SBgUvcEibks4FGGvlnSQtJrWm6QF1SLdzla9aoF
ycYdUz8l/2yXMb7mqUZ9k7uYIz3mfKLUc4/ELn11Tl1kgADeaza4wESAMm026J5ZZ+alUf9SNhoD
HT6eD4KXcVhKkQYWJG2ILfen47KYAe+kGMCr2KuIm39q0EeTVVTd8sAQG7D29C3Um5sb7bZmtqqF
rQY3y/mjIDBaNLYjo6kUBFZcJG5o8qphBsq5R8LgQ13vI2KESapYVzdqaY9tOkPu2Ky2reLZbg9U
eES9Djla9O36eA/ayPOt76QcMBRiDaTBzDQo8BaooN8phWqw7qXnXakHNyirmxODbSgDvzbdKwuy
FQDkYu6thECD4fEkPj1wxxxBvjrLNPpmMwahw8gIpBPVdtCZWTBUpLagyVyd0GnHXgbb/zIrAq1Y
s6MoQwhZJbIW4c3ldH0GyEBx7IeHRg/6x24QNoDRevlM2XicxwqxE7fCyYhk+7yBd7hpgJvOq2OU
57uZhF3g4Az3Qh+J0Xe3l96OuTX36kAxLjG41hmGpio4KfEjgHwaHol2F0E/DJYrLal6kQesC8JD
3LqY7QInzAU2D3VSv++BkXWpcci8xiZ36lil3cF3//yRJzptk4oFhdb7u5BKcFyvyUJFmmBBwqi7
/FclfYoyZwN8erG4/evNGrq7Zgz/ePTOhe7NGdqmJ1VlooFWHU9G11wkmeQ/9yOn4x45NL75LsSJ
oWd0DIBOz8zmGtJ69RR4xESgqOwJf5+DQGXs0syGr5BGvZ25Xv0y81faWWAJj0VgiM6o+iBbeUzP
Q4zyN/Y34t2i/bBB2ZqVWkgz3zQiGoC2Bzkihr1lT/PEJ5r1vCxqxP514UYPSLvfCpC3Y4hlzemG
LiiJaABEc8fRb1H6xdclzf5GtQyDibEOFCOodm/wipHGRP/8YMiOsMRDHKTJfar0GG8lWbeCY/uQ
BCEOQ2Xy9YyKcPEv1etJMf1PGPZ+8Hls1s+TRYcsnzoKSslB8/R9XLMaaUeCA+QtWnQGl8GfwOel
qhHonII3sgsF+OD144YLyDyLYKJ9hhnaNTujPRh57KP00K5OJ2SGYOkDjLgpCD60L9fLcDJqzwW6
hlouLpjc41Cmdr4hfi+fzbxR4CZfM4X4UwZnBU/Kha/u34SN7fpkJGATSreO4jmzIfPm+VUB8/x9
FgD35LUCGEE9fk5AHMRPmldPI31WF+HzvVFqi36h5yUIaCFodhgXJej9ZKpUnMQAZFZJe/dJVex9
KlTUksJMglM2xfPV8FAaFou+BSIMxXI4+ovxt9EokGkwxq5ky+9PZKQHvG8rnOOMN9eE2o6/+++9
1lIu9XKS8it99570Vi/OH9cndlNyyiDjO7kElQkyoYhzBm3J7tNJ8fh+9vgdHlLjhJqzKS8sZD2f
zVsDb0o08Bf4NyXQdrXvquujpx6yM93k/1t95Ddhg9mX+qnObw6JdpbLmuUYKKRoDG/IS9ucFmUB
bh+EIDjl2a6Q3X6ubZ5lm59HXXHERWihkEShQCH9H0RAhzVSRnYjRiRq7WnwaNx1Ak5MezaPUdyz
ODoN1BYEE+E+NKAijxGlBZmUoe4aja6Zt0PZsVNIPkzTL/Y2PDk4asfw02qjNSTyKVAP8PI3pDxH
lqhxWUiZ3F7JXqmcrNrxXSiFYQ+RYKustaT9FnnFa9/jA5J26zv6KT3nPJarJswFvMiFN8TV1wxI
302Czgw2u9aRKo0FPKQNxEbJNMgDzWtdLBTpQGPIKznPwSxuSyknIDfvtLABzAoFbjdwNImlrzLg
DzR3HBWndZ1ABQhtLaUT40XHBeKCVA02yj2NDdphSAKf7iKk39yf66HfL5BjeXqLIlsGlVUaVs/r
5tPoJsWyhytFnVQzj8AqK2b5WlO5NTgLVDqHvPoD5YJlRT4hwgtgkr3JfaG4XcDiERVxP0OTeyfO
lhB9caJjKVDW0yj8bdvUU58hGoAxi4ExpLRvfJ/TcF87vG4VlKvtP2g3BHTw0MVo9cO5hU5OBkbT
xJIbd77VJpubAvmOOyK/TKnOpJZB7TYUNCNcjN9ZjP6hYbDsUWJGZg2V2Q9JcL+S4YXoWy0d07U+
C7vU7eJvqOet/lpyA1o1rHZsXiAUT7iQwRmCmBZgHMIvjRYnbKolFxWwSL9knfs2AE0RWOsXm7D1
BSVtVfaj4ZuFpAg7zkyYqbxumKxAcT20EJ1VOyC3Fy9LTYtVJfvi6QxZ0KwV2zLqcO3uuH4s0hXM
cD5JOs2XakjuKjh7mVilbMEeN81v7+BP1Q7W4rtaokJ/UT/8Tu//JObvAVeVCWqCjXFb4LE7cPMZ
TpV9EZwZMN+1Cvq9VjCMFeio2CB4XUlbHAM5mhYUwoz4yKB5qJH37KaFSqldMvuJZsaxPE0E4zCq
37yot7S3Q9RF0t09XyHTnck3Edq7nlySjWoGRYG83lkVTaMjM5bdsqHw+lx9C5jrsVnVT04siqjf
IDEIiBHS8AESoJda+PYRTT1kFw30Tkz2lxlzOHrw35PK6GSj+Aa1b1YDGC1o/Ke23Z20hfQYkOvC
utdgrsRKwNbJO46HCjbtI1iV7fT4syxEHoZrQIM4FX+5vCGgAeor6ECjDpB0yn3hbAn+QQgvr8ok
DPFVEKZHau4mUQmtcs1PR/5SjBOeDO3u+/ktk9QKTLrgJhxPApRaggTxzRHxHFlT9bKqxKlbbWl6
0lYL+l0XVIHMTOLZIn/5v8KnZhkQXGO9qm8LqYqLVtgTbBD3WcULt+kE0FkzgIbBFjs1bWgHOaKP
IaY7i+Lb2+DHunf6zRmG9XCE9ZRpP7U21eIr5rSLW0UvoTpjkKOIgpmz8mhiTFDQrZ9U3o5d4Guu
E3c2EwVJyh6PTNOkqTLZGrNVV9Qpv8UVckWMKCqdKCfJynnQPf7h0TbDOgr9lmRfrDHzVHyftj36
T5Uqyds+MPWOSKDThPBuKDqpdv12o5HHVs2sLmB2Dfu3Pm8FFEMG00gvmGlRzEM0fKCyZWiz7cou
Ngj67J/gzq3xbgRqLHOXAzBLQAoEZXJ+CxtVg5znGHs9RJgVqxTlkUBHZ0k9m/ijcHgM3xIBKCUA
qjxudhAeN9hlHJFnR86fdZhAz8o6RYWs44a3LxYUjSGDqxRIs0MBHVMVxYMiDO7mMu0Buw7HTvzL
vykOSSBVmadEFtebldKu4cMsiySSwtiS15d9Oib8ENLI8lYzucVfrY3Ne0VwyijuxoC/XNDHVp1H
NSNdhrmdE8umnABmUz08Z2idE8KggUzTLN+aidZV/1USIMRyPzbI9vFV5OEUaj0dQJrYvHpK+A2E
c2O8DFH06ZKP5yxhHL5cxNLSN8iVNhVfvTRfxzsdlQZ9RDLUINX3SIdMoO2vtmNW4IvD7M9UBM5M
nBazYkvu+T7QNhgC9e1JnXRDztVWvRLH6hWx+kOsfO9RVVxYMEgg1IQAoLvFlC0GjQFysavY5ngG
HYPFs93RfdVazhgtx0OP1l2U+pylv5OjFk93NrlKuZg4wOtbSzxioRFM7FXdXWagrPUUoMcWHVdu
DyhUWad3BI1hJlfgL/cKSIynjLYQZQvxi6U8J+pULmfycIYvgyeeHlk4dLUeoEwzdEFp1T/Gd/un
m733h6/wvQXFs1PLBpuD4PB/Ut+e4kjfY3qz4uwR80JlEGjnG4byFnsYnz7u+XG/Tif/dAWt2Twi
Ccl0mg5K/AGOolHFC0PxgoZBG4Eew+npCBqYmnYvZ6jbCJHM9liDHrIKN0yx+4Ma+ubZkuqaQy1e
nRZenPAloldKiZZKE8zADOIUjfbfvIfghT5rfTGchCNZInjhpgK3bwLphit0sIU6fScEwrzWHp68
xiASiM7uCkWgzzzSKlZqKHmwXHqmZnrJvp+V1LzOvlziI5g+uDLyWkagZ2a9HjchYWnaykU3i0ag
uani/e7j2XA2OBdkV26tnA5EKzjKBGSD48rPZ64MDDBLY01ATl9S/a+x09j/QSyy0QZm5Artvb1V
nCvo5gnQK6M1KMfK8NJ0Lc1A5OGEdjCsf0+Pzx9HuGu6RjeaKqWsC9qA0VF6Aws066yGgcbPI0In
mTK3VF+N+xw0z1KErKuDlKIMy11jPb/jt/vcSSX6TIkVs9Vi292CQtbhT02KJLD9fAcFRvVbE/Xx
Mk94Rdmq2TNTdjrtdpu69LFPeyAXdPWZXPNB3Qt5kYFlY9Tz5af6GtrT/vI/lxyi/WycNaaI78UN
dD7u8rFqn7T48xMSU8NF8ebHqE6LKtLPy0Dfwo1b8DkDNTq+9F6A/wVndesPJqn0nKbqZFv4FpWU
JDSqARbIN8wmU0niCQLDTZY8zs9CJ1VzX+KPZehn77iXOjTr1hDmA9aZTyjOCEtdJkxV1mEdb/kT
vVTr6keAFoDBLvXdYr1VmSdjBY/DNYfRZqqt59D15RXouiLrXkXHZ9XEyCnlbLW/z7uKS5Ztk3HP
UEGJUjK8X8Zxp54jCo0SznFanSZqAxx9tjxPDgOIJAFQqJMY/Ry6Falgb5y/T32UGg13Bm0LReyh
eIFwHOsN3Og3OMkRwiqiRnHyW8wb+nRkA7/BlwojUc8ssNWqsTlc8hPWv0I7HAjMWPrt0HJpBD50
Lot0T5HJDYRZp15iJ2gRne7vlPceXJq0qlduNJjSUH1YXbsuE4rXmPG4D03adbBO3WTvdXBHMH1Z
r/I7K7EtuPXgUELxkfxoCk9eI+c+Z7dyxAlNHo/azlh/sze8cElGv2/51qhUshl6zKgLlMtd9kCo
HYeWCC0RThJ/UBBPxKM6ar3BDJXWbZ51kXi4l1GejX4p26I2fuEQEyECwAsPHmeZNtGl+OX4bVu+
diRyB5CXjEvBRS8J1knQVvex2DRYVoBV2EyO2Dcvbh5rH8TCyTYYqrHbRf1e9jLwDoQDyPfDqy7m
yT+lmycSJBTQ0wBXeiKq6C+u1oV7ujWFUb7j8pEeEmhm8JPqhbbkDMk2NyteNb2ebzNCAZYh8caL
fEy2kY+HmjMwaNPGqZcrss9mjl472831QbADFwFM2gV+iUM9ti0vzV6FrjLK6WF/X+89z1d4v4lI
TALsI7jRsuN6aM0YuNrQsFHDT8CP2D8nVFldE6t59wzympO6hvM+O8guQhbFq/vWmhHyPJTH9V4d
vUpkVwLgv//UH+LCR5+NqFpcBJ/1h7DFAt6ulGiMJQ20WI07JxCDfjlrmBClveklJ7Syv1R410gt
wOVU8EmWR/8FoTaWiFrD4LSwla+ileDydc/ySAmTFHyQAIY/Ax1RCGvrGqAMvOgtQbLfrT7xgWlK
rBRbVP7IhvKezsUIhDQ8rf1vJjNJPNuK2pF+5FWo5FLlTHoJT162wwZAZ2+2KBsPZfpOol+Fhkas
JB5Wlk+YdwmLfozozWSlXGVqoxz7oCEOiBSk5U2FVjxBqSHKyLaWI5OR7FATpjFIC1Cb2XhwrrGM
1XkwwJ7am61elI7wxJphXv53P5DXoajmcR29OWGPjNk2NN6VldqPzCNB3b1ST1EBC1pYKFIfcz4S
PT5sEzy+b7FFOXBdLIQDpeUFxctyXfe6XGtGxhWX5LOExB8LLK+uSQlg0L2nBozuajsKGEreBfxD
D2n390T/YXkrFa6SwTa/KTdEPnB9t4Zj2SYuTwvNw3Wse255Wz3TCRBoo29oHYBQnlPbWE3fRnZ6
bVYe2zg06y1XcUp7A5jj7cPYj7xsXkNvKpOVYVb1KK4/TOZUzWmddIPo7XfWfh/7nxQKG23aGhKl
DNLivUTj4h/z4PN5zlFEyhTCY+FNwX9XB3oNkHu3Gu35/7gfJxssR7mjtYUAuWkT7DYk40/TdXMa
y09ErsFNw39ayewDH2gobGZLP9yUkhbHuicx07MD+mNcAaJqfmwnvdkv07hOFeaCng8GuDGjfYXd
US0IBssHNaXwI9ZUqM7D1k36V4NXRqn8Ukcb1jK9XKnlIQJbYFRtlW6rY+7MKR82OKOut4lW1E9S
TW+YdWkwc0Y4fPnGeM6gLbVEYtGUTAy1EIiMx/mzzkUVGIkeIYJWGyyek/S9/W7HcT+1iia9ysu2
reTMF7F7T/AeP8dausw48P5ZUbgWMEu0OjeV3ntt72P10wbyGYbeDhwfMzPmQswZHnTZTch1+058
7BLBh18mcTQPywrFkU7Wv2le750f1REA/9Wm0rUuT0VizjYdptdwMXjDwumJnZxR0ntb0AQho2LO
avZhTMFqiKQujzAIlK6HjsmR6Apaw7R8jy0QZ64ZDJHQyTwb3yCkCnxBACOkOekjvkKV2HtK2522
9jB2bfRxNrSA1i/jOf5e2X5AFGaBeJ26+O5XnD28b3gC1xUSccdbf8Lo1xn9K+kOwyPjFbjCwnbK
HhVWFW3r4NgZYD5R8DDFdXX5dNeekZ96Bn8wYYRX8hc4gd3nHeQohAYZ/a1oV4sLY+h/2Kukp+u4
n3+Jgw0Q9Oc9KyW1ZAqINL/AOOrY/uAD3LjFXahYGUdJx2oaSSZYtDEKpwyZjEQ9/BDGykr0jUQf
38A5g5oMBEsdjlpd8RRxk+yE+TkdP7c5zGI4xOqB4Mrsj65BRpbqH7n2dQWe26XIPWmdx6snrD0U
fqoKrnpXNZKAAS9DD3CU6ONDScGF4qxOLIx9GnKkJXSMkmDtD7rXC4TBCvVWNxehgWnZqjaSyE2u
PbuUGMqMWJaZQhbfVlywkegEELHEKqjLpbyKzjgwFPKbRXNSvE9WG9hP4VleAbtFfc7JI7me0c+I
7j6ioampBBMhHgzXzbQ5PVpx2oL5KDxdE0SzN5GkCbNR/VT6D0qkUEMQzsu7g2pvD/cPS1yDkrFX
7ER0nsQ7ih1qlZ+1OjrhmyfoR2BQTlT/IJVIRTkIznhkBD6gvpGNIC5voySHlFnqpT4luY4K2dkh
XxgBLiBHua5Lu3HN0d7bBJNW4yvzKwnOKdzCvLdSH81PVkCh+N0ZNd6hZ4hBK10AgcD5hICBvy3X
dVcELnHhXz4TrbiuYzbf6dK5IkvSGAlS+e7P/jVIXiWZof4+GgJnJk7WVLyO9B1ocxf5H+WgWYN9
3Fdpv9ltDVRi6vBiaVFgIm6mpchsm81oJfi7b5/fsPhF0yPFNlkwMVPgNgAYvMqJvnRAE+kCHduE
4E/Amw2DFGMAuGUFBkNu7jIQ/hFgJTLKdNQSZ00jojwANTRnVcZcIQIIBbO8LeA92oepFZJ9q1Tp
gH8BMHSH/4a3zoz0/I/0qTOpOc7efvpFUFiJN6mw0jCxRuGmdqmBV+YgWIN5kt4nyi7kSNzJRZtO
/QqALfwhl41dVKos+FNWw0ef6nPlyhCSqaMuMLQlzxXp8IG4hp/cRTTrifVnb2OgOMryf6dzY8rl
wVAVF5wAVupzEGT3rEw1jRyZUKGkjtu0LHjHI+rCM1rg6dBOVE/gnu/o6bIGV8MCf6jO3Ku7yIiV
VCa9JFoaH8O+NlqNY8WyTU3tjdqzTPx9B+B3vynr+uQTmcet5xS2tOnYD0SLqEt0lPBMAKKOYWB0
aEhuhbfGZ0Pn3LsiUJZkTv0LOTCCywO4tqpt0KQlg2dT4HQV1VJjR/gexB+rtn2O7wTep+GARyvW
JQdIsUMpwdAL0YoiDkfap7g71UAQTGtmws2HTRrE1sv0gd90bhTJPj8Vy40mQJofgkOTv5Staxbk
1SauxRQtqJCj7rjBWIof5LDN/tFveHsuUVuNjQETzmkOyGyxYY2iDQDRj9oWnnZjL9vNYTMXjEvy
g0nUx2YSk+Z7KS1lWCQ96//W7K/na0w74dHtkcQR1wY1URE3XrG/oF74pgYpwyn/RwNg0k1++c38
8oaNaU7zwPnrzA4C85adWDjKD+1Skj1kRH3MFi2Vlfxtl5Dw/DzJxut8TKkFAsnbjRE9k9nMxtrF
NOEB8LJEN3V7Qzbrumu/LYEz6WJ5RuuyX6Zzbk2sKkee8JZmUyBlwlDAEKKzhtuj8JeyMwj+6xKP
T4XdCT6UmuwFwVN8wnF6S2hWHaJI7/mjs8+wFmkxWISY3te5z/tt/jwAT5RymZErLA8lc6zURQpQ
gBVvan2gAWyBvYvAXJO1BgZ/yv68gTvBdrUsJz6dtRK9+FBqhNcW0snLQjV1AH5f9r+Eay2Bh0TZ
6M59PfcQ1Qvreex5+FEG996n4VXhVQKRKTebHRK5eHDhkJzBnxOjC3pERVM/KHdMmUsL4tbUMJqP
VQbtZ7yDhqwTmnJa5DGhHof5XJ2kF1OwR+68guOUvPAG5ERGiT4qdSpaCJ5p5wVCKkMSK0cB4M0K
XQRoapGXEhGAHihdvuGKZ0MFFGbMdRxCzm+wuZ/rNeQPbrgwYzj2bEHor71g8KsFP7wZRo4tErtz
YZf3FRScSrOXTf8fJ5kuYM6c9OKAjDyYozS0r6B13OSMLyB9B/cBQNlCPRnbPB4Cw/y/EiNqcSUv
CUVrInGeuf/IxaGEUeBRGjWLCG3sAskf1g1NyMtFEcjr/Hm29xE+z8OPbpgjXIkRhBlVQ2cBHX/d
hqv0k1/hun4tZe+pv+T43onmSsLdxvzdyHjPBGFPlwQr8LvgeGxSjmMk7BR5308nJc6G1YO0iXrG
zh88nJlVOJrK2BgMxDcqOQYOzPHnRFcsk2GhHYCBMb6IFq4K960cAepXmM7idWSdnh75X6gFzP63
EFhXngtHJnIJqMUPss2TPUxE9OmPBnhT1WmW4bA+fRaTnBxGja/srcQQHuGj8NQmobVjKssUrI+f
H95Cq1YMAAoGjD8FxLI/s/E1OqmvFvZk9QJPI7rTFpi5iRCl28b9e1draZ/C70gggumb/1m63SNd
0+dpCamKc7uogHQzH9c6cJ/p8GvXUoLCj5qVrXQvBbuQziMBL7Jq/fvOaW3BjAnFrfvlVA3dMdJE
8kby9aMnkpO6W+B9ddfCzCOZFInYv50Iv/3DbjQzCfSYhjpeJQEgP4OpnHWG/m1c9Fgz//z+LO6+
jkm4n8w+JN8ePdleKu+IfadYz7E0zA9AhkbNsEB1Sv5PivtPcoOvKmrDgWCs3by9LRapB+mCX9gK
5YA4gARvfLgyWdF48LVKs0HJuIuiOLpqcWuQurmXdEfocifqsICpp/cDKmhxGDjW033xyEm7aZk6
jC9j9R8pOFsFruAgPSrRA9mxMnr8jb7zMKa3eFDg62YyACNrVTpEO3XQr1ehqVFKilua3w9TAAzb
QIOc00aCAcHXsruwnBMckztjEw4pnj97tyimSqd/49MwyFUqpyiYCgUjrdoCJe67pl7DjSYwIubk
iK2Y9cmhqVYeeW7fiwtKiA/47KDBPEmoAtJ1vd+7cUwyqcC433qoXwxxaa5yGoiPLAn6pOooMJqE
UWTBiYMMmbS0jVIyOLshbBaVCE89wGW9eao/c2m4gXGDQC1qem3epMsUCbbHJFRwKX9jMbWTr+kg
liYw8Fa1ZDbEyl77iW613fVL/+X8Vgu78tzJfHD8119eD9wjiMmvEsEHNJIhXy+g1kFp6LpnCJAE
4/Fx2inFCPIk/CAHbpa//mub3KHVJ6ogQDDD9NxrBwxSRUtVzOe4t5bckwP6iZx5f55Gk3RqBpxo
FQK4lX1uVkqZM+0f2y68PSh/4dl5HOzu4LfFzU/GYktRBVQ770ji+/WUEXupe6SglNW8vK0bY9qc
bHDRgLa+qjQXPjN+9G8y3PqCxxRue8oqk0xw6WSjc/rKH+KZF11rHQQmxqVtO1p6iDMZ+COlci23
slgmQf9Qi1FdNIg0PoBzGVKsCRbzOhsF+qqRTZ/wNP35ARLtrJbFmfCUAE6VAB/WbVYY/40HTSZr
5ozCLg0bKxJxbpEXfGQ7KK7wAhktJKIPtHuS+fmDSFoJyB+TjHmp5oXwBG6/MunE84OZ8EkACbA3
51YJVCfzbDXFMi4Yl5PMV1cNwlW7z28m+eiKqufy0Rx2DETZlqLjnIlXbqzWTJ4kFUIYGgS+3rL8
UC1XP2+9uMRGpewoYFo3XVrhmzsVbLqvFz4rUsPrQTs3Oy9oYEl7jiWncrpw0AhypvnqUeJxWgOZ
rpvACf3Zs5FzpfDXM0Txpq9i3wfCfIznxezNXOM0Sqc7Y9QbKrXODOJCXMVuQ3iy7Y5lz4fyhvRt
BM657DILyzA3JKNr8SXVsTaJemvqxJoQttaXqSvytaADN0Wjq9tMEJTEQm1ldCrMnS+TbHBVlZMS
jr6H1VU2GwQ1aVRUQORFxMpauwIvt8S0nnLtIHVbgICOeAdbjv4ul1Y+RJC0Dqp0UdnDy8ZFN8ak
8RVxqtVkgsGC2Ks3sXfyVXvd5bB+muYFuOHZtJDso3KAf5qLjtc5eegfHhCJL2immlm37OLmES2c
ohLmHgvV04hY3qtMhir40BmLBGdDL3Gb4u6UhB5lGL8c/XVmIL/Jc+fYR1bgtl3CsDBWauYI9uP1
Uez0nj0dnptKb8rVPovIP6M4uQ7cpPL73BZpYSPnehoKdAnMFvf0VfCLLOMDUvuxVuyBfDRuhBOr
DNc4n968QUoBwzDevmwYWRa7Ri2jHHKSsdYO0gdAviyn5hwW9fP++IXbJsjYmdwaUgRfZNpqpKQ2
3L8CPVNxk/WZTWBMI2Oag8rYK6IKyBrJl6PPPtc7qWAbBfD1M43CW3GKwFbDBX9s3IKlB87qrZZ8
KwnXarwYPJkROAcPepNWcfAQmA+PuoxdhcfIn9n2SFT3FTkgMtUIiJTOyUTVSMqjg1hsAQ9f9zdD
DvSsMDKZIRH5wIKkImNptvyG0y0sw2Rcd6tQMtuRikjND0W4UXn7MMLIqVKzjlR+WP9VTWaFeJEh
VJ5nwPwSWoGY7c3EyPDTFG77enf2GCLrycSKboMrLyMC9jLeLf3BNkSC+bUpvG9/pYop9BKQVlwZ
asyblbkSs+3lrh2HAJoBXeLeZhngxkPftxF/zQ56F682wtmgBQiCcN9nDj+DkxC2pqJd8n2LX7X1
vSRInXfu/d8wC+5I60fWQYzNNmGS4fW2mq6up4K4lvnWq5+P0TShLp/HM7uxa2ht9CpZNXRZgJws
9D3+fe5+zhMKY/mQpeRJ7XtsyStBjXG74AfuaGB0kqlYIZR43LIUbXS76YNMW74jGdrBlCnhVKQq
/aReu0rGuSRwEEXeFlIhBgqRvo/G6AKHSX3VNqIWJX7IvX88a2TfVtjrI4pd3Fpf61HFsQJRAQQI
Xvgu7+9hsz86LNPbXnnUge1iNRSxAXRHz3Zh2Z1EJuxOx3ppHeo1fqGbe27jV8Z0pE7WL5FPuYMx
HpgbUr4+vkAnhheKWGCbaJ/OIPIIrDCVnV0E0ZjBKZwupj6od6ZU+Ebpddf6eYYiWWfnHlFM+Qve
SH2/iyHWkC8Jq8qMinNc5c7LJF+a842ctiWAkeyDN1cnec3Ea6lz/Vvbou+G9aI5xr754m1oQTMf
jnehOgXLena1eQfyWiL98d5TbRseV+PULOO7qshq58glHgYPthOZ16bbNnYQA5LYutrPfvGQWJSX
19jTLxGg5dmTKE9ca6/NoumTOkWet7vEYSM0vW/YuQ1Yx4/BvaNurV9d5k7be1u+qhqLrJ6zaQx7
J9if5cLrnJlA3vCPpMB51otIj2Z0EjLD8TKKF+ebYcioPMiKR8iU1s6Bbp+wsu1tW45nAABFn1eR
rSw1h7mJvd67t8dEksUCtgZrZaZKgl9y+J2rP45EtELkjSaNDev+wvJvCW48PPiG1qzTgdx6Ojgf
vv1bOwH+8icSQ51SWSka8xC2OEd6Cvz5EDKZ1iMpn1o8mYQxCCqVV7h/lXxeZlb23Hn7zthpkCkM
vVQdh68yKveyXnc/3nRM57HSyS1EnWpzECcWGKGC0K1ZId6XpJ52XdrwsUa3oIa6pWYLVQcOh2zz
ifg/HwP++rn8f4aGVYSgjEZtvb+5fezSbqzWF93mlHNkY9nM7mPeTUT8GNlzOLRRk+DKtjvC25LK
+qwlnpphDZg9zfUziUMmRQQLB/JA1G4gFbNXBloBio6IF5hxct7P7RIYVhchqE/pSKIZ2yU2F/LX
GMdSKDXkVSQmnQwaS8KIw1m5WJyQ1NTfKQWnefIWwAcKtqu+gRnd8B1VsMmaIHITqVD3ngzhISIK
kyS0iHqDwAJfXT1t97ZnhAYZ82RvQ3u/D1VRGciOLuD9L0yL/POZ2lh8VPhhS8SASzuK9IejMo5Z
RT6Z8lr44NmKqO3QsiUQQ5bpRxUH0vUUXx6EX4wUUZeeBjkajcSsG5qfuZn8ItMYdsM44Mw2U/is
X5T4XjSNJTYrQxFKReV8xLIkCb2w7ef/czrlfZTlFW6bFCeehG8pPDcdXq69IKi6UQEEXvHTq1Sc
5h4MCOArp38OfDnh81sjJW7UvBJCmxiNGYwksGfBzo22bCzBiSYIrMK9f8pnf62+zpUpzYMNQXB7
zihqVkvesPqQiKj62CfE45BjWtmNzeP3m64hyByg9OQCebq9RpP75LP4nLCLzNYpbblUFdUW0RRL
6LbS57e90ktwS7zVBe0jPMzJZdO9FCz6SE0/h4vNPFmVBpQuiNh5UGuPag3OEyBFZ7xwixTBWiHr
Js5lMyoXVVHfBv+frhG7AEXSouHvUdEexSUHlwgTb/LQPsVoySMMvJtJ53CvvG6D6WjqOtS2Q9Gi
2GQ/DBPGboXPxYlcLbbyKgjOv3yWYVjJlvA/NGv3TSW0w7pH7UEFvXyQy67fTIB/pGWMM7+/njoB
XucyKqGiUctacprbpTMTxxIuShfWmS28Fx4DW/8PewCiDZG8pvJ3x/xVOsbvWRav089kQ/PIh46W
jydTJ5aK4n9+Tbo3K1QpmGMAhgKwwbiAaeaaA57ZXk4VVeBW1DW2wZS/GZjI3LDp6BS5G5+lqQ5w
fwDrvBPzPS+ZhHUwWnNMsKHXeCCtEHW1G7Y8UBHml6//19A9KqyVGWU8iZWytExSjGiI2t58YidX
IgW+KXoleyHvonYydyFqT1faCsBqY9YF3AbkgJAQ4FEC70C5bH5FteCIybxVeIiDxukuQpvM+dkI
v6xEt02q9xDBr0au/bGtyNaeCmXbwV2rqKOXVaeTidOCPklka8UGtZfLJ9/Q40VITeJjufRoqynq
maeKgFBb4BpyqYU6UME2uH+6XTjWvoNK1oyMza2S4aZr71QpI9mWsBvKxL64qSHzooRe1+Y76YgE
8aWcshsieWoHjwdrwXNgh5XBX2SHcMLvsWav5XuudwQL7GPSs2sPGHALqijlbAH2n69SzNNANPu/
WAaevdlWc2Af2c7dhfPBO1fTiBQrDSXpsj2HJXOYM41ifQf3MWv9/9po3zo2Xml6+YF5sUVh/jnR
tZMX2GkWP8TPez+F3Qw5R7oHUnfR9PchxYkYKQ3pYdQTq8Ktvr+YE8mET1Id//HKM3KUtTEtY1F9
K0gIYSBHtreRIXHfKIPBm3WhRrSz5YS3TwlLVIJE3n2vg7crcanyZq2nHR9HRmQ6ekQNPhZb+59v
lU6K97ZJMCQ1M1oVvR3o68IusaK0ZFNQUcrDF9ACZYBkJ3T0ZcfKPYihpXbES9r+HbUZGgVVbcj7
D7K0P18/CePQ+zqaB6kDU6PPXUcj9j4IkO6/Apcfy0ZoQAY8UccA8lpESs00M7ZL1QLyA/0f5NjU
WBnBAk8ALaniboRTWtt06C8D8iLaueimp8v4e7s05L3fjrLlMoAzUW9v/mtSYUnZEokb2sjY5yaK
2uPPjVVz8Qnqje0qILKU54wfD+aa3aitIvxvntGgAtkcYSHl4/8xuzYCkjIc6pcGBlYHVL8xkpzI
YJR7KuH8T3sFlU5JBt4rQ5pP+kJjISN4ieYxob+b1u6cYz/5Ag+GdhHLi7diq0Z9bmyw/6LYYH1f
WlBvjUp/wJMetGGEC0iJDOvKoR4Vgo1kEXaLLG0d+wodgoaHM3pjG3M0UbUS7tDqy8ZbqPV+amY2
x82RPb65doYSwbOybR0yWeCUspCQKoPsciZZydJvlwe+h2vtgu1dZysX9eCsKuh+A39qRYvBapa2
58UtSDARCrjOhDLQXR+qko49+2Zgi7jPnqRizUru8HMVv5FSDaqQm5SaKdH7wXL2hbj9HAnL38UK
dCSR+/sFw8KGehPVvmqrEb5YSfzFwyoMIJwJYFnM9+2uBuYmL+0x8FNcBLEtDFMu42tfmQPyRj+r
PQKMtkkRxlwoSK0OW5f2XpTD8mC6vbohmoXGuroQ8gBcIRCDrrIG+8lBlEXN6rNRhAnEZYhh3t3F
24IA9UcDS5sxKICaG+NsBYtmVt51PjxKeO8+nfL+FJyxZen8UiEF6GZLCGMNtuZCcAwwxFPPd7Bq
+y6eXSG8BC1PEsCFvkK3ch3haKA6esXroOw5TgJ5b4YJUlXAPFVr5SSLLEiWBAJPqSPyX+nA1V4w
0quoCju52bisTWd1m20nJQXzZE6Ojl162Z+0+nIU1KQCgORCDm23RNYqoC3b5HjSuTVAFE9bAyPl
5Ty90jN/XCH7QiFb3tcLLDrsSm5uFcpfXG42n2i5Vp4ye8hko5g4jAEeF/QKpcV7aOXbcpbsX1my
f6Oe7kD3ganU+WeB4OzuqZQju/5FEM+YVjEde1Tc7+bcpuJucs33ClYJs+UyXRGvHoI/Ro4JyJtM
j5VJTOKUDh+AqCaHiFD/GPtqhBQhlUldMViCF/1L95WAH9KdHxVX0oPtGCQ8WBhmlvYODMJeL1JT
gLtb6R341LSptduWjcqthEPPPACck8T2+aQwFpVO0xvs4uegOFJVpZBPmK/YoO2RlUf5m1s3LI1X
QoG4FOXuPk1lz/f8Ont8LAVBl+c1RdYPXCYwyMWrLoB1uz4hvPurNs+NzAI7oB9ShzQPEUxUvlhS
6MdAYBsIzv1x32zvCyezcuSDgYplV9iWlC1UnZwuJwR7DzWggrDIp/5CXfmeroAqkGJSssA+55bn
z29xtVkvBUkTZh3fEuVaqCDLczywyy3tRpU3/GBDOL2SsOHxPVIYU6bfDVOwI2IypVuH6ezwvgh4
6u7bNS/4/77xZ8LB/tn73H7tQ2leE4AUsLYvlJIi7qkXEqfd3wkkRJrsqqGPtdkCrgzGWw0UPRcU
Hlbw3csbpCood7EQFXBnuNllCNWhqjvIegd930IxiYouzD+Z9+cu2poDAR2KPBY85egFviy1Ms1F
RZUUBWnUARu6cjfc7bYGgckViWG9iJJl7p4wQQ7xyOBtwbDyzXeeOOL1izzFTytYW4ydo67ks8OL
5KoxZMfJmdlunra7LfHtzoionXP1zEVd8TldFvevF4Bc+MqR7FyZzRQgfwaQxm+7gjBZ+dW3jz/+
Ntve580YZRMujEb4xK4J0OvWpOuuYQeRCMdT0kmeTfbvNdhQlWn9ap356mvs35jwGnBqmD2mb25K
H9HyJrNjJ7ME2BwaKLnl3Q/qhrZ+std8NAgOIxBrvs/tBE3E1+W6f4bJU85yYz0UjliRW8dL9oWn
TVb6N27tjluYp4QKrAzVsgfoTxuKtNwU1SUp43eZ0N78DqpT/9t9edMviKOKHTvE/au/TixucAyK
dwla1xOGjPTIimnalmyg6i1ykkMvUklvZIXawINxrYaR+bPY8boaLz9t7YWuNzbObvaNeAqS8myK
puKBBopoQsCLjJPU6RlEdRZIBK4I6Pw0vBfQiJYyCHKVHhG/pUZLQfSHIdxDN+xN8vuLNvViOLWZ
naQcjXSOMHQL/sQ9pCQCdmZ9CKlXbvMh0QD2zt8MNf4CoWInharcGi/VZoXySDyWW0xc9y85dVwF
5PCa/nJuLscb34W4h5gEfcNUppQ1JdF0czln8LJAFhthLeI86BiOAUcFdEB/6EtkN7VoywRBVTUe
aA+LkpRghzDhCQLdjA33V4V7x8N32542EATWWLZcw4DtPYqkCsrp8Q/21fO6t+XyDKvWNIOl64qa
DWnMt3uT0y5ppeVoRLhvtafY1CXglSmFUlrqD9DFC0ZKYKYkdw/tB1fV6EI3M/KkkWu8s+R63OLt
/t79ZXp2qSGS8iGfJDDuwCIjlwLfaRq/9WF//5viX4J+7gs5B260k27JPYd8NcHmKyehXI0evvPC
S9MxH5EFSKp+hA0qHVj/AA4p2z2NsqLRstA1yyvCExx17K475GJspMpmYsblRYiwnFAx4JJntMZn
oWJE2Z/p7StL/pHyctnkBbfeT0gB9bQRaFMPz6aBCwkOh4qZiUN38wsH/kCl3Z+NP6YKjqkzq2hD
jrEy7EWhyqqRB5xju9KyKpzGoPwemH3+/E8UOsrixs9Ct3j6nKawDnRB+tax+Fxtm8HStZdmEJnU
cc5e0KPa3eDeRprqqKbb5Vlj4bIFf+UTXKQePpe2QuAUgPHM2ix4DX9S1uLUb1U2e70mon4CRLMI
0K5BrLT9H9EeGyc4PRVlzVj9H8eKH9ozXu6lGtgd7ezNUXRNrJFpI6/cnC906tcAKdKPXLuXUgdz
UKyldfWGrVy4IwXn0aOhwD664/HELc7Kq44BPBstWnnN0CHqiiscBTI81XQjrC1BTwC77L6iGIlo
+bE3giMdP9fTAqEzq+Rt7Uj3IybMc78b15axHCXUJ83M9Xb3yaElEJKK7Y/jrD6O2pj77bSYdYai
Iq2sVULdxKGwPeco/QFSGlqvkBaH/vP44cmCHTGplnIraIRQa6TtujOee/+rRxIcX15CMiTbied9
kc0r/GsBoo+cYWDoYoTlH1QDba9KuA5HG7rbhBcBVXOok+K+zlOTnm4WgsjKgQ8OK3QxkJ+YKvlu
C9lLjhhXoxpRUpmholz2crN5R7mA9ONN7SElDOWobB0kXHmXv5uEzQ72Wh23xHMe//wr3bPO20oA
KpLIUiMSaUpvuTLF9ZzzCz+yuIe+/KdwiAS7etabuJMMIBEl/Xdlh2VJPsremLgEQiCSjt6lxRqI
/X6/Cwhn9w/kzLJS/kcXCxYeH0EJDeF9//eJsG0VEyQlRu2760ZrRNw2d6Hxk9Tyu29vG8vcIpdQ
lVD7KT1EvqSs/YMjbqHNaDh34ipACGxYzg4UHeQxegEvhFIaayAUaVq2TZuUxouUdIBQE3cRECxD
79VC85GtjpQDhFdSXQxZC5PZKPxbjcJJ7FMMuKPAhM/vc5MiP9nYiKyBJt9rIYuc3NrgZDE2wlRW
rDWeJlVrVILhs8Rk4LfmSm2t8PR9VSpITkMIW8v8qayvcF95369LlrVnTRN3qO8wDSxq4vstGxE/
4a+OLCGcySWutxhtfXqju8p5pWkc/uUsLNGXw9D9DL6dbhgDGGwhSVtOBzA04rxlmht5VddtDDnG
+hRvXmTyv5NRay6J97Xd6kH75hE4wG6c78tqXlJR5dntKaQnGLahEtndNX11bVqv78VlM6T/R1WY
lNJqXI1kuoJyW54eHma454IJGZQNC9mXTyC3rBJKXoLYNzN2GYVrDwYuiSye7uo1wa4xRVkLV2W+
PcPKryV0B+fEz4V4AgL+r5ZvUtHABAtvOQIeK9HDKbIn4M9fOK4ZgREhixu+G/s7qCUuUSLykvqZ
RsaXwygJGmBgsW7dhrSPmaKUJH8GWmkA8Mbm7batuoJQ6EYcJO5NqYpoIHcWtBn0oCxHS4BlMSkI
ojJy2wQh1AsT6cw13HGvsi5R82V9hj9IoA9AiaKvowOX9z2fvpv1KVtWjSDRQ8eWV1r9dBIPZFtG
4IGvgnVC+fd1a3Ke8lEOR/I9sMThm63R4Wr9ihj6d8/wgBPo8JdSwBGih5PFZPnFBxUgvkr/OdWK
CzTGOkQLEFwdK7dGWwFlPxSFX2sT2Qf03jIbLS0MmNDOZD+dw3+9ktb7NvmNNvQNb0snsP+ZYiDk
NsaOAXQdQhmyV8NovW28ixAyRf1pZt7yxFm9bxWgDAZ+8ZXWQ/i9IxMt40i+Elv4Ofpx8ZsbunPC
zvU5XKSf2NaXC9cMK+qW1gCx8l+KdY1Oefw7Ptz1UI+i54/Wk6OgkNsGQQymI+2VjiiiHGMbShvS
1JWs+wERrS8v+S9aHNfAXrxiFBiiYvfxQ5bwQz+1KyWByqT77k8Y9hqz1IDsljkJaxmMN7l4f0ly
EorhPb54ZWvkJ9IJRJ+9hmWqDDEbEye/E1FYw39gVl2w4iJov2BwVowtI1AWGJwZX+ya5X+rDCIa
axOn84y8+NiZduGshkucqoWma6+9fEe5H1aioO71rdAK2KKUjOzI/+srACmI8t3fTwgC8mSCpbzR
yK7HH/VhloI//qoUETH5Dg134mSkl8xCUb5DOjf4yg9WPS6N+kWWPKt0O9DEA9EDpo4Mha/z7e8U
dePnrAzi9MtDJO1a4SteUR26RP27eoHHqKftn2GDXazjPI7lBEYmEAuelrnI5W+4JgiFK+Q2GD2W
ZHsp1ajx3QnsXzVHS4952wncQyXwgduz4m/xd70cEf/yhuD152P/0rfCj3NvBnsjsK5dv63KNG7G
0LvfrZ1UkYstNwQCcLr3+zeZcfmO5Jjj1tUOheTCd4MNMRLIuICSwQ0Nf4ySIe4fuklqPTgZetZw
WFVAygjxQo/uhSSt9FYiFsNJ1msvg/jcP/n0UOcV13VC4GV/bkih7Xiwa3iJWCMItgpeSiSwWzO/
oee+fAEERZRduV+cidl4FzJ2bj/2uyQZ98kTKfSq/JpiAs670PIzbwo0JTPEA4Ya701OON+Bz91V
RL5EfM4gsOuRTVLieXgLmJnyQ0mCAYVWWTOHeihdfrltgDpWyyU84fglw76SLT/SUfG6E0o1rwMq
cNv1Fald//axMeYECiY2/0GdtRRPZ2LZfKepQs7Tcvb3XwiulAtmo8lWhQjhKxIJfvy2F3hLVvoe
FKxoCAGu91TZA8/tBj6c15VJ+cQ0yyNt1ay0XgHKDvos4UYGSYrdA5GCK5Pn2/IvkCe1SUgFu76b
Ec9rkEMvCcUeKQb3w10/s43X8CnQ5j5IUTrUY888AjiJrG/ArXcDlQ5HHTa18m2KOGtt3EDACIAi
WQEzUpP5AGDdvEgZgW955m5z+Bow/J8uFccqUbCxWoxwlIL9nsa2sGIMVcy3y+nU8iNwnmN7K6Gw
UgsbYrHgzibqHAu84v4Qn0IFY7XYHpKaN7Ls6T02I1iGl3yOCznjbe4CheNjlZ5vfELRmSmIU24J
iVqfDZzEZ/kI35SAYgBex82jRZnDgDIDYkflAR1bbAkpSjOgo7wFMhPWIHjZXQMIiIp6hU/jnPHq
nJ0BfC7lyyPF9SRAMnJEBqv5bAp+5VFC21katbYJMQyMTu4Dk282hgLdkvZ9SlFyxaossxXFkycF
oLIXPXqAUsiES8Q4NKv018ywsfGQVQioTyvqf4SiwJU73Jp3EpTrziHnS3+y4H3aeuFKIaKkMCjJ
yaJzzF21Hky6djK0XCNdjcWuiRskUTuNfLZ/SWVbHClDzrOgcSs0jO5cjANIUikiTMbD7foMxiMf
qYUULY4uSY0jBK8SqMJdGvwpipnIMho0HeMTR4xpMnmGayweHrT8TpxHrl3/W5WOCVL7WloyBEgL
f+4s03LDqRnjPCpwb/RW7PYKQjITbrCi02DgQ/G1ACHA5kakfg7FBm+DmjVSgZQcNX0WLgrey+Lw
T8aCzvxsysq61xdgLifS8Kwh8t173lRzrclgrT4SEIdmu8VRTGFd4Q2QjaACDNZ31UQ9s+UILVlj
wssBG4qXFH28tLOtnFVe7bWaqxl6u+6f/ECAE0xmIEkT2Vm5kO1kEofozfUjwEPyJb8hBvR6d/Nz
Avmas2rSxoJVQMw6k0B2k44BORCV3r6YUjq+5nRtH5dJ3+dPamvxXhcqpgE/QAVrdm29amAI1rSo
PUuK1cXXUO3rmAKirPxiyt14wwCH5+XAZixVIEtKw0cWwka/8GiDvshzivevi3YfeSfoAakLonFD
ZIAsASAshCLs9DY4Pk2vjrNwRbTVzCTGQPZUNFrwoAm2MTKobEmGV3T5RUSCDyWBkCwzyYu65ehb
axBy3/HFpQL7L39c4+U8tCG0ShxmgX7QuYt3yKEAbdIVc4JiKtA13MoeJ2Slnxwrl/bCMZrsuHuO
PgEwFCMuj3lZ45vSeLJjMBRUCbh5X6jFZ4HuELwMxeEc+w5PiVYSO/zhs1kmLzM9yD+ITrV/M+4g
zP+6PI50d3V6XhvGj3wU6T2U3UcU0RoC8tddSjuTE2szx9seX/nNOhFQUmFLTungBhiqnvpWjvpn
cjy0L6HKzQGRG84F+1VorcCMhWVLTchf7fmLbYiDT3jebaYHC1s7Trist7xuznYiHSJL1otPwsL8
TAqgZ0+OS2u9HUxZ7YzZ6pQqhtuodINaY4Uq3HtopdRFLzmfBhPdt3UknjqyglB5XWZB/c6oMGmF
ZMOfslvaEE4Ae+tyA4MAApn24IEA6tFmJaBQLRZQlqk7NoY+w7X92RREd90UjEaEN1EQV+tSgVwb
sw3K0DstW8lrpyiQmdCVGMTfIETveZBtVk7xeFghcrG46+aI0jT+JA6+THhzWT0yi3SUw6Yc4qSo
Z2s0PUejl5bbxWpb1ER/Q0pJYFJ9KMBQJOwuMFl/hYOrjFxTt0wB/xbsyaayhie/h/HBgCmNtYmb
9De/sNblg6F4x87mq+p9XOg6yV8cZ32OJ7QTOdJUI5662jXg2q/uQffXAHPbAEmXaODRe8TRpm0m
w4164JrSGI4MwH26mkCJFYNUXvgEs06fsQiUFqIYcaAWAMKlLK8aBgSCnvNWnvEJClegVmSeOKqu
aJf8rmetoGKl5BQXasR1s5tmHhQFvmjRoy8c0I+9faUbJpEQh4pOCu6+GP8HCJiSEySpcMWaEmdT
NJ9gvgFoKC02w44y7U+3rMNKLLcD7sw1pP1TgFaJIPZHuV1Sy69Rk0HWIv0MtorG18weGEkViiFI
Gb3vdQW02fpBrErdkn9ZmCvmxFd3MgBkuheDx/E1DBo0NQ3UKHHApw5YYMjbFkFqMrjKv8NsrM+/
Ed1BhfTz67Y8yWI5/VKdA8RHieZlQOMB1qE2ePoKb8qorTdiSbT6yg9N30MGgJiW1h2eTvncyTG2
jHy/Did8yEpWoTI6R+GXchJPgo02P/lJ9pngjH2QrnFF8TNQm9riTAYaB5LKT6GWiY1tbiS36KSp
WKnymt+AbVhOFSo98BCAULJdOt/Eh01Bm5R5Ek1RoL/jzShne3PD8rKLZyU4WIyFTN+YEK/S5+b+
2l0vMJRWo1xE4vfVLxx2tMVGzREvq4RVFv0lTpcmilSM0WYrjAkXvUwOzWIJ8Q+tUZIAONkFUG1K
9HXWaWakIi5+MW202hqUwa4hYVe468MStq6PFa31Gv0CEsePGt3AJcSP1Ro9SqvnBRAzWuiRGHcU
Bg/Cpvj6hzgiWc4pAcuGyZxdPV5PiyTyZfAGKOE++ZgWKTRVQkh8m6HntkCu1vYyanL/1lf7OGPy
lpCg5OkPCM6waegOF3JKsASoLz0TtQ05MxyDqsP9F1r1fM3ZWCoQqNFLzV5TvrJvapJqAwxzmrf+
Jzp2Sg2eSqgxxUt5Hbc+aW3L/MtiJg8vodRh61fiXbqNj7XDshQRjwbUKCqUGGiFsCaLGjP+V1PV
s1WKu2BJMN4D9sgR/+ZQaE85otDMmf/eYgZKv0JCQkM9Z5WYZhDc+TITDU7wp/JOQR0MI3AJQwdV
V83LQwrBgj1lervuA5IiBdENR1yPKz9tKTGh3th5ZzIuP57I2MdRJoki73ePk457ghGQqHckrKgA
NdjrZ+THmJVHm5/0z3yoAn9HjvGUNuSQLdOnJXrdj026iPYNAhNnn7OZabdIwXMIsqx9ENIrzTNz
pI9lucJe5vbet43WaI3RdAnapfN5QADuH1MWrRTKp7MrDCa1dxHEZearbgs0vnr3q6+TEvo9fOoL
kEFQZiSKXqKS2OMhAEVHBLMtN9Yrbi4uCCi2AJktjrwVTKbVy7/rgN1UHYQOITYhty2rZzfT2fGV
dHNPI/pzmoNgJ1Pa4jhCTMDpv2+a04niemzYP4umy3zg1CR4U3xb6EZ0kULfoMW2B+SVfmBRQXYZ
bsb/KiKZlDkBkxfDjSpI86JQQRfQIfO1DeQVY5JV+ZvIg7v4ac1mWOBfb85WVAgNtqmc8NwKezIW
7FXLCMN4MgP/YUBGdtftz/FStz4w2/O7+IMGZDH5nzvRSNjGSC75SrEHNlViYAFoDGrc3IPLB/5K
WZDueeqhad6hB6pZTSpJifbnCgAKBNqmLA0MsyiJk7gIYYFuScvRZA+NFGfkbnvJY1GI/bEj5SaD
CxUloqMS5/K7RI0M3Vx5xsQjHBb0UOUYFPwzX5eixo4/dGKHus87h6w05ngPWHv59ZwcBO9cK12A
Wbi6sgp+8+rADUs/HffuaT4D0Y+8rZDlvuUKhMiplihDdTnlSIvcfVcwyM4JEF8is5u7EQDNeTkL
HEPoQyH9rsRu3a74W4857hGlpnaiY89mQnzGW23ILwP0/A5DlRtjeaPegrfen+ELTHfCYFhxqgI8
r4bArX+/GhxRJBCCq3K+0sicUGedgFrQHSxpnpAVK2kJqG8XuulDQz2TMVsfiasEKI+MKyIOzgLs
aMBsf+zH8PD1sE4SfEl11ghSm8Ndqpp4bIfJDdH8e0Wedellukai7aOMb2VJhF4fTT1/i2T5/JKW
pYgfQnEvMkGsuUJVQOg9fgAMPjQGvei/fM78tVjsBHJFhzUlA6bnSkfcMX9jvGiaelrJyQyBLJKt
hKU0l9NIPENvunD+GznKZ7Fjd5dP4pWHC6hfpDWKdsMhZ2m7t1VxhoyXEKQgBTYu1knk7gEQSioh
Z+IlN6ocEVng5SzYg/immEYivRktzOyiCtxs/766M4QE3dVuB5Nd1GYGRel6fsq1ot4SKaITMvdv
85XuIpddHdEFObcJ/iFNZtNu/CsGIPoGa1mSh0QGpeoPGxn215odVHxYZGe3WPwbxrlZT4x2yN4g
clXOhzU8trFmD4BTw6VzGxo1XmLEDKsoR6jGVmgtUuZVOy+eyhh59o5bVIv6Fz49fhhuU/5EX9hO
vV7vPNYWeX08F/2wMf34dMZ1CJNfMo6p1gFRu4ctyVbANTDFBLR8kbq7bQTIRNYLIXF87MOseZ4k
y48F3LaAwsG05KQjt+9KXZMyQ5Ge2uH32mj9ofxjUqplV4GJza+222aSReNejUTmkdE+VbzEyfzC
vN6ScneZD6c6GvY/m8FY8ZyCYFQcTfsN9J3YmQv87viKQrzSiuu0tSeE9boaEmOUWrXgvArC3q+X
Eht2pcYVgFxBV8v1g45+08QQCZx3XzZlhoa7E/RgZOuK26eTTngdvo4/XFAcICzPsLkTqYyMjqQV
v/Ps4hSKYuOUz4W+5hfCh3vA/PGophtHQFm4mzfXqNZENd5RsbbJXHUSD1Ts99UPXWZvjk/DGCez
KAkkRfnYDH/di0pTwc+e5P0fkWISvWXXLxC8ICJvWJLn+ZsN9VIi85eZ1jGvYOGsvjm24CgAFjiv
B+p0CJe6tdwjWjRpHQND8X8px8FPnE9ehclnUEWx2pQFZIc83qBx+kWRiCPzMeDDXs+GLH2u78tf
FqQPvMhTMgOsgCkozaX9d088TPOLnmpYG5rKNl3SxxnduxsIFyztbZNTaJ1kLJ1ttSRCK3LRqEOj
vIBBbv5H2PKIiwWi40FHrTbDmvPXl8t6CLVj88pXV9bbdQOHa1/T0uo2qviHT3oa4dgG4wDllzfY
voZeXLI5t+estZnj/L0mu3KwJSprWIGw+RIS4sobDOQJ/IA9sk2HaBhXiAfCxQUA20H6h0dKnUSG
Bqxqp7vNPl/Cus23HtQ9dIwm1ZVne5BpxVC9RNvuuhD/kYAhi0O6nzWvrwLPExYZz875obKh2aU0
dYwfCjTdzp/1FTwA0ID7WSXZm9uq+Z7UDrgvrP37hGgG7OA6Q3mtblQsSwd1QRvlyuVBTgz9b1j0
J683hdfNJDMwPiDCNp349lOgo6LamLh4OME4ckaKlEe03N/GlTP+1+0ngaQY0pJQIqzyL+GQI4Yk
5Kk9jZ8c4JWuP18Y3mgmc72KmwI2PS9RooN21fH/5/GHYdgYxTKrP9oTlkmGlRsjBevH/V8xT1vF
JdoVAk86cjdxmdSnozYpwT1qL26dF0Go9o8YEjrC5z5Htl0mTiOa2tPKhFk+C+fNlOE6dr2AmsMo
4v1CmRHvYVnLQl+OYmMQlhlTE3IUKwB4dKWiRb9V6NDT8NWu+vKkMA79GWIuh+65hzolnAGqqsMt
sz29ZLh4q3sxKWfT3RmbsMKGGq2jRB9YTyKF7OmTxHXZg7kun5cmSB2n/017RdZoLHkmImetT+Og
GCG00/e9EaYEvIfKwpF8Wv7QgBj3PtCNZtFU6WChJdO2Nvlrs+dsrX2laUTUKVR9Y8iAMe2Kt1II
nmuUGRnbGpX1Zu0o44qxntHfG4JKyufh1ziHff+R9jLlq7PnJwwmYntOO6olQiJJMOgCPCW4X1bw
ujWHN+7Nh6N7TKm6+p+npSiXeTv9fVKIUWiBfp5nn6DWE65SgvzfXgBcYU3T+QQmMggzTPl9AZFG
dH83FGrZa9XarYQbw5twapTP4aJK5T8XSNN7hlxle7sCrxNh5XzmLYtHWayL10Mw6OdAxqHEbp4G
9Zha1NppbMj/B9eCowHunX/JwEQ2tB1JbeeJUvTJYFsjpiqFQRP3N1NJYiAkygE0AI9W+QxbxAHr
ekeXu3SYWUX1PsqPMZVSgzYqyG59t/Helz6+PMqrMM2A56eBc0ccKwNniTOkrpI9PgDd8puX/AOu
imoYWKI1XZuUfVJuBtDuCrI+VTTv5TCG9/q9e+y3Q0KQDCjS1B19FzRkUIkg0QulewwAdVLv4B0P
OOLIiDIadzGEhd6xjPW5bzt9cLphkeTeTEoXVutJ2Ub9BzVygjfXUHdlyOJQdKEfM7aKbRLB5aNZ
DPmZM6GclniqfqmdKKw5U95YKs321SNIbFkCHYKqAhRAm6AWovob7Jkjut+12MjE4Ae7NBrKQ9OM
ux83fEdiZU8LvStwLdSdzA1B4QdkbmVB22q7sPS80WEBKHHkgKVOaijyEwCFcjUq7b4piF5XbF3v
UFwBGoj5poXKnr/fq3K+3JXWkSE5s3K2a7COxPDwVkxYODW/3voZ8JR2kY358jxjkiAqp8eG/1GE
LGSH62ZiFjcNWY5WkniHvuNcPMBOvyZOroEv39bnQaFj2SOK2IaFY+ESHSNO+2ZOKLEatqy03nr2
lbE0pyVUb2vXebDSsxjPYKf/XGNOVIPjQujshLoKJfd61AtN/5d0/WmeOkcFHydZtH5tXksNu0Bd
vIJEvKBA+ZJw1Ly1r1MOHzxUJlViJ31+adxQbwkIhv97pmTzF4IBYpOvobBQ2LME3JD3mD5SE8Bw
xfnymR2wGCLUkFOye/rjVQLWCUYWUyG0iitj+EVLO/1yhNzmdJH2xmoueJdWs41GRuJC/PVjJdc4
6kl3gCbbqQqC7anWs+Z2daaJPmsJXmJCu+aPHO5Rajrkb+wICHXy5cZDUyiRSR1tT3zD5mPUFYxD
Qse0GqsQqqI7khpHsrUl75fxE+6RTzhAsUzm8zYQqavsdhuWkLJ7LyHUvpquuL5Bt+6DpAgNcR4I
COfubPywEq5mGYaxjcleSrx4NnsPCWxjOD/zVR9PcDLuPMqfiP5TrrucQx6dbsHZD1HTN7eFgMl7
CCeUQH0vLpCPmHIo71s9c8kn+rr1Y0Aj4iwc20i/2zMiansihfT94tqd6FHwTEjgdrW+WgW49Ask
pqt1ZIx9z7z5Yh791oR9PbYibFvmmYlBFdm9YTj/OiLFQsVg+RWK5+/GWHlMPNhGP8H/VInhY+yc
5kL53KRWToygBUPXfcOvCxeuziVGy/Eq2q2kcZyEbfIA0rXPylyJ0WExzOpwRRygy+g3bj2rF7RJ
lvmWv/AC2qPlQcDdBGps2mXb83ZPoUKs0fLpzYsBmg6FdvnXZlYFG+l98+CNMrjFNocDymv2VH7L
HCEIX9y2jCSkp5o7ZgpxrdRf2ZFqYYOBeTLI47hIwccQxZjCbTbz2DdOsotY30H6n2vZkqDrQite
HBKF9wNKz6Vv1Wm4pUniHpPbmKJslmbSTgm/SiehEDxUBSQuoy5seJhwy1aWVbG2VcBUOYXEG1Jh
vIbfSF74/KvIezKX9qoDGBXRBMcenrTah++RlPgKjPPFhMrzwKyDdL+rTmt62sMZ7IHW4CLz9WfK
GswGkvDp0IBu0aL6T9UHsaTLdACLmQ90C5Z8CzODtuzFh1ebSB7fbI4u45wEcPd2qR4/wsZ67Rc7
KfAyJujsYWBSD/+/m+Zgr35qIu0xlNMIEem+kEVnf0MXkCuy/khCWSEVkahzw6c940zrF4srZLLh
/+b1ieDKtQ/WaeBHZN+RgefLfm7neZCuh6zaNsXq+O1skTDZhTIpq900+dXk85yK8y+SC/WMz609
O/LllD9Nu6kt3hdMaurX6xZoBugWW0tU9yv1fWVcBWM4G5WHkYoJ5IT+DWOJHzZz86DblZ7dwSuV
nh2jlDjly9L2KLmLYm+j8jx/ZRW8CiUxYJ9QQMSJP6s0yJx5z2tpnvuFaQPhX8T6N3LhzoT51Xo2
yVtojUnVGhc6/I/o3Hc9vDTS2W99MqDjBTziylP8UXjRcWpMgmN6QIevLxQ9cgLAsdpauqdLcFIv
6maWtNx1Py9hGAh8KWf7e4kpDL+w4NEHygDRT0ETd7X0PDzgFJe4+FPSorvf533BCpQIpR+bNdMF
gfqJJ3OXNFneL5defiBfVat88xQYriTzv/n1VgCukQNUpiDVGAccBo6ZXjtciGDYnfCPWps5TsAF
5WwajMcGpBJsOH6BZoFAW+y7oRzhnB2bILUhmmR4bl6vHd2SXO5cLTaR0SkqFyTeXmZEZE9QpPmw
+AlhqxjUjpR3Bc2YB3nHLNWAqrJo5r8lx0WJ9qvceQYTCrB63UEy2s6wQEqzBOjESyJSZpe4HhDc
M6mqOoIfD/7Lb9yNtWwaNFYpp8GXMhCstfp4rK9bu3CXeHWrG1csJOuWe+vo87girc6B/XIS5bEN
dmcfHdr/x5TF3iKEELJLANfJwwXEzHdsSTAr5fHJ8hJ38nGijGvM/y3A4vSXeKxOuGjzNZs+MAYL
IVVr9TPWa/C+0ZKikqGuPOu7bGvHNqoW+b+Hqez4sb1mFhmZF6J/IXgUc8qfLNY6Zz6sJpqI58va
bX4lmYVF7O8k3Y/kcgSfWaJm5uSfu1RWrmriYF++o6/IZGnr/ZNMmILj6Sih/7X5RBTyZYSx/fPt
JmqRw5risS5a98f9jXrCvANRS3rAxQTOMobyC6WAOPTZWrRk7S9nwxr+8e9oIXQLq7ewDsBni1O+
qfMjjjOZlVNjZvYBjwqlF5U2Hu31PIManwibfsGIASnCGjHbyH9d880xgEm6ukzMwFTVBT8I8xXi
KdnRoMyv2IQZVuCZuLHhXCpS1DKVzl7XpunBL7BEQWPJGyyqCQ6H/J8N0QYqCx2yGatkOx5dFSnv
7Ax2mKeGWKmuLYs3o0KxeDR3iJVdyIr7jaLwr+rD1C2B/nMYT4gUwKt2TeOrkzgrJJ7T+Ln4youd
yQKLFV5p7OQVLBTigcDY7LAQX23fW2zBhzI1qL6KWwj1XXpAdpU4llUSg+cKNI0s7GIN26HYawdI
RmG8I59dgQLdACZl8rwQl77ovEpG9FOGLG6r+xGb95aYkc9HtGWQsYCQvSqPge12l3ihbATzIoBi
unKLQWQNHjUrA/Pf5E5Xq+nDl3jqBSx5NK7F52gg3oucqESuYq/89JfVA9yWndOmGh+w4wx0fZC0
8FJdt+5srPwbP/oU39pHwerAZQXD3nxvf9QiuiKngwrnqf2sKGP1de1Q7HHRTX2UP1GtUdbW7FdC
ulbuJBipZKalFWV7KLe8PgyCxoJboydbwsAGp1S8wBqlWLMLvIqR4Pbj+YfcZikwrm48N5ExUGw6
nuwfKT0/HtBOXY7RXUGlhmNg0Ti3mWKxI7R7sJbPe/Ydj3Eootmnj3LcxIg2SgDUddbpcu5f6ObH
E+81pdX1P0cB3y7lxoPCRxSiIAavmQ5XpHHhqXUbba7Ei7LInkTqeccZIQMQDSsg5cCQvX/zdkEe
NQENiKhF5uaBR/AN67fGZDGIvGZ37/agbX9/5BQu8d1HFq0ykZAV0l+aWRgR/oVJuaC68YnNkmn9
5GojvWS02saFGWEAL5hpbqnxXiA5djVU4HrqNMzaMljxIGBwmWG8zYj/3nD60oDx7OtAC/lgre1c
dNaCV+wl5UZwOIdWuDfIGGFqkGBDMQ4OXuDaZb9VmbuP0cRSlUiwxs0jjUG/rWFC1qLJEZKF+29Z
hYQreTVAwqq6W4Mljat6W10CsWBF2QnRXlY8hm4/fncogR0b/XPpu32Gaqv7pYpj+0chxs90sCNf
3PFZ77YKutNWcG4VxZJsnYek0FEBZesPFmFmjrBoE/+4ED1LCYFlg7bsU4omtJY3+/cwV/8GFIjN
H+2wmWKf46e/lKQE+G+eItkisTeUrQQh71kApyVDCII8OEiJ9mX3JfHorieXw6n6kQst1Mkm18Ie
iKpivQKFRJ/ouFu4/kIuBfVUaYmJed1B0q9AscFGp7cJl8JFN9fCdi9SGg/sF+GyMXxa6nJ+iXJv
SFpeSKMpzeRmesKWPaxZ874H72Z/RhuCwwfClwoPa1W137Grbfg91BaxAvIXeif7bE7a6DTgTr6g
gKU/68DJlsppu0/jQThcbwJnLHvlBlOsjUvIFIxPCuGI50ch6SEZEgpxon5q36HdEAYDH+Vip+3J
Y7z6vEBi7OsZ/epdWMA6K1sj+1jlfu4D79ziF/LeKj2kMqTkFAl+XNhe7A+pFVVWg9hQgVp7quEp
xFtqy2esSpKXdTOjHNI7IGcAYno5DobHbP5IYirxfxdIcYA+jRYDIOC5cW0k0Io0nHFZfOVRF/+x
2Dx4i/sXDk/aoZhdepwa1cLMq/EbJtgvUHhzoYyRzC1Dgsz+SZGvzebi/RjIe62uGCjBTA/FihnC
gDe2tEK1mkO+rzWoWWNt/9FosOuR+bSo3B9c6nA69Wf8xBJlFn3vVDNWIQe9LnDbtV9xVbVnknAD
8kKF1E3mkczOiJ8ytfIk8700zSN/cAZAieNo8BE8F2wvIopbjCPTSO15B6qk5jAEZLAHniHBK9lR
kVCjqIEo1+lgXc8FBL44BSvXbisM4Uej52BmHBDvJCogSDGdp6//mPR4j69gW71adT6Tue4/ibFE
T8CebXerTOzg5222DkkQGuCXQPSV/9oNYxTjxTlNT+6ROgDiExhoO+/Gmd4sCuWxwIACl3DBX6FX
/Anl4o4rYy83QJF1hTdhiHsfFCDG50YLe7IivmeF0oXwIp3iP6FHuGQieC4jC6j6UxAbmoivM+qw
e+w/tWI3LRQPg+J6KPww0iuZRxTiq7uu1DzSt/Fh6MbtWncr++HH8oliU2Pvlqeq5jKvNvFb/Z8t
HYRvPUwN+Qyw2vMg2w5zWWrrjKllIGTWSl+CBXlQYKSTGtjVTt/lZuzofSiNLr5T982NxTKVadaK
rwoZEm+3LXZGbCTtDM1eW6qgn05S0pXsRKWNekjUIiGcRkRXz122JElpQdpj2JqABHbiTPsdeFL6
4Jb/E+htJ+7FP0lESW2E75kfxz1JE41m2Lfju2ZUP3IQHKKn+hxe0NxD8tfUV0uIVsOQDyg4Bj1d
SqjwQHWz+VKpOtkBTF29pfDxZ/UCOhL5gOXGWn07Iyg9hon/70B5zQ+LMaT4/KGO6YDeslEizxgW
FF94jrCybA9sZDNkW/0QeDIxtwbYVmEOwE6nBDlWYhR99W85c/S0BgBfX24L1rvUFUmzXGBuetPV
eIWn+hNFoVq8E/3P/BFcL7oE+0nRAQI2+vV8L6AhWlSUhB1AYne0//ZVr2qAWRCMYU+KzW5s7rzz
PUQqIIyYfCCYK9bFVBfKNOheNrhUgVDblTizvWHMkY+aKhnk0ey4Onqp9e2fjAhEnM51dh/Mm4GE
2gvzfMZOf1kJFphi4vhbViu5P5TYAbtJ9Pt/Rz86buzsX7mZxnrBW9S6GnE/It1FWkYsGuuXc4EI
58j9rMpSGY+w7O9gvrqeAomkMFBdObe6WiDogxV9OG1OEbSvz/cAxjUUfqx+nptGNBmeXLzclvaX
uBk4uD3O/zfOfBYIVnTlyxjfwlHzgHkLpyYNYWjDI+vCdvp0AubJEugsXgRsMWG+4Wd/FhYSkGqY
RbflkwMDmj2Z0xCBnDsWPo5naQGoSsjTVTwnxcgYwVnMRdCkFmzOpjqsvpM0hfIneU9LbOEpBY6D
BIm151PlSJU0M3KdAwEi0YxRuE0Pxp4IrVT7CfsiV/X0AXWtHCvVrgEErt8k/DY3iqG+BbaXOzQ3
s7u9n90gDh155Od9svSJGznIwOKitFnFtrQG5RnsEedMPoOv1W7m0jtzv0rSc5Uj/NtvBANQkuKh
i4BXLFCPFhd2MRAGEyaAgr0MJEC17HuJJUcaj8oCIU6cWvyy1HcsKqgSao5vVsFRDY4gtE2NAIoF
yajWHfu28F/J1NgqEVkEQB9TRgkhWL5Y2Bhe2bSLgII0UHi7fCZZGkct//EP+CvtXZc51zzAmFjf
qp+mqpfZI0rSiBQUW2xbIFqEjdjCmi5vjhCiegaPgh/3mC0dcO+HJbWc+4kVJcFMYm9BScY4qDi+
tD37qnQm8iIOZXRrwK1NXI8vHrgCXP0GrdCoJxU/psVbCWk+dAkqhk71iU2tJ2UuyZKzJnzWENO6
zOqy/2K2/C2JjQsA9LlgN/RtCZ7CqOU4QfGd4GWXjXmUZKRQH7pxLffCn1C75vVLzbNBg26e8rA+
RfYH1C31NRHPCMUIMI70Uu0PvZ7BvsQ0QjyA4QCOjEn54dBt6+pHQqWxhU1d4T+hRKdunhyQKtHr
uxWwZj37JABdfZjE//5OxM1VJPMCmzykpcDvY2jzm3p4fiYSWOwTODwUrwdsXoNZeAfQw4lfss+X
OMmTNbmbsKXLqqgP1FbiL1uw+8B7pJMNP+F9lHh5CoO2JyetyQqJaA5hjA/DEaafr7Sn5caKW2jl
zikumnIXKJypDtObtRSAT52pTQMvmdH8M/5Ch4TN7kErleBMsD/WkvgDcNabjnKkmj+jKp1zaNqA
N7UtBUp4d25szPSVZP2tQFdTVCGMjM4CaT/n9Z5QCv/7ElM4T17/vVDfglk5XDAA7vSJRFmDRL+a
Rd+mdHdxD4gQi25TBRNEwyDazzelXkGL4eLVkQPfmCiIoXsOsrmL+lWjMcroOj0wNXKeM3NUhLLv
vL5UEE/C1GO8O25s94wpiV9Lh/2elgg7nmiZGrs4itr8hwqKMp+2puZhU9uCcuZwukox828BlIcV
bmgi/h5RZlll1plUFd4LEAokSFnSNcv7pmjoFJLJLEbo/eMRAHOXwwAMispt+GZr+HdDG/3Ca5h2
ajJbMygdB/RyzR3p9oGK3Axcjf+ZFObs3m2YXUO0erLMhMNgMBWVdnOUuzMje6InNOJB6Ns3mMD7
nk3AcsIKVS8v3VycdHneFcgMj3sOnuFOH0BIqe7DdI6bb9e4Lml4OODG0iWFHYNNgOpHeEOPGK/s
DxGpxPt6P3n/fWgNezJQcEirDJd9PJY9L5jF9DjWZ3C6oyPiqBMGDGuxSd6q7D9aBXZaRoS9icZR
f05DGtNDStXwfKz70y4e+CTtKGpIO8LUS1XrD2M+JFMqT4TtJWu9G8FQKHndA6jan47I4w2LifjR
HCHfoi1Ol9ivRW32Z2YR5JgDvX0UzmJeMat+I3e7zTRZ6RkU/5Fd2yGFfbD03VxDSiVfr1y6XSfd
Lu98WtvLWZCXYAut947fWoN9BlBsZSGtfXrYyOzqFJNxkxRK+pQgdpeUkCyCr1Dzzu2TdocmbSkc
aE0s5rvqhrc0V6HO4uc1NtezmpyOQJ2Pi/Q/fagN/NPpWi+tWkZeKZaMqjrxaq36y+TSstF71EW/
aBH1w5nsj9CncGfPfGOkdMlJiT72BbwkOcatlJa1A2UKU0aI3UkTWK0soUh3J4xrYcyiQXWCYJzh
Cfv6cdHrvV19RAJhUCwLDWyIsw4DyaAB8jqAvQAGll1H0gTtHeKEguALJDtlqSqIednBZ9bSjL/3
c27u0X0o+Lj3F6msiDqzSducb6LOj8vgbnTO5KWBCCYuFs88Y7JeOg0T4pWx3fvNJa6rEkUjpifD
bIQOBU/VDnKuEoRO6UR7x/gclN5WXz8rcbybpKUJSZlpFl/N74/8uyqAv9z2U0CF0ueo+mRe60rB
bG+d+L4cVLhh0ElDATRw5cgHib7uBwR7Jodyn5eAYbuKuoSDk22HmmOwHEFL7YUV0xGRwfQpTWHf
sSlXwZxPlNtYLaU98T1fMoYKb6mRILZD9jQFKPDXAyXz+G4iaKijNe6o0CnrwQbAQXvhTrZPtNTv
f/EF9rNdWRnxwf77jP/tTwsjeaLJVzFCOFWtayCLLeXpJXeQ1smH2uUOLOtketAVAKl+60ZgHIWJ
ic8N/rxnzpnMQA5oRf+LCTWBbn+y1I6dRdP+P864D7jl5mlJja27QgmjUjO2S65rOXqayoNtcnde
FuSDAyfq3UBH9NpMqU2Zf5Dc8A5Qh39vYYcNJIlDxwdNBitj7isoU0juttFHJEeeC7hiw4lV4FbU
FbhZDSV7AIN+K7oqDTT26UCwXt70h09UfERQJ7WNYTlK1wJm7IxhXCLnV6q7c2P86U8MRgqwYOO7
es2eKN73I2N3mGRi4JI9Y4fykouxyJb971Cr1nfMB3EmKps5LgEnPNDTlPoqMrfPU2EElgbuvON6
Dl5u8C79g2VZhXkRAxi5rebVVQ1b3zhUm7fzDX+PAFbbu27hQAQaKf61w96iMHaaAtjad6n7odOD
VgJQRlA9lifyplVuyeyX/PPvpdaOnznMIVnkXPXw0x50gwC+NVRDcaBWqM6LVbA8EwWE63Kc8pWO
XtCPdjJeeGHQBhhlYP7AFTQP3qWoBxSYrxgMOltugH+UuZQmV0foCQdZnU8pqzBFd85YtypReJ1e
oLwqtxcwT2543SkCBt6a5jamr9/BKB9WETdFUGleKdNiZAPdKVr23Tft4sVhF1+DQYthkwga9Ros
e/HOdiN+kFqBGglUzDneW2XMQx+Cq0xIvWlS8ZKmJPo4UQQPb8pUy0xDsrcO4kJYFK9ZLz4sE56C
2o1Ls2iynFZzM44bubox9KdQzBRdo5xtHzTY+/7wdR+mUYMfoI0Y82N6a8GsVplsipELYKtZ6+B/
pbmqPoFykBw4i9K/yPMx8HQGTFG9wRUjk9O9lYFoceKgJU/iwtX2crINcsyBKjHPZpfBMDrcoeon
/ZJUV3v57b9lDlWz6WweOvZDWOkD22jmcjJC+obL+Zs8RYqyVe7ZJt6QdjmaRU5AVHYxzVv920OC
x7b6F1rPWXf8rdhWEG1Jx6u0hBTcQQbSh91ViDfRyPxCwrP8//4yiow07PKzX0yIpoJ6OSTRxAMR
vAWsZZJQhOUBvGLlmsdihu8BjLlyIjlBobvjLaZnHvrx1Ul2wdccTlt788WcX3xIDf/f50QW8w35
Eoi8JDm0jx4XPxcKoUMBi/O7wj71IquKol9lihimPorjxPpvERG6k0m0O+N0rwg674X46+2xCTL9
RC7VYy+JS7SfThpvh8Tcx2otv+crGumdNQheEF6U0GmjSBQAJd2/dXdyeuX2hGxQuqVBgWNEMQrF
QAcqHyG+R4f8jWI3A8cT+e7nMTyio/o+DaFNrldKiXAHTUPxlLdHVKjwAeiZjmjQA6kJ+d5hERbB
fNdWgSYp+4mLkYHvWBY2UHHWdOk2ene1Bc4gokT/62Dy0QSU6WDbVR5SzrY/vLaOF+HCVo917QSh
+gmW0YK4GgikvE5OkcVtaxIyJFUm49iKJrdquZXM1oWmcoOzjiU3ErzwE2QCh6kn+f83B4Q11y72
LGn4LPnK/QviwRK97RMXeEFttLBZIZsI3M0eLFpNoniEU6lovOaQ7LYJNXsT2yYxDGtXCiLk8F55
AXlJmLGr6uS7WvnHwTjiAOYv0rhgocG9f+XieLZt1VflVKgxBs1alB+eoXL/UmO3aNrqtCSTNGUJ
CLyzPNHc7bd2VA1iPpQRf4eizWZvy0UmVYBwf2nWp2Or1s8XtgvtfcHOPp6XJbjyaUDMXHjb6wUW
7PERlgCG9WngYeoMNy8TN/eTErU5cbNVFMh5DNOV+6BydDi57gtjOtWLbEE6PXj04q4vmEu9V/D1
l+kV4s8k01Ox4JHSs2HLMnNG+ZMIym7ZKej8sg+2VocGTpr9ACcVXrJHkX+rYtHf5Ys9AkI7uHor
0W0vSSEIogdB6Ml9suFgALvO6IiQvMKaUCOEZgiMTR4n1h7rcKzvUBbIYPTUDLFxJ8i6C5pdvCwy
phE2thaTWNFiF/Ist2SCqaW4/+Htr00sQ4AjfWcr3Wx3jLIpLFXM6bMW671oZ0tgNu5LXo7Q2LVr
zYVQhOaXi+qfDZlb+7mZYrmqtCbp0uRRnAZczIuNUjhKdvs6COatxh0iFw7m27Hu4K1+IGcIy0lp
xOC2LW3TzuB7mti8LVVjlAa1QHvS8q3+aWEEPTxvcvwYvG7XHVOppbOkmj9XKTXZAhissAZ4sX9N
MYWj4KfJdSaDQYBSnElfAHxTjiPGIMWoW/h6q353o8fXzjZ542P3hTu4l/oik6U83fT1Gsk9LxIc
wTcvUuxY4Zuk+IEdbpFs4mPsEhqlijPWzip3e+1iHGNKEdBm3bPeewtjWLfS7UVW5HT8KHjnJIKE
3YL4v5r3BJ/25zzJcfCDKVpa8QUEjPTUgsPw3tlgw0IoKHMQBDPlxZechyJre0S3CW1WsHOrWSQr
gq3UPLM7zcTVL3yQwK+V42zqztaUPmQkBbnV9D0UF+6BvGgEu70g33WjnV+rUVbDLUV7cmglPHOi
pM3zjlpasskzcTLEMbLUzDN61sTDBMnTGzsdrjlAUHALpFUQ9CQNT+UAeoBrDLiHic4accLitNJB
hK/d/agYDUtbLsoE+Yx7R0z4rmFJMwykKZp7y47P8BhDyhz7lI+Bi4alyxsEUHHRiBNIJOeX6N+h
xT/yZKbR5o8N1owUmGzw+RaUGF5ZZt9/7K5yYp7iMATt7pK2GDnaMSSuETtTTCl5g5zaQKOq8abR
NOoqCjwf27Lk5ve5P9+KIBHjKY/rVtGMfPRpAL3gDgt0id8ACx55culhBnDl+6U8pPJaR14VEGOv
XXzJpsdERRohgxDBAza0aEJv0+t51e6XkMr9CF4Uez19T2zARCBxwmpmgAAAtgJ677IPTltD6HWm
sip8aVznpNApjW6Cy0j28w1QihGEpqplGzXuL7U/iremgxqC1zY5PlIcNYldejeLYiRKtu+zqBWD
38pSSoudTZH5qFPpklKpSZpv4fW1JaIoz1VTOfa7LOL77a5vxcemvc40V/x8gXeDH7KIXnI2TArQ
58XDnga7++dkHyy/GKMJDT7rwy+t1sQj1HR47COoz9ZG4xWMniGvhxzJDrUFW+ZTEPsOYYgdhRGV
ef2IxB7NnZF6nTvvnhemOg7CNhAHGfYCBJqyHxgvB6u4rnrqyclVG+NSyvcVfUcQwCFdnbSkbx5U
AGY5VcDH/XDO3L2rFD9PZgs6dEik67aBxUWWrcYY49Fojg54+oNlUIPvDThyI1ov/mdpcjjO8Ibx
68FlO5uaFHig3CyAcio9e4uNzJxR+iREIMZHNVrBzi/cvl2CEvWB4m7oDXiV2l/iMYu/XzIM40Se
6iJMLql/In45R4CUbHkdHL/4gjuxa8bNVNtkSns4OFZwxbfujfitSf45+R2BUaK1X65lFIX8mvoa
zw9wWIj66P0Cvk51tiS0FI+0ycgHXXGjbAqSf2KZJ9YuFW5+NPxfNQDUQ0n+g20+GAElFr1k1AW4
QABC67MLZv+IQzr+sH3Ift/lYHa4n0DSjY0pA5dXEtkZ3XGuP3LrEyvMvqABsE5MbItj3iWou0qm
ML+yG6djPcEFC8QyBh60q3rX+NS8FgniffcQx9hWvB2OsY+s9EE2K+rHMBW7J3n8fvlNE0+xd72b
z4fSDu+/bstnIyQstzEIFXAs/WO8KBMAHoSABu6awdOxTFLS245lauY+aZ4/agh2rX19qIUl83dJ
oUfpXBoTScLxLApN0eNcg00XqeEFYZdc4VVWhy6k2u+euSpaFma6IBKuK6e4Ld0GRL1Eu3/GQhS3
CT2Fz34gjbEQ0AXGa/2QFu9XclA5HOO9zZkgatjB9kwcLJm7tX/3+mKFqhp969lbYnTzqszT1+wP
dzLqcConEHGFhVPbM3rLWBaFu5KtiUo+42hn75eMMpzyT35FVRB3EgAWRSBkQyekVob1xKFyshKF
DIGhE4PdB5et2BiRC+vB28GYf5h6MCnWSgq0OQRc4qDnd3GG3Tu3PKI8vtY2neFHsC9ToGqHaGM3
tCrtgDAe8V4go8ConF8uov71PjVodR2ueT7THJ43JFaMaTJyPS0NaCshfe3sKYTShpw1b3mxSC6V
aJssVKi1Pk/Tj4l3VhSDxTHUKPEceGCOYVyPT9H8I22ytUsGoNn73lxF35ic6flK8JTiV27r5EKs
oZmcYPSq2RLDxmIXsI671w4/ubMp2AgN3npeDMMbV4QAaq8xp2zDY4RrXUZRVugCTwiVQgP8mZ/R
2wx/sH+tEUMGXlE5RLeNYH+MK5KmTkR/ccfp2IIg3dRrMTu7HB62I2qc3pmuR+Cbmerzg9MRmuT9
ZAsnUN3P+Z2bu4QdB9rsHEC46X2G1Zztxz2rCAT8CLriQEAWT4q3I3Ia0lBcKbItN7f6U3H+eJdQ
q4HZIS0zMCs/a/KFSjzPPadfRDHhcb5cEWO5wRuxCfGFpObcqV6O7/X2Uud4V+H/WfmGWOyaOtIn
cEJmkM7pzV+6SFgc5XvmziSupdN0Q7DBSDGSey9lUEpswPiBLfNOm4UH0S9zMAAJu3tn4lP78CYg
kmW/woVbZYiFGHgUwSCQi5hsTr1ixrbPA/8DVPYRQc/m5gsy29zHCJVs+IgOfcfWVOeMv8kkrN4d
KtL+2h9P7V3MkTBZa2XLh2XJcGT98YPUGMt214rW9g8sLxi+N0I5LWRXvlAXPOZ5X2eon/sII498
C7Fcemm42nWv7uD1DJB+UUEaoRcOfFyN33UuTqsBd+eREF9T0o3++LwKwWkUuBafkLTPHwYBFg0C
RVPuc+Mt6CG97t72lnZ28fHkEH0qBIT1qyJldu7UgYl+abD3Rz2Nm02M0IdIb6UztAAXuy7ZpGZl
8JTrW2f18u3aofgf3l5PV6AJLN4hrQ9zxeyPH3lLA3s6/YEBPKYPgWE6/smMkOSPZyrfkmT09UGm
/m26newlaFzqqc2or6mz/bGcAruWc21obkaAdVlI38+OgXPOZD49otcJ0G7CJroudqqL6Nd1/yxR
qP0IDMI+kpn3vP5c7yc4KkS6NOupk5XboTx229xdJ8SrGy5oYSPTXwod1ToLsa7TIVpGUOMg3F2R
aqgJTta/U8B1YszlYyIAhSjLZrfJ8U/aQo4uq6dyG5iKbYlLGsDkXP14AdZCgK1YQM23+hL7tkNj
P2l6RTEZStFEMnE4MSY7dVcCy7ct37cOgg0fVl7ZiR4yr6+0qX2BNwOzyF/l/is6AareE3MsuIjP
Av2TwsJGIS5wBGb18FQxj+eOJgSud9XBPBMyssBMuUK1p1wWwjr75Y7rci+9ShlYT3pSl9aCeazK
7g57Mu1Y6DO7wXM4Y4iAqN06Tk+cze/katnvVJsQc4kL7hRbiWPyDIlp9FT5AzVKCqhCTAz74Jo4
h2nHEBoZKY3nEpBYm3om0XuNkUy+WUGBagf8xC87Ufd2zTg6HYaT/G8+gKGXYHgF359zqU9CeiDX
A/KkuEwgVkxqhtWOAZskFfj3nGk4J8EI9bJS6TVgmlqkYxM566itCazsuTuq8ugqBpQ3Ve/JaHr9
Xc5pG0B+FpFPaCr6OvpfoTe9VcO5y5LK6hRsH1bcbmQkRe1bR5xvdN1RiYkGVigCIXBbZNlZQic1
NhvHpDFgIH1Gc4B2ZCRxdiMOplWzHzY2kWAeuRTw9WR6BVAlN+H4v+5fFn21xbA8xUDtB+M5ufkm
AUwcybCYKDj6WFR4dwuYYYGNm3gbsZhWu9gOOxWmBnzo5rntUciryTKGAnzuTWmLjwmQIqFLAqxs
tb21tUpSKreEzl0Lt41dV1L4b5fPDtmCKPFkb1sUJ6dRUH3wxWOotgHFVAspjtlBegJrJv90LpAA
e/YEuwGQIP2qtEVRKyKoSAJPjw+f3Lz1ZzcEtV0kLsSb30h2EQ0ohXapUnbvNnNx9nBWtetXLmmF
bk5eKsLsco6PD++zm2YtPdxp3jbBMaon3D5AGYbhStwgWTFLB4Oafl6jqbCbMZS7YG76Z4N0hir3
culMsFN+mnLpfojZHIfoRZJ0Y2T+QM3kYhYXKDpjVcC3d8+CA5sYLmoNYr2Y37IvLo0CDLFvI7eW
j9RHdakSwNofAahENxroPj5/VGl0SPlhz++PRILEfAAocj9ZXxJdpMQK35SwU6agVPHNviaQKRMv
+h+MQekSKgNl8yPwbXsVb+JnauGUWW4qfEuThK7Xk3/pwnhElHJcMaSTRVHt/hfPibws5zu4ywXN
TjbOjruL4FfgwLcYIoue5PuTOnQrE6Ztd7mBOerVRqsAlKbigfsLkbLSMBHrrubqNxAhf4/kQBxs
JBOYbeVU/7KDdVwWfrHmcPwp57b4bej4thVsDEug0v8/0HdC2fOKfVAxGKMqjcJR/HDfFAmWtFON
8xbb90FviF5Fn7nIniPjomHd5ZJI8EVeQIGtte0fTXI6ijC+YMLmuLEIxvejXuZ/aRNXAfQQ83/y
Y5ER4LLUASdvNyAgEPsEQ5zv8an1Hj/9C3yFCxMXPFMkmJcjnDUl1NZ4Cq0awvSEJB7M7YnBeVF8
f5CVk12ciPSk/wbwcalQjGIvhFxmBbv112R6ejvOHtTdVLohCk+ryF3i2qsc9HVGY90Mjw7FAiOp
gwA5bpKye2OK3NgfYKwChIbLN1zxz8JRnhSSY4/L5uhCF6ujOFecz/0QzSkbTkP9lSNPrWcnPIBD
GWuS25koZYKxkDiWsJ9ZCvYII7R01xgVKQ1zgtI5mJPfeW9wCfEtoGALHzyfdDthftc+HAzEEzh1
D6UcwIoDXAMdVhiIbGmlSWRbyoAopQtO6Vp0/VRe6urkX9uwBYZ8JcdpKvudvXAX8t18cymAHNTt
Dl7j9FblmYC8gH4EmabFoJwUfceOhLHkpF2SrCJGnFdLSb2QLdKFzA14TORLHM7tiY7Sxi7s+/F0
nd9865HqbLAswk++oBmrV91bZKlT5gvv7bOKLC3mD0R1NcTtGDGZLzCb9pbNEbVesp+nwdDYhwfh
B67gFznOPoMCKCMw6YNw6zOMgRgE3EeEpTyDBcXeowz8wqth5nEqKG0yP/DDR4beUtNfKVi0NSIT
jTM/sNuRMIsldj2a8ag/xgAw3YfcKunU63d5XHxg0UK+sjs425QGDKaELqPVUL3T2zaWP2g68/A+
Ucfn37LxY6aFAqAm8ZEzl4vnhE0GWCbc1rQCLh4YB4txg2X3OVL6XnsfaHAwzY0KyKiLz3nfbB9R
pPwaIBhbh1+OzmjJoNo6525SRsQY00sJwu6MHxWCVXlZqNFkCZ74DhtD7gDFP92pS4LQwtdMDtj5
T0xFiSrzktmJyvPB5KPscMXb9LOs7D03FjUtTODtQ3Lwedk6Rwe/KrTv303BCCq7ECIAu6KWSLSe
D5iWBnQJdROUPkurH/p7BaQHWUGTsPX12JcJGs+KFtZDMtXUEMszprXP74V5XAtqQVtjhW2Uy05d
OwTjBILOtuj49sYpGnH7ODq06U6UR/THQoZe1qe3Jq03XoxOsU7qAGNiYnSVflwkXcQ6obbkSNfz
m2sU6+2VgyJ+OWHPrzo2CHtMe3Bfxg9znM4oCi1Sta+mo8BdLHUhLom9e6HOuoovdVqmf09esLJz
TIgaGy4sbXCHqfcV4Mrc0bHBxK6tOlNzKi1DdZqzho3aPTsmu3rkyswwXsJgL0YyxW+ocAZqkbK/
5UG+43Ntns1P9bRtcOo6yyH5eKUkhbF1/CnB5q67VRbjP9H6olYHhfkufozymnNyw8Ox8gfo1d6i
XflQk5HadlgEjQeLDkB/F9tLaXzq9GHP/ILlfedXfHlbblfRvzivBlHqQQltdHjS5YNj83pNUX0C
VfAKXqUUTR2rxJ7NdgnWxd6fVvNnVE6de990S+0N/KqtIx7wC/emKcsTiavLJbPe52vxI3GETxQ4
atBSk/oGYTiw1gu1MgIoruy09dUTyp55BuneuR9+/hZi2Wt7dlyDjmoHP1B/QSTdMAm5FSf9XTCZ
dlMvbMy4na+rhbsRQGyDwCx/vzcue93gPg+gFJELZgjIYUI+NtJOH0TQp33cpn7IG3BLx7+ZdfKR
/Ha+rUKtfzSqLoGR1duWOiFa5GQIh4XyQNobVUuco6jLPtJecqgqXrVyM+pvWCanTw4N8cdlQ02R
3ULmbikqKBGFOVTgJQie+o57cPEHo8qyHH5/zOB3pX/CUkFUL+e0RKjy3yKYI3XGgccm2lwE2FHF
PToaobI65Z0ccX348lRRKqRspLg3fvVujLRlFXLLfmzI3CDPKmx0xDJT1R5pu7pI3rnjsC2BSxjQ
PhCa1qPcvkSZuHQH2OrEfxUTZllBQT0Np5vpiXzLIxM/+gC5D6sBQ3L5TdY7Wi7mYpL44yyxAELJ
u0AxCh69rLKm/xCiB3kZJdvz74DHz6HiTbRmZyuFYqpI4bn5mtwp3ZFubSjIhK46l4fTacNDHOQF
iPq6Qjb2W4OJd32D0E47F+dhOx3LIr5H5KE9YvrLIqIPo8Sxb/7wakx3C+ACHVEJC5FVR1H84yuu
Q0QOIXYVSqUUOZ0hpJXEYe7xu7HQ2oVTG1f48UkJydSU/s6nQeJogJmIH0KGmEJ5ewW5+L6OfAyq
mqutODTen1NJvnac7b6M1Yd0pLTl/zRK1EwmtAFgkxuzzzSoiY4Nv3P61x9EySytWBgjrncZFeqo
7RqxU41ppRvxYkitxijbHhxn2Dtl1V9hk1KSBFt4XrKP1Cq8Rm0/Lz2/qEIuynIkioJCG8o15YFn
HdBw7OPjIS0DfLTZYjtWcNakhlXEGPEeC9Sgy0/QDwFLeK7r7AcAqKmrgSr/96HppDLmurPLqh1I
QRT4TXE4Z5qC4Gx9x7XzWwFw2WU7JnN6C9P8wiEMDy82mwVFmRlDkvROm/QCcUKwoTGg/i6qc9wN
hgILI3DPq/gF53ZSQqG4qd1+drqn9D7mV6J3HnUJYyjsEoS3F/3DfhTX6dYDRLfBK0ex02cE5XUo
Eod/wu9d8H4J56Q0AYjSbtgRNa9i+MuZCRvkMS7ZelH9Y0KroH0N9mF0dKapu8ils2CKLKJgt9XG
EDF5TfXCWULNIyBpgJLO59LsUEnZN2R5ET0V2h4M9+kJ1sAq6P6QTQqqOP+j3lJvXkVsFkMfzs5s
1sK5Am1lbfaznelPyS/RAYqCWofs7AuP0mAN3eALEiJ1pa24iTr6tIImeEjj91t/wD30fZSF1SNs
IqtVYowdoWfqdA4BoR8thO8pcc34a+3ghIsCYj6CccA/5OCBhwtAnRV1fM0ZS0I+i2CBQeF2iUC9
vb6Pwj/H2Ive4OtudbUDybd/WNHSr+EKuTEmg9sIIwAZe50kNG4hmaTuM65Lm39fpcjSsywpbzhz
HYpRM4DRjxUSKHGtLSiyE6l7ZgJq5RrzQJ0nbKOHN2M42BIgFVsAN6Ycpy+qiZ/X4eNhXAyrcHCk
X8oIg+TKstfQIETIFjqJF2ohLL3RbnBD0x0vUWO38Q0HKrg1ER15v79XTVZaq2dDz8yk2gj2ON9B
Yv3jlg/AOZ8WqTo3mta1bfgABVDZR/HXzLWYrppibvb5pidF/TThEcAecVfZCZRctQL7iOzEZjbB
Pr+lYPowKsguW6eqUdw8AK/tKXehG9LnWvlTYyRk69yTu4CW4akNh48Tdplcdhm0gi/HqrvdWByT
vDMlnRvw2Q6ZEZHqWqexgSKGJPIKYs20uqVwGj1DO09hFerbbWhSIU2TZuOJXi09SFOQFOH22+JL
wRiP3l3YWfvPEgKvrgu9lfEVpcDRk+knJFGrFyeZiYsk7JuhiHcvliCshRv7oJSNENQISAIhDs+S
GO4fRe9t9wcyIGT+jjqUIflqNcY2r00LlSd2UFG56KH5JDz5Wrb4o3QKpjTpVTImuOPQ885s6Q/p
UljoYZr2kqYy7JZ8izifEl1hJRn3EpBKjCkGLQJxvPUiDxdsIWwa3AKMUzoQLPHgc7eCUowOxmMW
avrJ5RcD1TD4s0XY4dhNdea9UtQdDxONT6g2jFDUdXjawH9lqVWXPqEw8A+tB0FxfqvwrytxHXEo
5Li51zWE/OphCsdRxVE4GHv1F5eoF3rcpKeidjbjAEE9+YLIL1paF8g26DwNAz7Em0hr+qmP0R6L
mnpx4pRhDIcxftKrdOIY84gIrrG4HgR/b1EUy+yKuzsYob+3jQna0dek+uTpGVwtN9mfffH82auY
As8ZY5ZwKQQsPKuPR7efY0O4IO4g0ZsdRV9xNB03V5SF6NHANDxNoXnx16KEKY+eNzsAV7P9x5CF
KNP2TrsrSMj4y1h4DPNzNfEZ/HiV/PwZYVrYdtXA8U+GGyTIhJH/Blstqj1fOvx4gf1f1svFLxP1
nk7BtRJnlyQWa3aHPyiZBnjEWvoicG2wV4MuhcIQ07osVxDr+FxqtO1c4SA44mCOvKyF6gzy27oy
1iyBo5YvJuvpCbiodmEXnAJAIJHuvnKQTZtAtYnRVAL/h3/yMYRZTi7gcHz0+Tu+Kz2+xVTGtQaR
98K4RI9lsfFCmhAhWdZtm/w4uV8EEtLaclkNcVfyKsHegoVGGr1xbtfLHfBZZImr0xQ5rxsOgYQT
8f/PL4ZVWUXt2Oqou/PQNpH5390POIeV8LaBnWXP1WwL8ULYM1h+jW2kuqmKJwraUHTImJUlM+RL
LtHoeC0mZtNxQodh5o2qUfAhTaug72hmL7MxharI6L3xpQkCPtM937306Hvw+f0B0L1ldZ191HzJ
JJMB9ZTP5wiF94VaxRg4DCjs8++J8n7iKPrklvFzLEWlv710r/ddiY9VmIkFP9cXswmUpJegb7d/
4xnnyEjG54KYCCp/1VUlw8UKZeL7FHB6GUgZL9mMbvrHoMamPXqybhW+/An9Lejk5BxCOW/0fw22
I/ksP4OoYEsKdBUe4M/Z4u7WIHfsGlyi/4ZR0N7mI/0s06BJMUoIW6Bovh/d5HmA4HWfKmBHm2Yl
U3HZmbfHGVcOs1OR9kVDFMJjKI4RaKf+54zN4+DlW3sxbCJ6V78J6zWkjUOTrwYrFl4yBjIZF2pK
PxVHWQanMoKVR+jkUiyy9kTU8eVFHEKKlNaRxEctoI3APbnDaW9EpEYcteTuDx6wBMOh7KMt05QQ
et6znEyOyA6o1bTVlqruXggA+UkUQEYsEqi5Jlryv+zpuPn5Ec4SM3dtHsQo3MbZcbbnmrrMNtqQ
Kyk0ObrEF4Jt2t/Li9Iah7bB7AQk09YmkasTGZ+Q29D9v/MzOOx/DCThlewaZcm1W/yqEAxpU3+B
g3S9EgN6AW+KABSxZsIwjySRWoa1GeYhdd8mG3Ol8mo9GAG36QMNgy7zPZAeRnM067icMQDRIqOt
DvtRu5NFRZjDMFZht9H8KbLX7eupvpd02XervIqb+RzwG6vd7AEEM7UbWILE9usHXxlFAe24qs7i
ZE33OqLyQ1F+YOFXR8rxOBMuNhNsb2gB60R5lZ8ojedqI5oq/aUn7k5uVQLhf1fYiDNaN6Qy+DVc
BIgLhrDAEVS7ZTILgsQr2YsgsrxEmBUYjiEwpvb/a6sQFSn6njieoy9U6XOUGddRFdHmhohuaakK
4Tx+bnbJwc683EKFRGcvSwbxPnxhueqgU5hqXdL5XVQFdcYYdjJL7txOrRwcA1nRyc0eodbL4RoA
MCG2YFx5fgo6fUxOikdllDFqpX7hoAOJFYd+TMVwtMvsb0vuqsPM5m+cOvu1l3T5nz+YaoJBYcAY
DwzdUEItwVeO1Q7kW2/KxxLHo7IpUCOtY8mezVrk2MigxloREwTRYOs4P9yMP4KNLM8V+lmxiYIL
MFv8JtmS1pyPPKHuwrDB4170u5PWC5KqHMKslrtgceB2Qjn/ZvTivU8FqxRE9qcdoPYGxR5ZTdFq
1sdc9bN+KrWM3RWSOo6UmkDgZGCLyVOjLNJ4SaMWZJc29s3VXCghOZABaH7c/ISlgIFQkRfvuEsQ
AQE55OcfAkhv+iTgMJZRROuXvdkx7Eio+KQK1ahEDKpW5iWf124KpnRfI9ssBmM9q2QYfzSf+TnJ
5aQpV603WYoauEHgV7pKzDSkI6LXVYC8zBS1J3ANv7byA2Gy53U4Al23HJ+F/13j0imJpaZW0brf
g5GlvKErAYhKvJD/02CiCE7HjBhGbDZUGkhWN5MxO2yyrjiDzQjx4uXjd7fK3pVsBzPdIb8i+LKJ
KExYgDDRCf5Wa2R3ro2/1OJ6kKiTym6Lh8RqWr3nvNt/7zB2VAiHf2DkCHIVBkdJ6jFNZXfbr2oI
9KsqgFkeYh/an1C86LNmJfB8MFEODQWfXx9jvLCs7v5b8ZLbTfCx4H40bVuxDs9bYXt5a7/OPGVu
21/fZJYebwb7T1/bb9cUVtVysUMgX6RuJFpw9hzIf9vzck4gLDVW51iNKGt8L75TpWZVu1E93hTY
ID6TfUoEmgywYFc/ZSIakKXN68HvalrMYkKBwPCu2w//Sn82Fqp8zZHdOKTk3JKLIjZfJVhVCBym
EdqeSrFxFn3Cyf5+fHtG5J1lQL5ARbDA8P6E5wU4HeOVL+GReKXXdZF8Ovvz4VOitBbRsJmm2qgg
usV2TPs+amJVuiFfSCZNr1Qvxl1L2bKOsqF3hZshVEXiBeEFJ5NiK4fbKU0kmFd7/ZqMASu6Qv3Y
aWVR0vIrh9LHdXxeijKzh9fROp9m7W1eAfjiUzE1BJisPcDX2lmPNVqHlToVPHaYur2anpucW5QO
Oa8wy2jb4r3IRIRCV7GbsO9XA6/K26Q3uLKhE4ljnBFrxmTv7PJYSA5xWDVd/YkMjQbVvvk3ItC0
UFFsTc3PV49TqKFzI/stXp+d6eEIyHCSbXOCbmOPdVinI4Rb1aeyJLchzuI/FlpOC5qQPKeQY5LK
Wolc/yuiRrFiV5lHZWx/UrEurDN/+nE6f9XRFB7yEBDKqlpKlrUCzSnM+j+Rkmft5VDEmEoNVRlV
UgxWF2t+RZXLsDtU7VZxiK75Ou4mZA3YfdK6kXieIQa3zh1dK0evCFG7j4nNZRpxBl/bqNyMEoEq
6WwMpvtLsb77/x3fu6Ew+f9F3ab3K395JVF0EXNz62O7rvOyF3LWMrvpBQkZF0pM3512Hfzv0CJg
EggxhTNdynLBbOogjDLK5e1Zjp1/WKrFYrmGR4YB/Oz9O0Ync4AMJece4nZ9dYE2R8Y/8dS+wGs1
97uQVQxj/9hC2nv3nE+wFqHRMuXHJX8coUjDQtEds+mr3XvzTLuNpyprqcrA9g5OJUeA2MbVGr+0
gCpXf+MY1dUz69ryWPj3pUOVVVaadD9zCeRTuBoi54gqkMSxzgX38ePHac1cYbU5UnaD2usyaHtX
cizZTHTSMFCCysfDM+ulzzyc4s5meVgnPRTB5jkj0jvQSJA3yt/8D7HT6zhykq8bbjXzCt4VXMWg
vZ7ZiuWnsXfatcjjN7omoFijAUsPGnS1P148tpshAVAdWCUrFwtIXXGNYkXMKc3gxY23tIFhU9nH
y9hfmb7RKC38Qr5VjsRFbOFg+kVIdwcnyYkCOPlveNiSHa0PrDRHDjHKuvlpgGrW5jymal++ncSi
6qHJ50F8PMFBflb1Yrpi/IhzJknknPtbmyrcVEkbpDpz7Ndprok/qwyejxehUkoFWbv/h1ne+I+N
HMPNVE1X9NpbsjlDosfWizTEq8rRBnC/hvUUT7q1hXu+zacMv4PgmjUPB/hQWIHnl0A96HFo4VPo
JOfuZGq6C4qiYWiRXNinaO04x3giS/4PRVxWCdDqPtAJRB48qqdf3zk0B8lZlNt/SZVml1wnEaXB
jJ8j4evIlV2odwGhN/JcJhMUH5MplLQZkH4L1L80gI3ZQGKYbv3w8T0cIZfLPncfJ7za+W0Nn67+
dJ48iWSVZMRF8VvoDYXVLQzcJoKkKJFPBc04D6C7g12qlcJdsP1n8kHHL0tyD7rMQiA5awYjiNjx
ssr8pVaGZz+0ydZKyMc0hCmSaLP+4ZUARcXD00qNVtpQBwaa0ZTScfcGHu9xlO/O13/A+PTbdJED
e3czq5t86WtV3sOwPiCQ5UR86aePHymN2YQlSS1mKeiusBD+ygzT+gchHVRBhnAzci5r/ooFCJvE
naBJI0a/1BuTf3lIqfqx2IH+jr5kgDJJZrKD7uLmec7ypr8akqNk/JEdLSApqUlevB2tWY9xZpD3
gjpHmzcl0kFp0EJoQhCZhzhJ0DmNnq0MdBGDsWi5FhWhXvonrKP27LkQTEeeLZEWCQyCdAuVqghD
C6hXkjxWztq2O4sBWR4UutYrNNlXNM0qi9HrcnRHTXVzXmkm0/yLpUUvBEkSRMrm2cevEnOPBno7
3xpSv1ko9ERJiKoAvzTbn5qpGC6mgrZ6v+Hxh/48E8Zg77eGQdqoAC000J+o0ZFyZEivf99Nm9Ye
y2BoL5qzfZ99vbAtAVncLGZ4wdoozPKBqatBXaAnllH0Vu800XUBBCPmEY3br+UQzxGapBpXH+Mq
KHchMUlKuMP4EXlVqqdaIvxUh9a9S/yoVpLztkOOowElC4UdVetwjPQ6Xg0ugxAWoxUCwJvBZGMc
rwH52HSPaQaoYzxaD4sw0+Z39qB8Azc+v222CVIPS63PLxct/CCDTf5Yjrp6mg23r3TK5kBIwQ6/
3/vh2gEI1HvsEcVhrD2onfKJFPn17fLAj5PAdkLHOgBBEqaRtipiJj0pNsyeZZvXhPVrJj8PQ2eF
u9nQv5Vu1Z2pcxA51308rHVk367GnVRm05FKj06g+LbrQUclJMDsY0P3uqo7RSQHPjUx7QKN3e7z
lX4f6px+o4X4eIo3Jn2kBgS8zs8gzIkJ5I50VSQrFQjvwZSQPPHUNBtuFwegzJQbo8QUAFiHJasF
HUE6cJ0zcGrvw4TkC/BttF0+xwkb7HX2+s489TtxSWMmOu8CkH+2FYmOjXYg+5GndjAllpikGHe7
1xS3LZ1eGGNhl+83G6u0C5Mx8+5eirKCSxGDA6YSkB4ZPM6MgY9yQtJmN5IkhswRioWpikmkvo+m
dOvxc2fXDHk7HY9FljmPm6AjpawCbCesu10kd8hIFLmrpHdS6A0+cKHoYPQUaKtBFJUi8ex2yoex
Gd+cjHxKoLPA1PNrDT0017OL1HxnlsE2ibFr+2X2JeaxRnVSCM8/8ZcyJcH2zbvZ8Gff+WZ2vslZ
E+WJktFmW2iM2SoS/xDiaHI1D/Qz7wcb82kIaP72uKAqZ4GTrskSMZ9HVkcxV5n0pwqkt+FVQBdR
gqzkm1hCXsAFvN0aFbPx6OWVS/eTQcOXOCmoqS8coeG9FpER+PP438EN8d+RUGOA+2IultZTfU/P
szWM2wkh3Y9U4kWKErM6evZb6IvXjzS+gk+QiQR2gjN3J3ZmltSQdtsVoIZUxP6cvhn9a+0HXM6K
lhEH7DStkWECD0j0pAhQX8xNQGjQa+6UOOiSiCLHvYdTpeMDYlzxYDLlga5sXV0SpILZfj6dgJxb
ZXxSN5YAZVJmNGkaDCc0jTuZVqYc7B0hr5WXIP71f/ziiqlYLByyUW4eM2uX9Tw+ixsF53E7y+XP
FT8b/RgKayrDVrLCkNGxxdOSSvRvwTPuwRQvvKmh0DkF9zYcKtW93ySNdTpY0ffQu1fDcJsxkmWS
ZI7uQgv51BJROfoIre9FPF9HegY5+Vb/YXzdbuP4LgV9TvyyMyz/NR3o1PzbXa5mtzxSxbmoQVNH
2XQS5tovHDZDbuUmj9uA6DJrq9GnbTbBhhJxgNB+zto4fe7iJmQCSgjC+iO7ni3WDnfvDONxD+DR
i7t7j21d4l9OTMbrR+JGh1rZnpaooEzXHPqv1gyTX3x2dRPhXWtR3MB43lsdt3tsn7KoEet6V20g
cJAg3domQNe2N8F1P64xFkDvkDNgw0qDn0QM+ddBhuNvLwjhNl8/ArPl/qNT4zKJKyxy+c5rMCwZ
3/LNMsiB+ked/LshNMXb7F5RtuBxRNTjA22O6H6VB8T23asep4rncRapU6xddOmhGo/jkt6QgchY
CTw1rHrksz1s6HTvO5ECNiJQuOvQHD69JXLfRXRk33Yr/H14WXirgHp5/knV0FkLbacX3jG4Dk+k
fCPOSW5H21C0s9gKIcnJbDAKDvtqwa2+UUntFnKbsxNzFx45uvqGvqcmC2ndxtefkhqS3zCL7tAs
AVCz54FiSw4JyPqRxUktA2gAnKsnnT46kIoOMMGepke2zkD5EPlNIaFQEfORUcdK4OdUSxj9bOJT
pbnzXBRhoFamSFgTq1JVf9uCMubGDTkT6q/WzFB/HT+CpkBbX0U7Exm24ESJGCL2CXblOx98ZaKW
YkHpkJwpJEo2baqsqUk7rZmWmnnHkYE4YX39cZyQs9x7lUHxQ1zmWaqhg+nr6PElcNSg7qKv7P6X
4u/fu2nF+IjoBbRuA7rjY7PlIJuqLTqIRoi2skfHN+JPQfTCB1QwTaKG/McsUmDTNjoX6P/WESsC
QiYIcwchsnUcA/5cWEVBylKUZEje8G2STVWiilJ2cpgAOzTuKjuzjQxES68s5bG/+MT5TMiel+c+
yHRYUIePa60XUvXxOL5589DqLPCwmDqTNTNQDMEtSGxyADtDbOWlzyzUsbzQoZwxaMGW/msGw/w0
ZvevRRApIuXExtQBRivK2nuv0GIUpBa7nMDVm9PTzko0vES64jbgVPGeaVy8fULRyNRSF+o6cQFi
J0K7EkLKRsCPbYoTKGbKnnY+GxXNrzWTjyHBWlDEmv59OXfAkds86Y+ixGsT+W5xkdTSCR/+VcP1
6U84By7jknUX4gN/+MrDFhEAcnliKdoV44she78x0UfRvpq0t8UEqKH/gsm3tQNN6a8F8aylONxB
JPjBzqNXVpZP70sCAiDJ/p61qcDWcmQaJ06XAsNYHXj3RhM0BszP51/kt+gfZ74E3LXmFtFeupN2
4njIcQ7QF+v8YFRm1BEDL5hVpqejcWgB7dbR8aCVgnOEkaFYUbzmTtKzet0LDTfSpFw2t3It/1eZ
VUyppx8nn5gqspua0LqFnRaUjW5gCprSjxK94xPS0cLtA+AWHhRrYoN8965Lcowf2WJkftCotK5C
Eibv6CB6ooIRuZfs+weeuesmO3YYnlNWyENqph2TbEblZSe/jaGvSTtaKJGJjzBa0VF+++cIM5dT
Dy0EGrfYA7HBAWGPUKnB+SU4JoVCpyFHihngUXM2G+qfrhIABizD7FHqxxHWrxT2S4oA8s3xtFTl
6T3g1UQ065CNLyM/PtxQbd2zkA+4GR/6uvUe2PDTLyvEedZYHnuv9x+/SCzJ07/llxXh9BjdSH6f
PuFCjWvWNeY6/xskl0sP3EhQ0X4SVkkP9/FbBageaoBWkESAY+MhsYJjiIqBvIsGK95FelLXeViB
OARbdtPnDnLaHJxYTGiMY85r8rmoHPzsYNGoxAtuYoMye1PPDI3Xzdm1d1JtKa+viIch/cK4/kJK
c5cEKKkPgH597ichF7wTgMQIJJXE4M5B36izEODPwD098/a/bDDSY/ItArB0kCzlqwVX/YTrDzQh
dVTDHHwPGTdOD8upwdE/7Hr6WHz8yLTUnNLbqxB0U7yuNHgRUm7aWkCy04AUeLCewglRZ2byPqwG
QlOD2PNtr5Z/myg1deQntTMuAhB82BffiYTqc5zIkGQAyhfaXXMsNF2+ezPIIkZNE/TryemwZoF+
8z/8M0vwiQwx35S4PLIvvjTZVXdc6aCLoJIc37H+WlM7xpAUIqTrlp7QDasgYwGE7jlFWCASSUdt
Q8bwll/fmhIZliP0PPv0CPdLpgHyXk6PpU85UIsX3k2GNNq/4RVQBVU3iPDt8BRBaqqSK6LK75Hb
58fDWA0/eWkmZ0DdQBMF/dUkjNm8FkGBMZd1SRkPxEArYjag4jBb8thSAge251Pp5fBguYwLGFX0
8iqsC+QAzxlt1R9ei8fQyT1TUGV+bS4Mj7I4q74djYC024W4gXPbv/ye+Z6sxEmy8dSkmXYyNBR5
NKgOiKa7FZ5XJgfQlzeKz1jLeg6n8ljgPj7e7L7VhopbcujT0nmtBxhuWaatKHVT4+TRsOyxYlHl
wkTmfg4wjy7OkVgxcHNYXyN6XPoIqNWAhfG4xop7y+Dbd4FkP4QUxRlKIudBo3KvtOyxFzDG/pgT
kQkXkyD4Vk4PJB5DjdwX07I/1vLpDryG4AtutisTe/YssO0FGv6H2a9vKS+PMtF8+B9RDvJ/EHZ7
kaVMnFn7Sj3Dv4tVI+CXTbxNrjSuZJwQvg49352R+k6yPoCgRzLaXm+aaoW/PSr9NMmRnFf5LS9Q
igSThLnDirRu92qkxNxyIpxT4fGUS1tJg05yY3kN7sTr2OOCL7dzSrEe5EBTtMriwArC92GaCJal
eK19y9ZWR2ItwNS+zTQCXDwlgmadDdq5d4Tf8Rp//BTPQErzGpfZkYsynQgIZnWOY0ZNoJOYzpfm
h1CGMShJWYWQB1kWaGgnH4fBfGshOqcuiRMVdrCcKIFqS6HKCl4WAreVu3b9b04HVu2zhJxzx5n8
TFbM8HB0zp/6ICYnnY14iQEPZNBB3diVPAIvzmBLqyChQULI6j9IrqcK3RYK8JYJ5ftDyJfdnZ6a
oOCD36jJsO8/x+lV3hcbHL7d5GFpeBue+MmB7psDhRAT4yFeX9sbWET4buu9iiUb/E8urSrqrfqJ
mjkEVVjDRyBSkW6UBiU7HkbQ5Ilf2mYlCKOgwmAeIZncREBSv7PhRvJt9wA6s5jXgtNbgcA8g+Pz
N8M88dfja++rEMXPBscxGjsOAjhOJzmP+/ylUDPopS/0XraI1h/n88qCQW/qoXvSUb0Z/Bjowwvj
QAL/pCTe53pXHbX/iN5b+pfzK24C+wC/aIyYqvaopVhaVVh1XA+YdETqySwTAihBbApI3WeLQUao
OGhjISujiSvZHI3U66eaQcPS7aKyqtM1O8BwAKkuUP/OkEC8mjuinAYKowREqYoqa/BeSRwZkatZ
zSy0kTUkcCquf243lyIqrqT1sy9Vov0fdYfF27ymzAuxdTHKc8gta8VSNVTiUwoSCwk1lAGw8LFn
1zU2LzfUG0axDH4IeWY+Sytb6d9Py4fOv0MXGPC3J45INJYS+N+7KciefzVQPFYpmRPgwU62m7L3
earaN3uiElkja3bVBMAVic0xCuj0b2Q3LL+2ZIrapJt228pXHyJe5gocj8C3RJ4yRja9PV8RQ/Bj
P6W6TEJCUsU823NKnzVfKqD871jhLW7KBPUjkoZnuqzOpnwx0D9nMy2fB6gSbyt1NfncNsh4tfP9
XMkiLGLvT1tb63HOwBelDN4xtTCz/xHy3sSJNTIA0tnPFbvR46Xz6XqxrvrQ5pHuyLafpJjBfa3/
QukwM+lSUnnD4NR2tdxifC5BIqaXwD0QTI0aRGvd58zrB2JrRCps5492pnXiURB2/AF5plyeJc54
fKmExBy10i9PAP9ZOBVmolLNPLN130x1beQAHX+cuI2iRLwHziFFG/GPynUHWqOJbYg+gZkURKed
WDHBsmBem4uVQ7/rzSY63uW7W1aoW8aQJvvbubcdlWbkFDNdp0ZGu9CwbGwrOGJpqZxWuBCc2lqI
N1+cexGI6PFTAHzrXe7P4hSLgWqK/qLn9rUJ/rkkjXPHGYf/uzuDf5VsSk0+Vg8GYEzbbHa0cdVp
0gkq82Tht/mXMOCy8dEAsQPQL1G/KmcYSw0LvdUOfcIz4x4eUkAa0isN0wT3gOVw3vv97lEU7T0i
Y4emVRBKQuJ5M7znjrCQn30Qunc8ZjMAx+HA0fSIGtjxgemMfosi466kQMq7iYB0iPBP6ZB7Jtza
NmYPvK7nTUNBto67gjrjpcBvXmOYljk72dPdjZQRdKlXSD93ey4vZRW/4Mucq4GtKtEYDq4mteX4
8tansNgDpKO2uezMDSswqVpuvYrpKfwqTxpMALHGHaynyON9BNqNAiU6v2B+IRv+HGLZpNRSZwt2
xb1H0g2PB3zM4tRvaRVOho/gYl76GuPwcj/Cj746iOmCB74TyKJTn3vTWeiMtuTpRAc4e7OGrpwk
zYnsIDpluefOs/nkR/+HNw/Mwv2T3dosvRdhuO7taWzHYbU3e4z1A9XECy+6BI/WvtmT5un99qvP
wBay4FBSYID/6hZp3PpI5L2ZuEq8OiSNmVgsRbkqI9djpXg96LFHLGyR/KrFpzzb9VIZXH0KFaCQ
8AbFNa5+GY3eCtDFsiQTaKxWAnhwTT0P9r0KUsREf92PLPcj0iYiHgeG3x+ORditfGUVTTZPz2of
T7MZrzRr9s8Tib3Cjbpx13qpqJMiZrpKESuTeHYAcPMLzDCBeoAK79xJBc/kW9HIvPE8Rfkc1iWf
mUcEFMHsPDQ++x5kv0ao4mEb/AxI7B6vYNPXngtn1iQLGW4GnDigzQRcJSn4fYYabxdyDCpYcs5W
7pm/q0iIY3CeAvW2hTgXiaCz2RiqFIg0lxPpX6NDhmQutXwTDgOz0+5l6pRXADGnYBggUE2EO9E1
9IX/u6U00y6Hj3IH2CpC8eydP9e21MkVRCpUCB8+TOGxnloKT27aNIB9apJEtgAPPV/+/ISiw2jA
md8wMLe9GIGF1/1/pLU4/jLKwYpofTTPXNOBrrJ9DMkKqDDuKo5GUQeUnoewG07OWC8Tn9U5rzzF
ddVlCVuS7ZeCMTprvRvymdeYf4W9mlIDCqITBcoaVEXbAVd5BApD5JZVW9NK/6NgWmyduO1OzuOX
OtoFHJy3qh1E2t+cbWQwPrcgInJKhjqZ0fPbNz1C/QZRfE81hE6qFLURqTbbYQe4X41o6k9Blxki
KFhQQlFTNi509k+Z/CWyMwCkWRB0+88Yg8w947h04TjF3smeIP/WCBgDh/t7NHhLHOspuLRUGULT
NyVTiziyJ9bhVCn5XdZr0lnMhyLdilecs6EPtf9Z9qACWAYxrdsQmvafyiB7a1FWBZnJa8W+xPsW
BB/bOAfnItDR8iAiMJF7nEiCx/wjvttOMFavjJRgSDSH0XgsNSlRJPr0DdXTpE+lGb+Raew4x4ZW
s3/VnQPLxJq7Udfemz8iEyG3hR1dyCJ/HX7k8gyUxaQAoBOJsf5Lr/l+kuttusZYLHg9CtE/Wi35
+4bJU6rNnfp0od9osrhGUEAg63N/FbXACvY3FYvTC6SWgE9ubGMPTlfqDxfSJwjYjv1MZO9I4HQj
0Ze+TPN0pKeIBm5SMU5VUd6+fRxQutrlIP4YtlRGeTMyDwug8TV89/o84gi6iA0BRom4DQKkDtry
qErSfl2DdXjEx+AzE+T7OqA+2dyQM3FZVPhp8QAmCUlJvyJYoSuQbJ7Bmv2KVD6h9nh8LLXx84pq
4UFyXiIK3AL5DtQGfpRcnadUgJiB7b/ugNw7MdfPayQzpjG5ctEEmqqJn5koYcEaj2l6bxyXRZfG
5tbOPyBhBGx9WShNJC+wzRN8VMOGE2D9f/JPFHZw65CTMhlba6vw7DJuW9knr21IjVUBJWtlEa6M
2d/LisWu1mJctGOUBhwt4YOnLdjF8qMaEQ5ekTxjtboamyvBUkJ04V04IJ5RhGdXDRToDQ22QCXz
RqVPSThUMG47Eb45WE3ykI8BBgckDmE50VhZ6XRVcKeabd2tfA7umAsS3N1RHWU3Ijoh26l6H8tL
n4MuC5w0tJcOTf9wrJ86R9LSdfdrJUNHPHRZpGnwj2yKj0BwAAvDs7eCVGDerhaXfkLB4FNBkK67
FM7yVSfSizAewaG1sp8K2K4VA0JdOWVcq8Qntd3fk6INjphNpU863biTNBzIwU76gfeMRDg+d8FP
eDcekDI40oPs+MF4euuRGEVqqbx3yOqtkcO2lulY8qiIdw3pBZCWD9jxq4QRRD4P6yFOcUmz4b4p
QVTwHmHuEUyeNYzerUTAY8qa3cWh/iZL+CE/nJK4RBdAoQMlWnrt370EHL6pnaCIiDSdUx+oszPk
6cuQcuWIahF7GOALq6tADLFH1xDdOJ+fSUPehxiOTMl/KHsCgmLe2pcPNPcYqKdFS2DlJ7GwuV7i
w7IEqQTuBXM9QcPdJSB8sPTuqbsMycnIUyakPuXUNzMuQ++4lqvElu4kfYb+Sfz/dkZrCvsxrEtv
XHT4+2tOik8kDm191kpp6meA2WHWkcloIHP70uprM+o/6Lv60vMrDuuChg2PKfAHzuGicUsGgg4C
iMb09z9odmW2/T0luK2Ytn7hStmLXArbdkhuaMAYpYmdWcvfOMRZgq7k/bFV65cVbH6nRKT5rTUo
Z8gaHzhyD6nPtE2IE8pKBgfcnybCY1urFAiZs3E8Z5U0zvbrOqRaZyZ0GoYypqE6P3YDtJBxpsu0
eU49tYksU6zVoVV7l9LWdTm+5WkElI99fWOkDPZ6ZMFSENO2oiT9ZAsc6mcxOy4l3b4GVfPj9CDt
g4ptvakUpRgw7ntKrHQB68AecyOq6gstiMxMOs719cCXQIZDqcphWXr4s26v7ifwPJTTvIKRJT8a
QUOtxYXA4W/oHJD+SYSqCPE3HSB2bvUi+2d00CFIvFw8vvf2ZFBcJyv7xBBwOiaOwPtng/GvaQuS
DpJtoF7pgCKmwR9TaUb4iYX08JjWeW3KFMxL+30uOQG5CHAIIMyPC/dmFQ9lh3HZ/ue6T4AA71Iz
kbvDJ/KDShsXqXRGcp0tFH0RqiLI9vnMIUT4P0lVl1Qm4JmmeUEk7+K2YiT1QrOsDUD4xnLQ3zs5
Zg+q3EM+J1KrssLCO0mKdH6OZy4v010rVhQ54EkqAh9Irl3q6cUtRzHdC0/dXbrAAXvgk9IDIgqg
xu417du/IFi6JoFCQFnlZ1hrphU8vfeqKCSAxTwce3tvB3mhD5wlf2fNPz464afJ3rGVtO2BZuVr
8A4TbI6np93jLsC3pU3QQZMXyFKT7BLsf/5L+VnJ56H7ms2DaguxFG09OtNowkFiaKPcp5eLBTfy
mCxC59iaPvTwA9OVz7bsI9jzLfGbNXfrI3+qAWCEKvkhytu31Hbc4ChMrpP4IuRsV631RoW1GGh/
IhuFvgGIKCZxuATa9RYiP7/agMZurEiSsLZlHQQlg31RoVQf8lGrIH9o35CIg+ILQVu/ZSHu1AL2
QOgEqdjFNUJ22I1yUkm0e23BZiKasiPgsYXJSmpv4PKdahtKBNCrMhHWv6+O5SQzb2MjWRQqBhqH
Tsi6L7KuNWeVDqVb53dMq5qVNCuYIO8ZkdHMW4O72EZC9FVHDH5jhqAZysWrPHlvd4dRC2rBvAHd
CK5IcjAJRvl8Z0keO0H+VfBfqtzrgGA0vaOHmK+UpUf0lLDol2SeyolcufiBtKntkt5YFKBt/C7m
L1zx9LlQwqhUhmHeO8r8EkVaMrhYz6SRIAqVTpbCBJdQmmf2chowaeph9QgrDQwejaZ33GgQXWY3
PjDX0MoWzl/soE+3AF7+eb8uxlLgWtFsYZZz+FhCLHn4+mWSbRDKainf29ky8lehIgeA0PUkQXz6
29WBMd3AxVxJ5b1seqbzSSmbJFB8/oEF1vi3JzmJo5GXHFwgXSNI366oiIUwlqMyCw5jSqF1YN1p
LDubsxDn+SwJKTLZ294SxEU/9dvtexWn4CRhP4ghqL6yOjSCWqgo2uVaBiM8THZl1fj25fmzARhd
WgsYb85SRRWSRblrNKVkdjASwyGx/1xM6opLTC87yQviGtDXrrD5z2jmMgfjoCX6DvA1TpnVshsK
pSOhNZ3BpTSzyLZEmOpqBh8qEGUtcxY/Iy5SoJSZKn2q4/Vt0h3ZmAKOoYrVFSvyAy96nUjk0vjP
Fj6c6/uorjRTnqGI7RbbyEM0IcqtyL/WftfspRPhlfCT5oDuZRWuTcxtTpvmY2YVGvX0Cfz1C7fR
7RwgaS9H4Ivag4G2rrcBO5iTBWYT75AsEQGh+0bKgPJqE6GVXJnVGZfvQKScNa8KjTat3mLQLUNP
HvpovbPsDHIG/rohx2PoIWT5H3Z7F6Z4rovAq23el7RMqUseFZyhlqLBttuMhy/6QJ+8OcBrb1Lg
ji3zdg67b8rbLsxk8k7kGx7Np7g8VK/Lhojo6PJFdtYly7gRjjvUH+58rcNPsYSlx0L/qqfw7wVC
BQFliGXgVglKVqz6M1A+pHUSzfpgD3qCPNRQhGjDF3WQ00rjQtyLlOl4WSf0zLW+X+Kpn84VTyeq
X6HqKm4uVDhBUB2qfrSUfI8yxC86opd63eJ58dHHMnKcXe+hcp0kTn92eWTFUQOwbUztQPT7Z1vy
lGNlKgpPuxSXUvWdGWMWtkeiS6LzlsTwXDXcwmFjEpay02yYiGEby3Rwe/fcGwhQMY17NeNiD46g
ZO/61MHlvGgFkr0JqESRqCnkiHl09VbX0tbNuS4Iy/TBMl23Lt6WTnNQTk54pVJC+djnswOfF6Cs
8QGoXOMuv+jEE0rqYQo2S1D7DQT4FLi8utp5QJw3P9/1C6NG4doinrEjHKRrvHgvF67YEwJHSfoE
/i2JSy+5u0mFbbxVNDSYRHmbpCPvXTf4VflvWqIkrH1deldK7WcVnJDuPbdUGDPWqn3t+KmuyIMk
+IHIxhagP025K//nkIwgbC1FWffeY1rUDgZjjB41CywNMrMcROUBuxQDAOsuzUxMzIh4jA0BYkyG
1DZvs78OhMWkt2zTxYQCLtsLxHVlFoWi1EBiTqu6dRdApmfDfq/fhqlrKBWMLSPKj/INdJLFLJhu
a1sSUsnkX5M9f9OxJE+PRI2EAqzqbaWsBDXeY8DCm/Y8kykem3VCHMlujbQ+RPRgz9VCg4vsoPd2
QUGZhypZBgALkSkwrWObinM5QLJV94QILYV8bi4Rjesbcf/n7RB94qvIe0Wpq5WW2m1cUshuSiU4
gYcbPg3Q6KFgSIdZ0DlXJRFWiJG5iWKuTFOItgSHuVlXNAQSKO8JWXhCI9tSj5wplvy3rvT/vkWB
S+83MTwsXpJ5k5vYPp3asKiE5wfsnzLQcG4sdsw9u9O9495YbIByF6BfdRlxspxypaCjQY7hccgV
r+o/U3hDpzg3E5hGLkT3Q44/JFw9ojt4KN4n77NAvM3AUdz9eg4fw1k/tHhEwaBPR0s918ZLNqM2
cMAdotj6sFleFv6A90c+FCGDW8cEZ8WN43v/mFbEHpzy8kkk7tj2W6WATEaQ91elQlueFQR0R8+4
ska56SGh47qDU/tuxJ1oiQvOcPRIW/Jv0onjZipa3gOM+BVhnPEryoWsBVd/B5LLbwELZFWRcmgx
Mf7sQM1WUZIBeZceNp5j5vwp/8Sqy65S8PRibzAJYh0wjMIhnIIa30YEvLmR7BQFf4JqzOsesSDm
UaV5t/oAOgzeJiAN5CELwFoQ/z/tf6MEjsVEjQKxxA7IJTCQAQMZDbSowRE/ErvIF2kPBJSZG3mN
L13JaArAHhqQeYNldyUhyBUiX2DRhvgrfu/1lpI6QQkXRpVatJPWYWHYMmx3J1cAOP9s4GZ+QEfP
04MYcEb0+YPWN/865DCtkPAOMRvDTprCvQJceQveMfUG6j8Fp1/E7TeMOg8WoEAZd0Jiiub1a6aP
CcTvtMBpOfATs8YPxrp/Vz8kddaWT9KeLsCwT8VPUfDKiP7wRGzTNUzrafrl/c3iH/j1feDoV3QT
GoMgrZp7iWXtKGezVL50VL2gFV9OTblUoosbDbvQ5n3KP0cRehZwqcWF6Ah8wnKaW9n/A6QbEgxp
rJifEzrMos8RlV5wwDswqmNFtKp9gU0WRzZZV8YU9bQRZEFgoyHB5g+EFq2A3Dd0Q3AvVLmXrFdW
IWOa4OaBGpV+lH6+/WEk5X/+f1EC46+Q6ItB1WCufNiaFR9NIZVFlyNa3TItd9cAbquNNX9Pjhoa
3mPLfv4x0uwqVC/qWHlGe8g1yoliaBVjU7JFwo6rsNwRDLofxEsFXmrYMKP/iWKRlKeIYxUaCrfx
6SQp/TGii/48GLeowlxDGS7hxHYAnCyk8yH1SDghi1ScTFdvDkw8pG8F0jwa3ZR8nnzs4u8QnNf3
jdyq4auH2ngbDT4sMcG1Cs9YavO7p5LBzh7+AFkezbv5xaOeM3t6+pLJWdLMnWY67RO601mP+6QR
OFnwTZAKGOeaZlIStflhWzTR0EH6YrvZO9j5K+xZ//eKk9DN/6ZzjfllOcQ1Qu+iA8qJfeTZmDBE
ui4OR9bXWYLXibAg+gTeXNsl7m0JiQDCd+4//wOkBOD2U69XH+4KgDYcpBIZcxrO38oS6JgiTF+g
GvhxPOMKfzOB0UaJQkOxBzDttNaTXhM6lh5pltT1aRw9sy8LqC6x8fK25hGn80RIKEuHDsG0LG9H
1lJ7zkoJNPkaeTItgWED7d9/80EgO6TsD7s7J2D8RFZOeHKN9mBsYf1N/50dVXunaT7FtUS0kRt3
+vhatlcVhq9g1J2+DAM4p+Ld0NKZUFycJeQcquTdxV4OLQuTShBykq2GdF6APE4y2egEf/aIN9H2
KvRYzwgiFAPiQX6vzpHDYlEJBQtUv4JCxrGLWnVcyW6hzhD3AXTOa6JaqSRMH8tY/amtbuGIb6jd
/Eyz7hfbl0JOBS0ulWqzXxARGQCcx5UF/o9QKAor0l2xRH9/9QItIkqG3IRoGI878rm7luoEutDW
ieFRTdhk3Vy1Ki6daxbNRs0jbySz5oGjNiTg8OdbTq11uMGmLxGKURxl+ruTqwzXxAS7Z0kLAF2/
XwijOg8C89fqOkVI/KI5aLk0f3TqJp27WOTyoUhMRdPknih0QSGye6+QQT4hzePC8WtNqUCoQcsF
KpTMeEd+APWI0oggDJmvjkV0R73Z94fW9Yb60icrec43l+463kZ90yObHEciZveuKssdKLDPtMhI
PXN0l9z/b9xAqeXkyVdIe7jmWonKDbQ8+GgWxwOuuxcgeQSmhxUq84a37zNFD+hjmqgtGAzjAKom
AzOithhnZNy+q2TIcaeuKTTin074Dil3tCRLHz9u4jKJReftzkWVtE+tWy0/m9VjHxIl1/pfkxnV
4Izqu5/LdYejBL8Kp+sWXOYjm+PosUz8XPeQAdpIk+tUr6nM2TgmTuO0dhKh1Yb6YWWbrNHdi5Vv
GWTp8v/5tICRTCRrabuK8KipsDkj4WUGyPJD9/EGIr1/desUPCl/inCK6HxKcGsQV2M/Iyrkj04i
vC1mvKT9IeTU4FyGJtSb0sZz7Fj7Spew5dvB1thJWlm7MAhZhP2sGMwt0slhA5w5AvJfY/WD6t3U
rKD6Ar8MZVVmf3iDf6C5jeKRtaOlrW4i8Cr0v/hADGg06LrtEWM+GbDlT5p2w9zyLUQWOu6eCaiW
obp8uLA+9mEjBGr6j9bhGBenMPmDzLfZxOp4OCajiCTLyzF1JsLzpXF+QevyjzEQU3hCrd9NtsmU
Abb5Lo609WdH2ZVHKR4EYyEf6UMAJQd+OREhk4csQhSpmA3df8+zgTvAVy7vyFd1rJGUsrbSMKbR
FEV6S7LwfctvHnQpAQ6W26KzhwAH5Sj4x2GVoIATFio67RlPHDkjuWJ9dI8dv3RYwc53UA/6A3MR
sEvfjY3iHQfdkhTXXk2YUCJBPycZxntJUxQEE9pTSSVzEmeacaOFDzeHKi0++clZorKqMCqS70Ep
z2cAeVhkKxq8NcdV9RjUgeZLFyTg52D8wVSIveVA7XDl4HVkE8kRvryRo9kwdpHYP0W4S/t7rpk9
86G3KTxrJA4J5yn4GoHK+BGjgvPrtjHAxCeR4hBDIl5Gn5COMyD3RCXzQZ3MgbIKMXO7Q8BoPDan
hDzZcNEVwzv/VNXFj5469N8kT63u96b6wJqBe6Vazm1sHRU62QvfNirHlI4a3s5X5EiIFvNV8oP0
CbQ/OGuBoReS0Bcz2PCU9lszUbYdHelj4nnkeUCC9K8GOkueMtarEWA73Zh6U5U7q4peQkwLBmzS
QuzYDQSSH5gb1GPPe7vWCeBMm1mybsr65EGZhWZBoCZdQv2uhcqa1ovcquzCu+f7Sdg7RZAJqdlx
DtGL1qj+a5L7FcOJbadBao7oxsJrO0uv0j9KG54MKuMk4P26jVD4t3Kxv4xlOf7R2n9WXFUvJsO8
KLq+J5XOYIrUKtyZVcICsvhTS55i5G8zzyvcnoGBrv1Gz5v6OtPcQZHuhsIMyuVJa1yJKvwl28DL
0rY4gc+AnWvJ4nxv6aH+nHfTQR4JQZJVg16z4dzm+pkhqAFCFDhYJlxrXNEnbl2GlzBvPjdsPfWk
4pLfuReWeFuPO7tB1YMRYOtfwfqIMuNmDM66Ndxx0+nzc31oOGCTRRCYSvYEoCG4eo43LTm5xg2c
uiWmWAOD7+IfUSnVUQTEC5iyo/lrKF7cRMQhDMLPtwiUJEYZdMVVBsP82Ubv53sukzAHoMdpSWOd
RUTu+kZVh2WgaZmwYvEQoJEEJ3T4+yYhMkUmm+/CNJzeVxui90Wpuz/n6jZ3vqxx4ucORntyZLlk
PjZugNdY/8bq1DM2dWbQDguxCKbYcN5Q7s24n0zJrmm0DKhKArf5T7NjquXrOZEI4eYED/PtqrrS
hjND7Sswqvth3khNUrCMuG8+LqM7xmHW0rJx+De7xXXn/LxuHu2LLxjuBTn7GZ3XA7czbOmGhoPm
a/jwA3dCRr707wla2OIlQ95XC1TQmNs4M95hgEGwl8BzU5DZ7LGUA8f5ZnK8EqPaPpnkIrS1Iyc9
PtrJzsh+QTndY6xJFx0ms0MM/iI8JNI41P5eaJGe8KhFmbvF/YtWi1v6N2lr1+jp8h2+JLyYxcxT
8lRrsBzkoK9VbsaHCLwcD+hZQ+viojLNnxmv2WzeXaf7hHaswUt78oU56IjHk3Ty6+Jcyge4MYIn
CuatvRescp0UH7hBoGsSMYCdz7ExYJA7ddyXuVSexN9YwgNyGXeRiWH2qzeF3R0Xbn1vY2PyWRAo
bgjDPw2/LmZemTmtQxgaelGn/fZHMdVGTvbqvOPKVvsVQqpqFiKbEF6zPX0Po/28QWAaUOCOOr56
S2Dtn0NhI3CDvEYee7K6AAWuUZsnkjkTIUXEEbz5xp7fF/ue+MaAoAR71MUGWhiLIPQXrHI+q/zB
2/IFnjr1UkPJKKyrKcQqBb4ISb3+71ipXEQ3ixGVgSzVu5NIMrMnWPn1BdzRX5vCDo+g4R5PL7Cj
9OwZKtZUf7i5ie/9/0L78gx4l+g5+1j9/p5pKUK+yOiQscN7aU/Y5iFxNdu2TiPUQDCtro/CvK9F
ruskPQynCNlmTHnci4lD837fvwSKSIrAwWXkL9jQRgngeqVAg/onyC48g96EKEm/XaCRZPGAWL0f
0u85HeINvUPdEUX9TAFoqO/2+UF4sI/djemNg2/OdvNSI0MbGj3vuceLvjDOOA2O76Aj8R65NrEg
j/tIyTSQy0YT2a/Pelg3NS9FCD9FLvWJdP5zmeRT43W3Mprle0BnwCaZTFlirC6YimIydjfWTW/q
qGQLg+LYVkjh6XdJXKsQoPRaAJdwzVE4HhH2OQcN9gW/ibVXsoJCfcVbpa5ioswBw+L2N/n0ju2I
lRWeW6W0PRQk0q3NvyYU4xgz/HdjsOoQ9FNXpL2B+sItTVo+bhh0a/Bn/DCI4plvcfOZ1LR1hhKb
/xRbhWXXakPSiR/hfuyp+AdhG4iG+K9plq7wLMp1OEk4DDEbhtUudMhb7nB2CTp3MQ7tHDObw7Rt
CIY2v2U+x3TOZ9KeQOOM9TMk6rjFbqZroUHPqMPT8FDHzlo1Upb/gqExdEgdtvetHC0yk8mcGLK4
Q0SKllXsq6intscMiuNdHrfiEuuAlYm8VmrGkPIsKoFpu00Ie64FZPoSvAhCwcTjSLRYdpFk6i+H
OWFNpawN/sHVFhIannuTwxZCfO4lu7jL3tGPvzQweVTmMXi5ByIOf9345xt7bbMdcuvxr03F85iR
NzgmsduHmXmau5vy1xRxAStk1fnSeJwM633DQp+0GmDqqBgiPA/5kIil84Aoe2dLdaaRm7xeg4jC
+jmY7fANmg9iXhGOx7zbOAAOED9iQ+KIfiYTY1UF7iJYxUmmVWnXV4o+jVUUh1VTXB4ZjHGYro8V
yM4dkhoHiARexTZrwT0mn4meieIm3xqwtsnExdDmGf6ZIylZiG4AXEkr/OmN17LKugukkubVJog+
xmMn+5HKHM66/LS4yd4s/AgsFmaDbc0FfZ5VmbebzlXMBXi4MEvhYRC0KvxhsOdd7VHdWRE/80nu
XyieK8ej39mTVb6CcL9R/nXVTKlyfyWK1N0SfpPPciiSYm9IIsNY+IF96yNv9MsbFOdCBIaRyhjz
lCCzprmwrzFuTj7BUEBfejCTR2Nm8XDxfxF7wLbD9FK74a84tpMm41lEViVKY8NsDjJcadPylZ7z
jyqz5F3k8MVCO0e/53HiHzNtKCgBrl2N+Syk+5e/XU/PLaNWlaspi5vjw/rvNMPtr+93E+JpwIZQ
JGTKTieRTME84wzvEDK685CKi04OTzqQ9CCrDQKcYCrQQrnw5epf62H6NE3fxwrl6BVYu73S6AUT
zCXnq7qRazi6gDT6/Nn1SD71HbnOdvdiIAHJTcKxZEORfA1vOWKCgVzp5OVP8vHEUmAH2aGWd6LS
AjUJVTlDMx4xl3ZpmIPjSyNOfrxLPx1dieX5ghBz6Bv9eVdEOjkyAUsrV4sFIJNINLyJomJ+YO8M
pvuHzC8q0gW3aEn7umUTy7gfVMUV2Ym3WNpgrmonrKcl/rWv//gT4KnOreUBDrgaaJMZP/nvQQWD
Q1yALlAp8+ZDhWyhYeR5vklhb4IKIOUMGcaduX2pYkhuqKcn43z8bexJ0SurV/1Ccar10JCb165C
j5JE3QV7bLnRTQi9SjXRFigbTsRvOyg/MXelwBEcPizD1gZhWIbK9dkEfOL87qmBIBfEB0piYh7a
/d3eOMbH6OWJS5GtC9wKbNAxaZgKJcozWlU40UCIL0+5WhjHXSmgU2krB5WRbfIzsXs/0bgn5up5
a1Q4wbkPVQxqJ49u3LIc30rHaTD7386fnQD0GFh06qarbf0LI25csLSVbc4m1s6O6SH3omfKLmWw
LlDxkO1kHpgdijKK1Vs6UdAAjeDBbIiiw9R2qT7DIBsmN6FW/86FhGRf6odK2uVJDANH6aoPhl7/
g22piWagUuUWmd9MrAEU8H3gG7rsnV0eoPp3BgwK8hCHB3LUyN25gus9Tjd55vskmvhblHB8Kw6V
uNfmb4z7D7tXmwn4cNNKh7qaKISHVSt1j1kWOzp0lmlY1JTjQJ9FuR7P6IFq/EkJ/gdJxu6GbpXi
/GKUrKU/z893SYpbOdftq1KYenBhLAdaJuRaQjEJwxGTw+XNfiDMVmzI7TSuokQxdUzHW3hky52T
K/zncKEep1SPuav0Sb3JxPkMpdROoP1312UH4iVTE7Vq0jDdesCrXtfmapm943viWa2iRQht77sZ
fXE88v2spt+ZxdGE72IaIUZpdb0vCd6ugJdi2utzsg2iDN/3JvAknz2TfMGL5knLQQHuU6N6N5QN
b+6wXL2+FaFq9fSsIe0QOgiOZZwZZmrnftvgslNmvHN/SJz4gXXAospyMaqezKoAPsK7UF1tX/Ec
WocgDQrueqPjX1R+eGe8L2yp6d7sjdD8ZWpZpBjfYnUwuovPpDZjQZFGLfib+QyZATU0pQgpi6aL
lD1FLd8mVZdqlgtYwIe86D8+KjBNTm6e8ooMtwEP2SAsXtVOh92SKS0WMkAXdd/xeuPxFpCkZeuc
ex+KHHFDQsMFHJepQhrzUzS/M3rhtf06IoVlqF9l/DNXKVTaH95+Bg4QeQPFKSmF65I+66bgTQCG
98y61uU+oQhyQWhiGZo3zdhE851dD8wqU7A4tmUM7Te58IKs3ImV+D7gox5aX6x/i+VgEW6r1fcQ
vYzo8c2uSxiC+EMWKwVmvoxcFNHAWDYRBSgajitcV4FOVZoDjqV85E6DmLfR/aAo4u1OJh0OOqaG
XsatLi7CIkCfZ+NqDWyx0twQgnRoGcctBjH1YqKI/2nGTlbGuOV/N96oh1YsxnR8JbKB9sGFH+zN
imwomPwVm9TaY40Jgr9q2haKB0LiGhdYvA2GZ7BTvW2EnHOc5f8/jB+7JyZROkKZK82GwCu7ObVO
Uf1qct/9bAU6QMLPk4GvDFO1dSOI/eV5votcKh3M/NL5UKdEs3DJWDlEH6R4FOgE+VRiVakJmj8e
aCNeDSoqGN8/9qe6TshwjRNFyB4IYRN2nX+oOX25Ge6HOQ51HuD1aWHP69+ufvphLmyBvUzCvJAA
qcM3FGyi4R1/VyHtzvnbkdmFlC9NVyrKDJrDf8kb29nIZQvY3HxqvzpvykDepBu67+dTDk3PTxS3
Lpv/tyuY75w8wfoj5uJsi8phopV2ALLt85fwKDLDQOYX1nHrb86/6ChfoGCYDABNOCkUnXwb8LiG
eS6yzWuN5oORPKOF5kfzRjYZJh8j/5h4xx8tymBWpyuO8XB/9VQfH5Bc0a9qx9XT3rhpktL68h8J
EAkkpudNWq3n756CHCTwzYRfqi7+cjU8pfr0IGdjalli5NdvHrTX/xIVh/v10fkJZoaaCaoON61u
v1F0MArjhol9u6o6dt19deZAQDt3X6DCu2ZJta4X5vpSjz6l2GbOlpDSERKWXbjyheH77VyS7kdZ
Y5OjgDU+my0kWnKACqweMV737aBijpCgxZXW0HZd2NkLRMUdHAgEzwHTiG/nsy/Ak8jaPxODtpEd
YIPAt5EjtfybipA8sVuNIVauFW8drPpsnMzPbqYxJCysrCfWrzySy5Zzh+ZrpD5gzKblviF4LCuw
5Arp5Jz5JuQbW7NqT9RNcQgtxs9ND9PomLfnPRow2A6SdD3ZXS3BhfzvtMtIWI6G2I5JrblppLY4
icDV7wnOHW5M9AUs7az6YC8//XY1xXx6QCmWTEpVypddHUteWzZB+CuM2I4hMSm28sVSlCmVuPRM
gcG6EXFisbkB1XneYDJC8FvcG+1PC909Gv6hJY1Ghmw3zqtjaGHYg+n8g12shmdxDBXephIcnZ35
j01aDjZkLJnngwkDq4eCnwQAaV1fT2UMuPCnpyHKX8w/d7qE4RRhpSY3Z4XPMECCvgcoshL84PHT
agZ73dY9FnP+735v0sBmkqT1B98np6gGQZI5C6mwkxeCNQ6fvdQujkapR3mt5R993X01rfquK/2R
rvqnhJYIU8rit/a+bQMB5mu+bPCZbPTVmbB2207HkTE4izWoD4KQ2oIYxHUGD1F226bkyFYiKyaz
m0kfsnkpztw04VFtuSN0PKJo8ziFxlYcZBafYcd2ijAFp4REY8bO1sTE0PfDE8hvgzedGAjv7HZj
uKZ4iMxi3PxACT1DBbTC81KCAs0PP2nRDmf5FcE3gp1jg5u288tgcxiovcF4FbK4eaAcBmDq/rNm
N9nwGTr1aLpIiWqMzp1061yxLJIPXwTfS6uVPPjXHtgP8uPmZmhxd0X5rZu5sDRuNYzh7p1FkMS9
ibPCcaZVhaAgacB8vfECSxwj8Z+MqFSLqHXLw8IV7X2PNTFnNQ4+HoYuNsY9m0JI8hCs+KHTQBbe
UOTijqWG1zVSnzudIsp+4jHWh3Hv7oiuQqVSeLU4xwKmVAqcW3DXxGQitn1dRTAKRE3DRe1PjCqf
PB2gJteQFL4yHVeKIYhPDJSdjkshRSmTewiluGv3PVddjn/wgKBqHG4S7f+oW5bFQRwdn3/2DgID
eu/Lax4YuzYD27MgtJ71KJ5WYHauiUuMY30sfcHiQfBYtY54+moSL33/EP6QBpc9nYlScXWvJuo4
yI7XkRD9nT/hw59B0vcrqX/srJ+LjaNzXr1T096sMTuq8OQsV1H2nbggZIyojkSLEbm2YjaWVtqw
Qc595FmzpTqi82jywsiKfLvStDoY2p8RrAi0PTkLeThH22zDZw8NNKJ3dWwqBP5Jg0uVv9fEdjWg
VqTLXzF0Mijn9AyIK0oaD20GB23ItTDcA0+64+DYKwKjfoEzkuqgC+w/9FTqBBaL1m81Nk1MQPcx
GNw41hv32yHsh0qeQqP2nDW+3f7dmqUBxgkXiyP0Pm2AJ/c9UvO5oZsh3qXNGkSv2Ka8PoPrrXnF
imxl5qLkfwKItaPbmo4T6vtS9baZmX+yYr4fTd4JsACjKDrtmW+UBy89KCAMlfzZTokN/WJmzKg0
R1nBrlm/+4tudF42ckAMwhuf+o3r+linPI7ewL/S8ZljFty2/Ef0wL8zEHL0BCSlah14G+Citoue
UvzPwKzVmBzEsA2HC4IKt4jpy22ozFzYJ2rd+32uL7KE31kHF1sc+hXGjltMtmJXVCe/nE+plAV9
fHbtTcmSnDeqld8LCQPGuujxE5PiCDBtOfXkwqJLYqlBDUhkKfdCILW3cDVbp+lZG4Usz26/hMv4
RWlnvn581MDSbJmwjNvUztYOprmMf9cA6ANf9fI7YroQQfY3P6A5tM55zngXnw2R4D7uP46892I+
aKmt7ubBvaWGJ15evZjSn+RYxsHshndzuhBLi/tJQl9cI6T4QcEPxU6A8beG36sNqxmpwYOsFWzv
Qcv7g3UrAJsSP4QbgxkowvdwoKcPxARc3rSRqhiQBrTXsg9YjwIrSP6lXEXdk0qJsk7f6sJk9kKV
6JUwavdt/mPyiPyc2P9Ad90FI4R8WDFpePt26RgxOSmEz9rv6cnVELol4xLL7XHVX+OgXbCDZSs/
xWLhVhvB32ShGjPolz0ntob0IzSkUNWIJFS9GOjaXuqAx7NjT1NjrdscLdR6Vy9Pt6MkT91orU5n
xoFO0HX5KIUBF2+HI+kbOcmauZBgPqXr78uoLKhgj2K7LbJgXcxJpRjiX8MAsd6HqSmZY3/KhwFU
65sqlwGeJpXddceRbH0saLo4hQ6111dIigw0TgmRNqsrE4URyP/uS1EqVuhPtbdDfCbMi03+n0Sb
wtY3DfJ77oahvq8m30aPFMs3OezGPAGcQ9rWIhs9RenjlHWGduT+PkclXKT3nyaWcCFv8OlEcM9n
aqd2d40yW5tNE1cu7xCG5wld25dlqMfTwBSu3fBbJKgk2voDPNJ6IIG7dIu3lSWNoP6FvBx3HVWh
LKJxZWrrG6sebcxcgl0SG6j1wlyYO/hb9poqaSVl15tvasoRjQnFwj882amAPQhuwpwP7/86O+tP
GNRBnAhcm5S7W0OXfLLkYpLHk7Ic5JGaT1ueHDXbxT4aQ3sthTtXEDUfh7G0gGB1DsSYXAweaZ0V
ZA7JwQMoMP2wumo2GeRLJYkS1Xaxy0BoOghbTedTHAsJN1wUXA74D5Df3B7Y3SZm9EYRqZ3m20Jj
qDBByQAlQXKE5HIJlOjeBY1lmS1X7xZQaFvZyfBecv6IC9h+t36b9UdAcRUgQj2L+6UYt1gqL5c6
b6er/koFJYfORqiIhO6mu19KnqkSKtJ6e+SM6m/Q8EKUzY5VcFgr6SWwvQxvK1QXyReiFLFxswt+
3TCieQ66bQ9JQ9mZ4MOIy4KrXiZyKKgz4TVJCcbEnR3bvpwBRLHVKg3fjZkrZ5Ow3MFuGo9LwFWa
Ly8C5bKJZsvElTNJgS8gD7YztjPhxDAbYpdDKgd6bx0X7Hw+SJTXUQ7JAh8HmIR64gGJ3aMxkkIg
eLVMw9ZP5Gqu68HuqDrlpKEtwiGiasxquTx0VrxdKw3wh321ZB+X9eGk8nbzCTP55A+7ztdvKtnS
CMU4NGXZUkK6Lh5idC75NU/SQODbtp9DxxFH73UA8UvOtXkrbIjzlbyGhy5Em0DrhEMbMhbtEoT+
g2eimytYKZAUnJeeAI97rIDKqjW2goq1ui69BR/ByZgBIMDlxUlYujN46LQocAV6hDRpnR5KCjnn
q20+brQ9A/+c1bttQi/qjeZrKvkQes656+CKMWmyRKkpAijDaOOKD4x4miWSvkPDCDIBn5s/i9Fe
0P+6/Fu25i77dhCATOEoRhDdSIeeo4eEnzPriVquh4OgBx9J74FFpUML3l6XSPl/Tdj9HMjsNXd1
rq8wCzLHFt8BbxogBiNnBaNupy7jcsTWDDCLN0egJVmnZDfHBKPEZi4I444L8ywQNOGwudnldC3E
QDVgsqunkQkouOuz3RBf7JfPXp59rAbI/PIceJav1Ln9q7ZPXA3t6VCCXs4Z8LSDAdZ5W+gpU8W7
QjMi/oAv9FZS19haG6bA4YuB7/lhoVWptPQloadMuwI/oY+11aTZPFgzyCDMaJxPrlm7lbPuvU6W
g5LxHjYF5he32A4onQ5IcZALMzCjpFlmYi5K+8gjkqvDKzQbmPB8nD4igk7MZ2Voz0RFIvskVAYW
pMrNaS3ZoY7bXURPX2LhvWQvJCuIZ4NnxoMZiaNw0U6s5Ova5xHSgg4Fzc7Iv2GaBpf10++LGo0i
HMpPFdjtY69cYxlg8uluynpupcRPLIKt8fIq1RQeAkHUGAK7CgEwYDFw2Iy9PhXLj0Pd9gei7YhR
XMlvx5N/puG+57g2ygHHD2NteZznA3x6dcUPnqArBtyOfTtMq02mWffQvpUTZIBVPRqO5ucSQCzC
dpp4P0Fvj8+a478MESSvr7sVmOuB+q8zK7e6ynfkbdOHDcsbPjd/48IIssboigLPMpDqLFOU6T8Q
Uyh1HE4U3UplWOirb1e11+OBAWc4r9xC0w3CFjGiO3GEV9JgicnlltlY4KoEVvweC9pgAik9UumW
nWpQEt080N1H8vgFwbQTwE1UPWpSg2tlZin+1z/NVWysY3Z3w+76nX8KqTrz+9fJtrTGthx2k0fc
kO2/vFHJ6TavfIrcM8LFx2NJp4Axx+GVtXOkj/9pG9xmnmxjkNRuVsMBV9vpk+x3dWYdWqqH7j0W
TTBzP5WZvFSECDNmmLDBKCjqEPb5hHLQb9elB6vl4jQvUFNj6JpUQ2BYNz4cEvIRgP4TDX1yYeN1
XM0dIIe6kajQ+Bvq9SPs7PlrEjyPaHcUUpiyGYQok7fD7b8r3EtB+3B1jG/MG1URXFR4BfBHE+mz
jJKKggiQmd3HQ67XKrTUmpjA77uwbDCzy8FMlKw39YfWQSPCfJPNRxCTtPYoR+YTHcwTD53QKNnu
8IU/KxjubPrKlCy5lPhm7WPiUZ/ANWvPhtT4EwFhZtda+Fv1jG5URFLnBCfFQNqmDPtQ7Xfym7fO
qIF0l9g1GvOGCAfyuX+DpfZJZUyb8avoG+9pv4JNNKl8Hu0SNiP4ZMSFgL5JjXraDIbkX0CQy5Va
Bj21WfHNGc815mDTaKWDq0JO2nUbbaFUsxIph+krpeXZDUjLKTxk28/2yyY05Djd17PSgm/1bY07
Md/O01D980i1oFkHYM6X2W3/w1XxUpaFnqXx91dgrqJnsFJEUkwFTXX8yyD7us1wj6hhUATBkw03
Ybk8e8X5aI0/gk3STXpaHfNRLfqPL9jnUuQkYC90NUlJv8oduNJBz4aMfTGzJofULMN6B0EcPJQT
y2gZzL4qPJV7cCuS2X/1OmJpZFS7L/TO5PPUBP7W8w84o8FlTvxXJy6SmfmAVlbRb56zUdYfsRbD
Ut/5ezLFdpm5ZatLiWqzi+xAqlGnfNojVpCEeLZGirl3J5Xyk0ipzIXpEUdl1YkvQ/V0ynlTioQN
uSDOCblkVQbKEMTFHLvyT5TGm5iyFQBbhXIa5GcStXAS/MCVCJLZPISxjdrqjHt46Dkqyl6+bgzU
l3UkAxtb8PzGiSDLl0pNaih64MnLCyvot2HJarV8MTueQQDsA4DPfGkWbKuliRazr4FtYsEvJvaU
4gQM20+kVqvMZotB9N3U6AEXTXU0Mv4rhEY9M9kTQ7FvjJcJ/vDptcAIp6WS47H2If2j/9/9dx3G
7jwFCGsKuoiGwM0HCWqKkHXnIC5nUrep2m52WgMXHyzvG71Uu6P4/5rheDrcSw+3bCM6fVsmwlwS
XN7F+7lNC6AOVfMKF7pFA8O1SNYKd46ZT4Bt5iOkyhSpN3XLYMwnbcZY4IC04LHeSmFBszkEqmve
tOPjzhbQBpIV63/iS985EgFVlXXRNhAZZrjOImHydFaq2+z+BiJkyS8Zcbs40zoi/QqiCzrhcYrK
cg9Brh1FM4MuSN3YPP8l2XDr/vBdlWZwpCxFN+ZQ4s2bffBteows54YPAK5nHT4RRUvN1lQ1vpiD
5rKpOAo9+wZB+BiRRdXZkgVjQtFP2fQIU6ufQ3ApJW3lmJhBk+3Pa5ZjVNtu6jjzaN1TyLXPLZd2
1KLVga9q3mC/tgui56FXyAGPf3qha71VCEuoqB66n0+F0cXzwj1XxFteSmUdg7NkiKJ2uNr6Rtv7
GSOrED9X1VTA9lMKwyk9gzZF0YRN/jUUOqr9+giiRnHjlKHITHEP83eEuDoGOAJQ6a9BWZPM6JH8
b9nWUpeWVqtV2SSNU2Rm1xikDkLMw/b3osBnOA/Qqf+73ULGMetxh2UQfIdgO/LU9I46RMir9X4a
dr8r6br5PkcUWlP0GbfUL0svvICNmsyHDbQHZf5+4xHv5h6I2Jqk3CU9+rk9DZxxOOAjHvHQ/z12
CfWcbZT4bFcL4GQ09OoBcQS5rX66qiXeBRerzO/1nNiXznFtnnSBvxRsm/9SWzyQ+phUWp0tQjSB
eVYJbNlRO0s4qsmzbwtV70PIoWQ6kxVo0jKxZYjL+O8BSCWOV3VLrvkrxtzw44l7tdGGrtH+32vV
iLMJ+gcE67mmgGHMXC4U6iPGQajkDC3IjH+HxcKGI2hlkE3hRANnomWZTr+rtwmCA/IyKiSeJO1K
VijpSVTrvTJX/QSFd6NmavhOZbLGwcJdMc5Jv4xSU+o5Z4eUfTWhnnjckwQ5r3xHO53v5xWZRqMn
QEE21NVKTaC5bLcVz4n+yxRLD8695Q7y6qRytMo+OxaM0+UbXef5NGOQlonmFDZT99nPFTiRKvbX
THV8yXiY8CEDyUCZKtxy7y8MjXnYeYG0pxAWXzGIAD64CdmawNJeduoNlh/axMa5I7N44gJPjARG
MF3GkCeCHtZsRa1W1nd+WnnImMcjBy0inpxfObV5XOtmKcLHqtvvDKKOvXTGVWsbQzRO0hUSgB7l
s13S3EKjGJdlNQD9ZYYLVzryPphW/Q3LbCmnwwQlZxoocFxB43vmJ2prOHgGFAjrRUudtA2SAatE
Kfwfh1BWIcu1OjZB4PjxArRfRAILPVpehmUGaHrLa1qT/lGuVQEDyyRX5nkja4jKcefuoXVPL32K
BAhJJxmVVghSWuSz+2k8MygomBDEw0amvUeBX7WvFvNzTgxYrZafZeHReuA7gD1PxYIomk36IJXb
eb4wIGCmLD2KXDju5WJ4HxlZQMyV4vc9Y8NUVlHjw/HBN1n9XYNGebZPNWGCdGE7Sn5WaQ704Jac
jBtuHpzpZvdqhVHiAbWJ1LMDGtb/1glt0ykf8hULi5ppOOllhiIitKyKRY2o0vOzE2fb2cS9C5IU
rmCXQScIZuKr3lZ9sh37O4xljA58Uzav3DtLJQawmvDWIjln+HJDJCivOAq9qHWRCnL49j55Ev9r
dAx8cY1tamCBeKktXLP+uMZrUbchsmBtnL9mDJWBB9uDd3aYKiSfVyJQ+tyEd0jdDwfGPBcpCQR3
qEH5kjqcFOU4CmmLT/WTvGW4ZGYENFuh8JRbM7/9iNXPDAJf40I3s2UNGgQ7+3OphxF4rWkF0u73
SCVzEQGtuhDMpUjHXGDp8mZhzvRakcvCz6c+p8TqeeKQ8PDmqKPcq11Vx+jYbEDYJUdoq2Pw6SrW
x3YOCYvQUljBunP6ef3GqY4CZbKVkUAkIzcxwEBua+4Hh3PlyEQaXVDNV6ezbS0EAzOennjBIzF8
prXevWTVejK+bdJiksSrp6FyRusPqDZ/j8fsGmB6eRYJFKbId2ZDnIIb1fNfwqHZcT6lxrJTbuFv
8VSq5TeFsgJDarPFvAMwxFm9hc4BYZxPCZrXBtMQe5sErxXzznIFUKX1OVJVkCSiOAb+6JcTA3A3
JMWbmiLwi+gu3XcfC8vhJ1ug7me4xuJOaG1zjbw6yRAFmQMRGC4m6WRNt27zKxKbLKZbE3IYWdfP
pfh3KNmh3E5yLPsO7a91Dt2ei/EYDHI4Tsy6QMPdUpB/a+Ny9VE+osp4FGKBdNIILCtDiyOHyL1O
Gw1LZPfX8cJD8BqE9F5zrYmpY+SsLylCGgextWuI/Phhl/GJHnSSQnXaqbmhRadF+lDEj5kBPeBb
0IStJaK+ziN4ZOfvAc9uC/LqOjPyUIVHDKf6wI54UKkBkuP2cHNowC3L0rh3Mv4C5fLzpH0+vfce
yR69NHbI/j2cGgiCutoeHu786kwG64fg4DmOLzec2IqOFtG+4wdbAAATzv94/GqrbDqFmZKw+Qed
cB1n4SUt2wrtT2OTRdjd5K3sE1mm9mOV0THp0+P8vg1OiDoDwzpI8RPbj2rMiZ3c8gy+3ahbNVSf
ZG6nY7POPNBizhjcztRXljnX8D8AMI5yg0+BszcHsyotpazqxL6hpjXTFh44Q4RKXXgyZ61wvdLc
SKYiMoAacWZ2QLrpkGFLJArmmkAXfv6m/7xezr+eQtVlo/iPwMGhoTEjK84o0hm886zjJtWV34E3
9zvEkq6qa2qjatOHM1c7q9mkxIf9wH0ruflLSyHl6L2zPc/HaDaj745ThGMpq3EHEwNH+18+SQ6X
54dAxzO9oZydNKnRQkutPuz9WhwoKjJJpI3a0oD56GME6rA3bGAZXIhqYsz2dtyCcGZLwxb5syYp
+uoQf7tdyAahDbOcNnOD06mT4PiFjc64f9dpMQfoc5mbfPmonmzRQ8riArspH2SnhpKGJHcPCZNr
pokT19fi+Z5dogjgVZVD+iTghasIbQi076c00dqri3LsSFbQPyx7IKhurPw/T2awAeIXqGDJ+r0y
eF2Eu2sNvntP7pjHQc+8YOWc92tp2nSj4xm0jPu4WPWEjy7vdnYvIFzLm1HNp4CgVZKCv7xFWDwx
j1FSfr8Xksi0B2SGHTErjCnbJPoms7O5Swc70lkhZnMUORNwuxTNDVRMVU+W5c+BlhHHRzJ23LX9
h+CEyHpePhMLveCFNW6guXAnhKfEL38aXHmxFpM0XSSlG9lchHIX68rKfo8xDpbtqNftlAjDN/qe
x47qRdtfolmifjBOKSNvueerpT5sV3m25rptcLBKpUQfVMvQn1/ju++2SxND1SmaBEc0ld0ogm5Y
vkcybaOl1Hg571aAuPPWAkj1uYK/bqDkiGVFxfb+rx43t724/hxVgN21IlUl9c0VJK015WWLXf6o
7D3iS8L/jcivILhgqBCEKiQWXQlb4NQLMKIA0oGHNyzdYV4gTnD/vJWwn5GdFCWUrvhZP2xUQL19
OPv7dTp/qw5rHspuUIzjOBHXgS2nokPqF7nUtFa80qvf1Nvj1fGw2ZaiUPTG7FUA7Q4WnjOLZSmT
u7xXYn3tVXFvoGMdo9LCvqcUghNSsj/pO3S3avqxUUB1knO9alzhqpuJvkNava5rQ7Zxahbszhcr
P1zQFJDWO94uHSeC7uf3mDxyCTIQ2KqQfHejdaxN4GLVlPt7374BF1GVSAJQBQBgdoHJM4yDrFEx
2L3wT/7obIn/sc0Y3IodcKhKibRXxV0xG6Q4K6mwXW7TnN86jrusFdWXw2yRhvBL4OLGAu+xC3Se
3wjs7p9vNmP0rdCIGysJ0hQMJhjA9CYQETzI1XnxBkC2R6aEBDxSCiBFElKA0lHFEvvlQtWX4+au
Vmbc8w0A27HhQez/swgyPc/WttYBXcQkaMp1bSjnQEAnBhl92cxzVqjzhcE1NJoxymYl2dKDR4ih
uQbdmT8HOyj9xEJCxTqHBabacEHymfai5RRRMnI8NarxS0j16YL4up2H3ELQb5cEBtr4lRgfFRX5
jf42Cy1jDNSHjp+4Sbjf4kmExMXQAZRGHGIUhCxhj4w7MXe3uab8ODM1os22o3F46jVkIlFDZ/Fe
VM96WOVJUrIKq0BiNZXCXbv/Q4cNukA2n6Wwz5N1deNiLTA9HbUmc2w30y0tNLV0V0abYc7D7gC5
9D+/LoziGQpje5MEL+D2/2fXOSfCbRaFBPCQHD9UuyhQ2JNpm5NP0VWwnGCSL4p1HLTfbQYRLrvA
YlxvkWiU4gPjWfjXQwhkeHqLlpoFNauwjtWafxPpYkgpogEowNZ1els4EutPyRo8OWSgKAE7ZFkM
kPhWOu3Ri8tRG2yBX4xU6jI44sCANaT2otR4uMadSBbzYtjbxZdjLm6eJMxYOpQcjc61EKD/v2Y9
FGkJsWVvn4ZdRWkU7N1Ox6/cMb5SNmO3RwJQHayuyWrdPfCc5a7axFvlVxGiV/yT2FcPPlGXdPE1
3zPj9kCkTGzvktT2hvAXBQAq63AIJHeil4KQqiZnCYDLT9XxxTui0ySYo3d1paISwn2xKkqZahQM
uWbHWNRcqkgyjg8sNMJKTpICVaimgtk3V9XkNs7f3rzQLIRU7XKVC9rjNokzYcxBsU7xjUgnYUZV
Ig5V2Kx24iFdKPwDXtG2EyYjBnBt+Gg/FM7/4HM0/r2zzsT3IRWsmL1rBS1OXzDDipC6pRT/KS3+
kjbjBYugL+xU8Mpqh5oFJUm3vNSJse08hss+ntUgtp3Yhb9gzToYrSNc2bqb2O6omrSNC61FtBUN
Z7aL4CfKOXMVCjPd/z1sC5NpMh4c3WfWIYoYNHo7/ssqaETCg0/ve7UPPehG+9Gm1DTzRxEgX70E
/sCyK6KpSDZXA1pW8OLjrNvi3IAQfaJyIgk+DrtZLeBa6q4fQOWNZfe/bTwcFDFbJ6BFoO7B3ZHJ
2YNGcpqbkYn7V/gf7du1R+mbk7hQLJbHVoDoOf7dGo5GB9qh6iiEor910nngaNF3Bbv4gTHq4O+B
KY76xmqzQoUByYqLvt3yXm/eOZHaPEO5bR2fURmX0vBAwEpybCpqa2zIFzSmp+quL4qAHtR3ErzU
z9KdgO+lh3qXVt+d50kR0wcTWu6pXVPjKvFd1yFkyl+dEoP64X+56HTwtdE0G+eTs90wSw5pOsej
ey2uqkyuhSX87C1jjcFNyktlkSqpTEag2b/2jWfg89e3URGnvO58szYvgKB5GYmX0HOBIZP41wP/
8s/ESk//azK/CkUlBbxodnB/3x+l6wmbzTrfXQrFbAiQmHNJIAGe7cmW3DvdZAc9rR4sYoCornbf
QEffocNQY3SL+DTxc9Mc3Q6Bes/DlF+9/y0dM8L3cOv2e/BOWSrnA9GuJYixJ3QybOWYo4neGSNF
bxpiy1AdpoY+sIWq73qKUqc5sBrfHbwvx7dWvqWZ78DjSrWUjlxspvaxKltxtj66OiidIu2019yv
xYs++hFgiTUypgOqbaSrxdxomWqtD5diD1ueudldvqGuJM8DnXepP/OPNfjXTuW9M9whaxFsVGss
JUmXj5yplxtaxK68mKoNgKxKfDIxDDZIBGYl5JKOWRrlT1oeeRkijXaFaNRCYjViTIhYI9fP2UW8
xdO3/j7Aax45cTOhJoH2KnyQOoD2oyVDDFrO5ZDpMinJcsdEucUjFbkUWWRk7GhCSRN5ZivL6M7/
LBLRN5D4LHs9bTXsj9q/6k8rm/rdd+/LDBLjSZxaBTykgxAMgf9ZGXvX5RH/Z6+4TKJpNROJAcY3
sp/a8i49onNHiex5KehAmlZ2NSi74jKLQESs4RKI6rjXttGiTzdPOyAt91X4C6ny7PHYyaQyFN9h
sOvLH621delxfxY0/7uXsw+5K+Di+KljZTmRPrM8VtPh682Sfh/ubG+uyiuvjSS/RJIcQdY6QitO
3zcK+/bg3fwWqDkor6wJlxxX8dkMnjZHaIANoTFfxqkgNzY+obtEbTrwzTrVV+V7Qe+hUT/M7GTX
ljADSC0/BgU3lMaW4dmAn3fdk87wFGh2zACnj1P5k1oV/pWF0hWcrZq+enPx9TDWqeIhfKLc8NzX
doWGSp/V4pNx4S5W4OejspTvFGQ51EEZeo4c0xujpe+6CoaXOJ2Rl+/CvqlIDvJILVvYUbpon69j
qfAqVJ0nQe/4v8WoJcjNF1ms5jO6OLzO5Y/HHDShxoXm693HIUpebOZqn5tzIfwjj7/Tk9KXQ4kj
aatG/M7yFj3D598NbzLTt/Mb8V9IR1CJvmiOHwk+3TXx+MTn0QOkStMN7RMe4VBNCPdSmiOFh+vF
FWKL+hYcGrlMxVd7kn+cDaawUIo6AeCsz/3B4lOMQvL5KAyMDbG/4OHOqP6Jh49Dn0NUokoUOKZA
d+HigytFwAVBwFZFZHNlc8lEZRFth6m2SHgViFg9C1CZHV/CFb8cQkemEb8nr0baHuJhXYo19o5U
asL/qqggp2+OLIibWehrRpZ816P7xgKzIeROsTRLgPXFIvsEfISKx0tNMzRodAnfdcGrvM8coA2q
npB8+yAp6Wbm5FmVtUKTcMFeiw/8oshmvRt45qjxPw7IRQZYghZJ2Kt47wHteIJp+rdPyhkp5Al2
xMrxVsaKRuqSGZQiMmvcQl2GlzQ0LTapDMs6+ydpjrzieMw071JzA3PktaeyqME5Rg57/4WpEHxe
RWMYeNCoAOxRPxY2iVcODtauEdURhqKCFsDJCl3vE8+x2rQQ6JHp87gUJhAo2X1OmaLjdUNUNMpD
VFYy32r4LhkuPIUSW1OC553/DrXoboMQf3PrmZqZVy0/ZUUBFNCcFVQn0jgtWyaZDR4JnlfF+biK
QGxeLPqz6zGxvEXIhny36jrwu/IXCBDl1nIZtF39x5JYPt0rnHMuBPvev3B+yLCLGrrrBWghwjf4
kygh7fTf5RlOlCZhzaYMAYvXdSNYViTDueOeeMWGLYfXR2u9K+J4DpKUkcRqnCgImcxbbbklu+MQ
ROr/XrMHo/8y8omGhOZjY7oKJQLjpEDCF7H7dwDi0RnqRuaI1lvkqBG01d0WjRkjp/aonHyzlRfM
7rQprDxu1RDMNHnTZWTatJr3z1yyP0CFLsHms/Jv1EWFvY6XURF6sDxpgLvhKG22T/X+3x122yLr
WKIvg8aVNr3eog4h8vzOmStgheKDGDlXdPG53bdeFpk/3OaaGPTfd2z0cOtSleQ9qNk0qIU0A92c
bqm22YKfGQh1az0KpKxP8OmOoDBhCQbvKuCrp/2WHVstk9bFkwPUu0maJgpkCBtqPiwhVi5Vi12I
Hd+P+DzJPj9XX1lXnVoQiiPUEscf+NEMJ77p6lSMg8Hp4G+2vaikwuZ/8orpFKQ7mFACaZB4CgXD
/QAteCnNcTQPW0coq8oZ6l7xs3He3Awt7qqe2XhjqeglYovpZ3j7eCgGegz4favmuJlcKxwSixGu
zzo2SZb08getSZ9TJ7//ezMvLhMrh3p+1YEBn+EVz6i2t+SjocFhndxJ+NgqHP3WooX21aPHrU/C
XKi4Z/3jDbGze5ITZ86gGHbx2bSetuUnH7UnJkZxvzedEsq+NdbWhiES2D9tkJ03d+grs1JNM+Wq
asJexs7oz2kSHCfyk8XztKDOTB2R1Sdanqba+m0aQK3KColvdblZWlSRuOIooiV/4qmEZEEEat4g
gKRBPvqJL2cgWO/JTRb5P0ld67mb2TyH7zJO9qMXGmVKaVS8cu5PfKnY25BChE8J9DpxFMUNZbTn
2qsjpHN1GFXDilBTIvDkVqr40kes27pRAvWhpXDe6BVPMX80mdPVTS19Yzx8Dex5T0s+umZjQp80
yB479wY6l6zqHSrS9/bGKUnwCbvHhsnWpZNyS1bUqhc3jdQd5GjGNlovqw9iWOA4NpC6oOKuAR0S
D/3iKseJLUTxQ20EKXPACD0OC4mQZXVxKlkn3ASSAKqHe/vR2m+IdMdoXsHZKQ/QSvWrmrOhcUVB
Z9tapNYYvZdwpJAe+Vpmb+AlowlhIWFJQO9c9uuhfR/+pmWJUKsbLnXgjDWyFeJQym307fB9PryX
NwxsWSNNhknLwry4vaMMLKFy0UCW59fU35ZCGWhai/1Z6kPOEg/FnohoYh24n/+7O9YOo7Z4Ppdp
oE2nBC/GmN62Lk/HZxfI+q92JFi5vjZg9viVkCcW39+yDXmJMPUWYiB4CiMWPvcqlWY37HeZpc0l
PEg2kyAXvPlA7sA5ca0YHgMGYPQe3Lssy9USb66CgtcBX7T9ynlk83auDte6A9uO1Ys7zqAYf9PV
UBLNWY6dMJw9rmjOt68MGA2ZnAoOTvBw0ZJve6PAx7cETlyRFW4Yue6x4eIj8USqdE2cf7TyTV6V
Ox1l/g3TglXgjr7YQNqkmSYl1FlWgKN5Ugi+2yutv4IWgcWGWeDFdhsjtWIkPFCimsHCl4gKQFWw
nb7kLDf4etoQ1lejvzwKSWcKDVMtv8cVdUcwuORbxgp6fvUcwB7qQ/0Yqj5KDyd12l4SiTJZu3kA
cTZl0ln4LLDXwmoa19MBBoMBG1vIufN/tX9ImiOBpbSuA097EWB6bO0qhuI3jdHsLTqidpXvluLn
acCpWuZtQ6NgVDLyVqh597jzye8AUkk9kgfMN0SEkm7VVdzgnOjGQ1BE/K4zW+UPgW8A7FhdHNxo
1jbvFSjrCdjPCPSTxNzfsSIH9GCzxEfPtPxNucO/XbEb6DAagnqgARO6wjlohPfU/nvAaKTrfoQp
yPuAwb2d1weEp0RjIo0HkNCCkB+J2ffzca2eB7ph4KIkZDQUSw0RAqD79rNCbJqnj7KPjCRUf1GC
XZhpHApFxgr5jTyPBEiZ5gIp4581Hc9BD1bZLXUhYYwBMpfkkSkncXfqssa5ka2um5bBXHFSarW3
2N6Hhln048z6Ord3s63RlZ5Blx+cjuSKTZB+PaRIBspgj3ANpSNTf8LzdS/ClwSOPscw4NgVI0He
8vPYq5AOQabK98xzCqZTfKi7hYxh0PBTuVbxkYsEOLefSAAk0IZfx1sLpCpJcqSAQJnOE6v3MEZY
0nBc7ckvZoF/xKn3/EgPcuXQG0q9wk8fG/6kUKMeWv9rkFjK7ycRGUaUORCVrO72o+NszQd8LChN
DUzMOpuA+MmY9/bxKapsWgt5ufr3gsy6qUCeuCThREyoAvbqylT36/l9iZyZ09YY7ihlQ1XGFEkj
4/cKRiXSO8s8HobIwwqFDw/uMvfE9s9dbAcNycu+2BKPg23WDBhohHoTAUg2yNPUOX104EokVogf
0svGMnTYt9KZnSr0gqfEYdZetQQev7XQvdR9E15xlRZG0ZJZgAcJXtPTjl4+Uooam2747vUKCiXx
Yy01BcCJ5GJ11oLSxrQsCGQcN956d1O3ZXBN7Wt7oSoNZ3FZtqAYOBpU8UBV7RH9JmyeBT4EEzgU
Ckkp6hg30d/BN3PPLi62jbtBKWmYzstUbMdLX1laXDUiquPsJubrIo6PjYcVDGZ81JaRrHcBlHcN
+vAnmcIhdlPvtLGJZKFEvh6KqjUku8m6vNJ7u1G3Usg5PC2ivCHAnL1X/ISMjSUZTuT6rwX3ODS9
vzDhERzih+8L8HPNA1oVG/khVf8PVZAMiywUlu195D3T4VK0NTLySkgPpddRDtYkp41v2aussCec
9xXyMezagq0dWphCKeu9i7eqsqm9Ibft3r28+2rIAgYNiImmzB2956i2v3dOpBCm7gjcoST682r+
LGKejsHANJW+ruAs4iUMkMhh7uPFu2RU40+bRKjz7wR5WWvAdJeFpNegM21mRLipIBnxZaFhmy1e
gMTvdOFLWS30Qb80jOLXurjPakBXDZ/mmX7bZjhcO+XMQdNG2X+j4NwbgtF8vdPTeSemeUN2JIHc
AiQ3iSDGDZJ0UWjsb/tpoZWnOFpdgA0N8btB+rpUorrfDbJxu8Z4c66oqWw2dU12F63PMXB9J2vi
i716vZYTauDNE2KkK3iRmOKbELzSRd+rISJ68B04TynVyk/Xqkmqz2mpxczJb2th9ICwOiPrWJj6
AtL1xgNXnMbgogW/GkN6JVgh2mESYQfJPvMOcCelgSYzOP69440A+L04Bb7GEgDlcm15B1Etnqba
3GN3q3iuVPLMU056S/+wm7ywNOfpAllCn7G3ab3YjcHYVYqRMtOZ+3mLnibLMQlg1VnnfmWLrNiw
LDSLioevZ77ck2O96oAiZENo0IhfV+3MVN/6ZTfRGhQIak+Z7Ki3L0mdmiwrgTNOLpp2YwtaY8Ql
V9o2oQx8rRTZkLVcTLRiHF6wUkM3GAdIXgCZfsL0TdWxQvhKTvVmrZqIY5ywhWDi9IAUvVgARQWM
4s4kN0PCsj2VATrRazZ9wDwN9VLHSHjnW24WNza8HEwstJUacz5JEUBlGKTLWsmg775HaD3gGtzU
FnRP0sXU8Ul3KaHrfkd6Eza2HoM2Z24ChLYzcMJO8Leyo9WAmjhUai3kxdEm5nSOd1ehJKFXrYpq
2OFN7OtibsHZJTkJVEJM2B34xWK4e2cYt0FrFjOlQdScKe2sr3aevJNVxxB65AQrPnWQecbFUKZV
BfPEQ3Bxpn7BjlveecQGlvA62n8ty4279XJOikwEx+O8hIii81Knvf07jSy55S3qToAO+Hs3lkdm
HdfCQ5nuL5y25C72MhXaSFMuNgH7CqOF7B6NIHyGO1/BCboZjaaWJb8pTL38RdjSePw6na9DVB+6
KMOArv/ZJly85G/I0Z2FsGxIPIZvSHFuQBRck9K0tRy65wb3w5Gd0Kyggvr9MiAY3XUG4gbdpaeF
hNnoqsh/rZJh0hb3xzwDW2pmXLRHA6dn73GbAQ8cptHcS3Ikb8+FvMEMftm2Kzcj810/c4E///6Y
f1XvN9FQM3lfjSHn56qbb6F6bhwL9db96wY+peY/msc3zovqn86OqinPoOBi7Wso23iSvmadSUBW
JjPo3/vzbDKMkxmMMZCxtJyxfvMA52ILfEt0giBYe0VQFlZ44DlCFqZSPaVko/niKoCkR1Z13s4L
uvLnOQujLh4NrXLesiyn1l5APXK7M4tyIvhPwRe8/D9EwK1qu649kRP0w+VUBgG8SyUu53w6GS2S
1F0dZjBfhivZULEopW3McLXkAJ0X/JRYB94ON+XyKmt4cnW1bW/VoG7OQYTiori89hgOlsLScBND
OEsqq0izgV04XIHkyyjbSY64pMNXIk6RxanjXNu1ObWNY9J1SGrssozMbfCscWiJIn8aIIBIxl8e
yhwEfIBmmjqQIoBb90Y3JQ17yVEPEFOKx9sMqb3URrepY/wgwqxO2+L+i1G3w4Uzm++SENcBWfz7
R5NUxNxOfGsFD6wHKsFq5zEgl6zt4fhRhokdwb0e8mTvIh9TTa3GOPKY9oOi6ox1x+1Rj2dyLayA
vrroLM5vsppStxpL/bE5TZTMwXwpJjA69+OejDO3xZa6N38UR1FPfdNvuI3QcGtq5Odj/8hQGQ1x
PAaCMAE12vV36nnLoy0xT9Rdy+Ffub2ihMQ7UZmL1MqkWbolz4oJiSmT6BXZ6KbD47k10SkbfNeE
M0lny3fbNnZCpD04OtFb6Be8JB1+ff76EsQOMI7Zf5wcHWSepZnoYyS8yLi3vR0jPdD2m5zCEPWy
sAi4XPgCoJy3oMELvbAxlhxRnUfFPxqWhD7xxx7DYZM707btr0uOBg53B/10VYgP0KXftx9gCyr0
K5WXCwf1lubPdzFZ9svcfgeSBOj6g4x1lTR/D9P15zgI9BZIyvlrFWxwb9g46ww71BxhC8Or0yO2
j5ecnDqmT77hUj5rvSpv90gZVjD42aZxODxWUzNoFqPwZOeeTxq8dUyDQD16bt/n0YT9wHxHvIBz
lxFOtNFlwTWzPjkMuG26SmfWPW8MraybHg9+YkOzvj09svGi4TUyy39ZGCD9w/Hc6xhNS/PSO+2x
K6ndqFUbUeHJHFupssR3RlY5wo3wPQrhdUm1dtLAeKboNLOJwDNbLuTYBWkw+EuDM6erNMjI87z+
HfQp2KwH+AnA31euwEyPvhe/FqTRevB/Y2RMPtEi1wEu7++3FlMoVYKqI2691HCmi9Xd9FGVjXlX
E6Q7RWLsFrpLwOrWo0hDoydCyXy8ilCggWgAhVGJkVHFAusDM4JkjcKacvXi9Bbf+H8TmFZrXYb2
tVQr0szcqnKQmyqfX+INoQq0ecuG1skapvT1nFWqZkjHwtS9/nnnRrfKZgDdmd99XcC093X63V8R
9ZS96yyr1GAVrJ7CmtBooJTMA0MYiSduF+5vbJN2Zofz2lHIfaaLY8ezWyKtyzYHPQs4z1aJhYFE
Qzh4INASflPQ0PNHQu/hszDuKfnzmdCopGlSGq2TblIjXmXPH8mL9HXkT91puXn71OKNU3Bbo2hn
yVphN49Cexfv0j5+TqQ8yN4Dlh3uyuhtx76UkS7LsTNW547biYBCusfE7zHGUYnhEjCHTG+h+wj0
pyQa8bB9UFUOmiyEnVqDbVKyKT115uItEGQWpkqTYWRNEP4ejrPyEwfxXh9bwwCdOl/r5UIEN1/S
WDQt5qMF6GpeOKfI79VZfLRVJSuc5GF8OHYO/qFTiDjA4kZNI40jwbzYQUUC8TzwnEuEFaMck5dj
ergGRyNhlmu2DnMRmlLbLoKFrEf+Pbd7GXfhUY59gTebfNpu0qw1AvM8hUog/iFXFQAOyy4/gGSa
onH4Mfpp6aDDDYIdfJwLRglJNzQKrSacgSSHvEYVjWh6XmwIxvFgFb96gced/bgxMHfJeAddelrn
fkTwumbwnAPkcvUJp+XI0UOybi94/Bwv5o993skmUFRstKUaGJh8pOrpWaJeEqwmEqvmLpUSSW1M
ut9G/FbesxMGcBMBu8zcI0qP0qxZ1UKJBMZ9yaSoKqe2xV89tAnhl8Q2whzwI+Kifjc6nD9jLO1F
praaPyEkQXxo00zXtiRfzpk+Au7NCO2Y6WVnVJQaIryq1X5DgGwisGIPASFxRKskxqVxtMe6KCQp
nkyqM6f6EB3/N+88LJ45Wg8eWPuP7k+M2maFbbh5bK7iBT5kXZC/PxdDwLEKgqyMyC4cbBqxCJSz
EEMTot1123OBCa3fsgvzzzA6uIY5DFAdvLcPw4Y1CtBloSO3PnU0NocG8nVnz4aRU/DMyPUGJHAi
4Ww9wLFkxhgiS5q1DZx+JREbU6EcG9nYdnuZuyY/paxXZrYP7466ZOAaeD6+oGXkNgp0GKXqJM5Q
+7fXWld1OsuN9CQEwmp3Kp6tBsBRKD5RiG4bDwu/KdS5p2XUorpMO6vDN9ix2316WrUY6oSBVYgy
iamAXvRPKRNKWt+8ClxJUtpU4QjC9MmFQU0Nc0sVahxt8gITs1Bg0dS3AJ9jDnCcO+zbXi7FN8oP
Xlqu+NjV7gkud9XJ1vs2Pu1I63VoX2SoVXwFrzTuPsJxdE6ADywvF2N3laTA//sZMqmjPe2OjiMH
QP99/m+fmwtUfVee0Z+lC5FpKY9n8oX+fm3vGdsaR+OFgbmgLLxjJQXhICYpzd+3XoYkQetwALeL
2K7tZxN+SHpAkGx33O8vewcmCUU+cjMz/GVLi9aPLCldmux9Xtzxo3Ery6fKQUe5AIoiAcXArxoA
sQqdemUP+gftNRxEKoOoAZw0/GlepgxUhl7emBqoosTLXLghQs2F7tcgc4waKH9McoFaboPqfWoz
1tvzyJdP06hAlhPb5fdS4ZRb2KS4P+U0tRvQGuX3DDtt+IFBIeZ9p5HKD/i4nup1r0F8iBLfz3Y7
7JWo/AxEtSzPnnOdNybZeIgGlWk12QMUW/zdXQUu9BcKCJVjtnA0IVUOMvQmURKZGjtamOquKzR0
SwsffazHdKA+mzgAwrZPAjZDWhINzpC/Ox7JLq3VivBAxzDsDzGoW9h4zcrLG7dGzYLcYT3U9cay
B6XVZc+BUCzUlMhoahcMbtZNF9+lkldbjiWntRHvujL3/EjgBXRli+nwoKHeTcwShLr+iwGRS9AX
nXdPjztipYaeyv0tM0CNJPUGaCINe90HPxFG52fdKo6hYoCL2rvmEe7cArEdURVV8b7if+I/qwVN
bB6m6bV13Pq8gY0aI2xv6WQog6624KAeTmKfKI+C0GdaQXCOU3EfkQ6ry2ygvsUILbkqFxtbkT6o
Z4iaknM1zJztk5alJKCjy+2mcA00Jow/laO8kigI4sqK1PGPhdQPUkpV2L2Hsr7tc5cFHqLY85G2
Tz3toz5D5JRMjGY1FcOuDCF/wXqkWXI8QBAlQNljDPwHT5FLGohWZmNMPdA4POkUalwZKHjwJq2K
UGLvxzuShCAN60JKv7+RpAKKq2W1xts0/ZP/LBhasoFdCIO/1rJ2YGyIK6mOR2M6PVBtglvgy1hB
CrkPkMfs4bm9rAIe62zdg+nwaZhLuG/uCddNAUSMTyqdUv5LxnHNzwEW/XtWu3NEgKB18OpOLBkh
yScGhOFoxmezG4ou/zylhsy9cZLO0SQqpPVwSYBYF4k88DpUxpGSg4u+TIpNY+RgjN63K01YBoQV
6AJB1lF9RPshcrtoIAEnnWDg+iCVsPBCBZBi2PgoOHCRv2rXjM9V4SB5ER2IrGfHj+Yj7jTNnRD0
/gATHiLOSs9x/3wCUyw0XfaFlB7lj2Zm+kzw67yq6klsmv94o8ukCwC6GfIIVG5M3+x8joPHt23S
o8/5Zy6XJ+ZPOPX6IiMvU2UDCs2MvKVsJVkbip+QuTDHMiqB1AOFQQGdTT039gBaRzjcEUaxUz7a
lWqNkc89MgAAm1Rls30WRDLkeLQH/aVt0n241tHAgsN7yP30meUITp/Dr4fQD1gFjoMb5xPFkYrO
TXqmIeWwELyhQxIUukkwv5z/G4b2mUbjKqqsP8PJojOlKHmXzNk8RA08b+Y3j99T0Fmq92nfa/Qn
BHbAW0RS0AuBa5Wdi5tnF3Rzn+H2N/tvQIOS6vRNynkfFO1N/Oy9m1jHAGL5guX8oEWDbK2bv0Vy
+V0c5pRQ+5Egy6zkCKaXNu0/qjcwl355aduZ5n2BBdOhPeOnDrpT5YiL64Mko9wRNo9EY52+8JFQ
/w0clPbVytb4QEyl2hFdlK9NOa0arrgVRhls6Y6uskI+35cOVQYfnV86SKg62MjdH8iXBcZSJPss
cTAxJlfVJuzoeduVclu8D4cFaTIwEKqD7GajGAr8CVFSuniJ9cBgOhoRqlXZVoP7VU9unrHj+E4u
Iost5sKHXvu/5ZTw8IrxQ98iQ5rzg4asPvBF8REG/PLNswau9Szwxn+yJa0EZCB1Oqyl5fE0dGFL
MyXIAwo8C3Dne6WMifjRr4ROjY01MRBIsFH5WFO3K7eUvWg8/1BumKH2XWG3ck5lRVQ08AmU2byv
PuLy0dm28vpkoHt1u7lwn8kahDveJUcssTfXxxhWeaS7b5Z8CtDnoTvaHWtXMeimUku1146Pn50n
OPXEcHsnBybhKu/MXogZIRo4QMeQD01strZPhpKoNAibJFneMy0Hh+GL2EIf8glv1qrp0CyJmlB2
AVGBIBNCac3eaAVTmXMBbFe1giwSpG0wP1lR5VUisifYfwBLc/qT4ulN2W+JRQ6yAPLFBWYwk8ub
2yF/CgWDdgzJNh00D2R1yTGHZbK0CATpC2r6a3dztt9tU+O7DOsrskdh23axCAuz1OK8DQod/rTb
CclbMWOmKVYYMJ/FdAxd4l2CE0HUbxWDziNgsCJmUN9/r7iFTVEZ7z6V7cpdPx8ydNZw3E5jG58w
4nzWvvMapmTL2tpCafwGFuAojRdADXqYn0nDqdxDQEGUMiobArD6PbP1fbpBDDc/N9DSXQyKZF3B
OorbjxTM/6xVT/EsK5Qh3k04+cZ+yusHy0bN+F6dh2hewA32PQJCd40dUYtbr1RKs6TtH4e5Zago
k3ZfAlcV4OqZbP3+t2NojbFYQpbm/pDIQNEi9AZh4RHSuWb5VXYYtvkqB/4+rgZv+IVap10Sc6d0
d9sCiUq815iKzOCDOmR7ytzgD8QAM5xj9YtEomobGsBArd6AdXU/3mN1YIZUJlMQDTG4GOIRZZza
xiZs9BVj+s5D4l4tc9hBBFyuRrZ6VLS9sKR3bHrGze6MzbBT6akLnfbVS1RBtXLSXppIWyrYSGYn
R2jNGJdk275uhQR3sbu+iCgxfMiEFRlLXrRCfiqoGK6Ce+8ORhEDhjp0TlD0D1vfJcmtXCm68vyH
rb/js0pKtpfSf8XQrjOxsE/MLmiwyrfgniXQFyoNDDkA1UFUdmeP9nKiLcjE4O81BSi5k0HF1bhc
ngZr7STmdgSrtp4z6QtZonIEgQf9FzXJpPMJgtV3hti4BPj7JkU1F0qlAYMXArpIkJ3mFM2beRnv
Teyxsqo405qzC7FA1U1BLT3kT6f/mxWz5iW7emfHzkCxZhOkp/gFH/5N6IgN/I+XemMLH1zfC2WH
y1R3I8DjiptfYWcM6gTOKlTjkzOus9i4bZ9XAUyHduyS4Z/Tvh1vw/UPm5PIwB0B7fbR/msTI/y1
Or6x6d0Bv+ilIpbf2bMq2oJw7/xbptvDjrks0f+TFmYpcxQzxpBiwPiykD1rRJX77nfDQdkQLfi2
dPXnH2MxpoW8smjBP/sa23m1ZZVCAM+qxAZx2oS1GuGWhjMTmF4fd8PqkBFVDDszHm1IDUv7AF+u
rETbG69ac/GjJJS5k5UkMtwCUGWbUsuvvKq/8yDYlfOWprDysqBf4CnOt2XJva2O9nwJFaVservK
K+f1C/V+AeTYsdt4MqrtPbF/EZECfaIbyBg7GKnmL4khLRvDlnw9qVP4ptUbZz+AavinsZarDB/Q
QtRkM6bNXyMR+eAJMq1IJ8xGSQU0SFVk1Av3LBKRaRtGzw+IyByJnFM6iBlQJ7yGCZBQ0Pj/F40f
Z9gk6lbfGP/s1FKG5ZPO2RPv6mXdSWnf5vaWoU5uH4WDZQsVUNvAzKrEUtehNjikJPI3ZxjI7AC2
3iPARbdXWsziaRu890FABzcyX6brVcGnAICBjZyv1UAs5JSYONVjBEy8JMxWkyyHGt3MMEuZOjrF
aAUJv9BfFufY/ksn9cmIEZcPJj+tA7iT+6k/W8k6vt3nle4ZNA7K5g6oxY1WGWkKpcJx3Smz8Uio
g2wsGYNXHo4sksffJ/MxJBV9lEspPUZjXj1zJtDmEYzCMMago4cn/I3eOtkTxv3Zk3srrnmRXgH7
0gT8iHZ6dbkLuxA6nN5GgiBPPdXnfejrdGhAeku48eTX/uG1QTbP9Hx4rij2vsMtwheL7mk9q3Al
cLUNaSDcyJIDaNfoD0eIu9+rZgmLh8WptXgYQ7Bs9Eeo2GmaqWnBTqZh+C78yvPFYolK1/4Oe5nL
Sj1qu5Y/6KBxQjeTD5qwPRnHNM1gIQctoQ63G2I/FV9xZijimqen533OFlOkKrN3PqFgY7qzGmDD
JCe5a4woSuUEOA2g9snODAmAfRvUPsKpn3A1YpyOdxO6m3YkUhhrExeIiyInu42S8mX0luG5TCtt
5L0SilYbEMYRHOwgF4shhQ0PSmAOpN+3P4e8mzWDo2W7IcqNHvjC3p6dXcc9xfP7daMShGnoVODC
2Ba63nCjmZGcxtgNCiJiNR87iSInI6gwDJdSo32O5nSstsU+IJUDuehxuI6C9hfTV9JmS3cYUqPF
jW+zafgS5NPvWWAYZjELortAl6NbXIEfKtvx8bMY4WMzk90QurCjKXs6yJCNNa7yEaNq05HYPtv0
rm4cuF4eYYmePh/+D7todx7cSLlkXTQnN0upF8/oFXoX9L/04k5hfvzGhBSIP0useAlpYGfR+t2Y
iLt+fo8ZYsThOWlWKy8af4LCEHKJcz5OdfCw3vODonmvlzo/G5I6OMNgX8Lmc2iUsO0Ca+5CsIVo
z0rJCgps8LEIMnfgSMeNFByA4hSumLf43Rl33i9WIeHVpISEY1ongG8LCfwCEBbU7qOfIfg7AKgg
UyR/1aeqoq9gdfzMDjer/77GCaGzhFrhhNcaU460BA5Uv75Q66EzcS8DmFUoCRF8PwjsE+pbsXxp
mpcJTTVM9iwV4ZikvYGTRL6KdoV5Jpx93r8jWdppbPpN2utvwhUJ2do5ICNz+qgkI/P8kSX4JaN6
EI6WDA/4J5dJONI0DEhFXGbttryL4eILT7fMu7/D4a4q+nDjToM4ogN6b28LQD1fAk1IO0BHWgCO
XHrGWzSFph2sGxB8xgT6YAifN7FqLifb5Q3t6NftE1e9+ez9yuc0Q1MgjffZMi8jRXP+CO2eYaKk
DW3UnkmJ12kBzw5PAqpKOY8fmgq68uOHn26WlmVF4FKNjCnq8eafwN2J8hMrH/QFewXB3Q4CUl6H
mHtEZjcKeXud3FAH6eaqMEk+HuiJ9agrluIQnoYdjLtlt+pScaATnbmOCI21uf1Cevx7oaObuQ6B
QRDDah8V1FuyNgq2sE3lOYPIuOgAf7cBFnaG1Q9s7/6/otrLxNSaQmy/UeTgkcE2zNmFIfAIGlY7
MRRDt81wrwg1U7Q/N0+bonOPzJDC8QaPSWRtwaw9abm4b2212AlO+EIqwX2M/TJ5lz/P+9ICeUNG
pH5bjh8GGYzJklKQwmQDUh9FBNdxr036/vHBcVO3e2HTEOotclUt3hzIIoaUCCPSSOrVyNGET2qs
+PiaHLUh7u+gYqN9dJ2W6O7gJXSeB3J9xQgtd7C99TXHLl7YyEk+lnu8EMJNYnqm6VLQ5IBwIzb/
ZFBtSuSNGzzzO9MX6ROoZWTQvcHWP3ATqYg3sMLE9ZJGAYKf5cLTW/8yAq9VpFceTOtEXPptsClN
IiQJhn+JxUxuiyHR5ZhQ2dLC7jsbVoRBSa33IjeAqK8DP2zdhOEH1OLPATlLYPhgnmtjl3ob/Uq4
ful7fN+oFcBHpNjpBXP6+waffrKkfaw01xHTMgAUK7FJtxX7DBXXHQcz5vuMRkn4EaX2B6kxmniu
ceqqhfn5Gncym44ED2E7zE4FvqDLtEpXUJD615KD7hzR3AqlX76OV+OzT6uBQgIpdzkodqlH8ZwJ
m/uL1ud3KBahfyTcweQ4vMhQvXHBObjw1kDP5ogoW1ypPMR3XDldxc2sfo8TkyI9Yri6LouWGHbz
clzn/HGyjVvVGHhYT+ksTkTTDlvqOCJgpzUQxzLedlvxh2okWhHUWfkBrwG1tIdEA9dcXyuZvglT
DRc112RF80CUypy53h9lqwGvbTEiHfJne8Q5ZT7l8s2HXT5JaCQRR/cd869pUtuDyaLRfDZ8iY0v
9U+Fr1DvvdkLQxz5W5Mtyot6VfnAnQZWn00xZpiIKmPTcqg8iOdZ3/x6kaepQy3yvVb6X238VZ+b
Ku+5yqmsskssHdnjf2+q3gNwdxXG7/rubJg3sdMzJMjCAbfmT8uEdrjsflrsBm+tlcfrgTu1+d3L
+AJpgOK/B8vRMFpOUxZRwuNbsWizyZf0vYhnib6RNSW81a3pYd24RnfD1rBVGQXzkEk5HFSMdK/g
XvqO8LWuW3YBhPk5qQBbqf8tv6Kbilf/remUAZZxwcQ0JJSLoKsng4TMx1zZk9RQPgODj1zTzTwa
Qu8wgAsTibKZPdPjGawhVj0pVJ7DEDhJZjYUgtVL9sJLn7MYzUrFOs9g1WFfgM2jniqj5+iizJIC
iC1BG/ALaxGSY3+ssv2T9oFCkK1mbuz1S1v5LgR8r+d0YWB2cpe5NJwDuu4FNBNeiJZ60fYVp8XT
MpRpixF5DKKHxEJL/If66V4ini5WRBUGftTG545ygtwMfdUK1GegCbv6Yp/60ZPWDjRi8JrcCjSj
2jQWUdLyLbXjrhBBwSuNVbDJa/ONbPAlfmaHFf9+NX/MPg0IXeXKdOhjWY4L4rrFjmffCX9lXgcj
reA5LEwqKoraCFxbQ10YJN0b489YEd6XZ2Iy66nZF3hMWruYl4fW/BvZtUf7p99qCzg04G9dp+pQ
BT6Thn/FlqJooeXrAhz6ULPt8jCVwjGbN7r5ym5IXbXOZymOVpXmVthFK6xdF6FC7bUiEu12u6Z5
ZSTQC/3bq6M2e889C0eN9GMNQHlRO1gHQngbeo3nzNNIIfD5nkSerILsKo5MSI+dDFizLhEr+1WC
lhadUSGmz5dmnlxP7hUJuYGoDxPoCo9grBtzK5a0c8Eex7oZQxTLer0aZklgSK6923fs0EyefFvV
aZ78IbI2qtrVQcfcZhP0/flA7HVctAERKEnBEJLgLKFneEOf9/CvWrA3DYtE1JAL0CGIdfyKr9Oo
wdNVAS9oHh5ZhxIVQBH49RI0g7DU2L8Dei7sPshfuPifjj0Mub26swz5q7ZkkD4lxD87onT8giNq
UfLpDygsgzzxRzZx34uceC/UGRKRZzIXQt6w4oB5Or9D1iwo27L5tzhGVbu+UCITOhxKoo0WWBLP
a3PhqKTw8UapoP6hpPrzsS0qDBrC64AIWCxL60tmLRmfi0lJ1MUVgFt0rLqy2q+zZosdNyWhdgTy
sXyuYtX0TcJy62YarpM0lsnK4vbp1mSXY0xWkrY/L2ZLJ4t37QjGyg+b8mf8YjQzRdJgZaayKsSC
HnWnHsZ67wAynM+qecLA8s/8nkXDMAAo962m9Z5G51h3lSzMyxB0llMBDzGLMGb7YKO6+oiB1wTL
cS+gzfcr9wts8F+fToZPYBJtw//EkeZdv1CU+Wo2n8UEUXDhezvbYytwkNKaya0Qo/mxz/h/8HQj
ICkTR1Jtz34NWPp9Ny+H+zPR7mJGkoEtcjufpLLc78mrbnm3/gKGA35z11GKwcOr/Za9f7wU6yyb
HHObfgCut74XH8xf8jXUJRwPOThxSQe57Kg+eqvtZvO46Kim30YaXa0BANJztKeMknBgs9qOt3nu
I5FBxStMga9GbqvWVkuVVPw8/AvCsCxMwAUfypvBkV93ElRjUsZAKhxHyztiWkKwT1ItSlfgSpH8
Dnc94qTcnjYgIS06R7V023djFXkqlaAVe+POmdVZIpx2ViKtKDHjYPvMtLUJxjBBoaMm8ftHJvp8
5HQOIP1GkbzQqMQFmU9DxCMwhKwt4UJDRqMoDMuZYiaJaJzBZ7/6jmgmKX6uMtb4P/QrRHV8RrYm
sjKjKPxqyP2Xv5kcNUw5j7SzbU5qthr5pUtQ4JyKxczFIIk3d48Dh5sFwDsd9kSfee4CrvKd+4CQ
D2yfHCW2zDXaAv7fXyARrr7Xg5TEuvFDbRnhVUqxptdWBKPzcA7ks9ipQdCNR6HGwA1OTE27cQ/Y
l9B8jFmDxPfAJLQMk5o52M8Lf9nzFUSJ5hJ6E9my23xa613SMUI2NUvLcB9rL9+cqxCG5U0hFoWE
ibBksbxVcdL5TMT2TgMoYmj9IQ0HNXnKA2hA3OtzJTaR0lXYdTl9vmVEL9OKchmcpC1zu57fdvx8
ZHwTGrln1ailZbSRXVIxFZ1lCC3h7iMcjLelF1KyiOyhChP0R5Vg9/gXNY6DOn1EPfI4iVgUbzoA
8VYOWdqPVRwD57rDWRFbb47qhddPgjhkl7aMcfGO7BmYnzRQt4EecjyrC22/4LWy9EMpsyunM54Y
/qwNTYK8jII94jnrJuOLSpLyGj5Rz6AEf6d4x7lvA4meZfFkgpDd+9ZTty5B5ZCSGBIt7pGQqUYS
VfSQoGQvf1T2BuDg7NzbCDvR6rH4Gr7RENloedAyIrwrZ6Hqutt0ZcoPDSZEqrDXKL5Ek/tXys5W
GjaDiJKeYJnsQfoO+oIoodhwfrBW7jqZhI87dFz5l4HeAGsnrnTn4ibABX1lGy21yss8y9Ulvvyu
5f3OlCYpEIIgQWwOc/42m1a9T4iA6lc9sTtvBt11z2u12nPdNVXF39sV/ayqyQUZxTKV7Ze0U9Vn
fH2qbFq5WsIUUIDF8f8Zy6d+OoC9lzyY7U2B3eoyyRWWilwcsN7+wFH6a5PIY4FkJOXkQyVIA8kH
MOKlx41spLf4OB8MdTabR8rrT2VgQ3z6bjkxFIfA3eY0im/kRN2UuwHDgVt+OKjbDYhfi3sFdbpF
c+Pm9ajk/ji1kTFou0lCcd0C1GnCNYZBIhTeuZR/tnF373/ZhJay5qccRablU9g8Wkiz4o2gH6ag
vTAoF0oAGSgB+afQmef/2bg45EWMcNw6NuNcW9F8QQ0nlHd/DZwDPmw/DhqIS2FfoH5mkG4pKijb
YGK6jngVcEhFjkvSpEN+bLyc46XqAQXkyygAQgh+AU4jMZoWXJ8UZvuGtF31jYhEgnSiOYvzXavg
yc7rE1l8KCkQd8kGO3z/UbpyNvGP1GQ7e0/n1w9z362ABJUyCS1Sadym0DkLnq8PXxWlMgU+qXSg
HFT8TR+LVwAnKbEhb4WHgU6OKqDSs++ZThVJ8Wbk5zvNJEUzlaObKHvpbzI2zev0zI2bJjYpSAVx
x6hsCc7HsqJQGNflSXHPCxOp2suc819sESXt6nFr55d0mD+Cs7zWI7drt2PxuVrMEfaW/2GaeDJ1
2xWPgmt1XZCocEGYXYi5rS7tCX7LoOdWKgJmtxNomxu6J64sfy2BE9huDqZklLEu2gWOPP0rNw8C
HVrdm7Y8bHn8y6ZMxVMe2RcuqbsI7Eu2daqIyeNF1T1E/sn9Kob5nTIYbYJf0tkFKIfXevrfi2xD
4bmADYLX5jzeBP3jLf7PwqF6Qv9vG0Xq5MB3vTZcKLuRvXbq3c8WBBs9qdAknHeQmx/kIqkJpuSg
7uTw7qBPfPzqzKBwkQTPiRBgWV4dIwIJy/JovdIt6PHsktm+TdGL2tnMqZH8e0r55knUYwXsMI7V
waFeUIk5eJJCc4U4S72nf3WHr0/RA/0WteKNVhBDPwRydDxz2Pqf0Ws29qXBB4Oto+vBUvuQbWfG
s+yklOsPDyvis6MRERF6xzBSS+/o9IxgW2WgwSZaElbiDGjhKQfgBtJSBGrQpxy0NXKGEBn0XF2u
VBPgw/OBxjYLfBIcEU2pNd81OCx9epIDfS+wcQYfQgGe+wJy24sI41+ZbI70EwDOGhQ5ibC3MmGZ
rLeGckplTlwP1Rl97bOmLxgScxw9i5j1wL5SVRb6uA/wve378cDBt5nA4hS/5dSL+igiS6gsvWly
AuHDieDJWPrkzCLXoOXfUC0q02+T4iVKfOTAKk2lZ0+yQYSXXi0gI86IZwX3J20mjj4yxBQtsnmJ
JBPo0b3RO2MizovFQuCzNLWmO0ZJOTczYHvUghCtTkPxh1l2UXmfvR2YkvqgVkqBNpd2BB69HU27
pS2OZvJb3AtiSqJpE+ypxphqVPb5d2xM4xqk21HIf77tMnJCRFOSheprQJxMxCBJheIRzW1U6Qqq
Jq5Ck1SfwnPvrqg/MtzbuD02BPH+yHtwxwO9Vq/sOYQJV8ybbe8OqbfvViL8WKx6hwTIjtC0PCBO
CT1kQkOGk+pGpN2iHhhGS87E/B0DwdG96X6yqsDQ1lhzEOMPJ7emLx8NfK7E40Z0OCwmB5YP/K8l
BSQMKsVRXC3f35c7hvPNjmv/GsfzUPB/cm1SfdYwlKeC33fG9KUHYAG8+DPMax/+f99yiFVq2BqF
kMWnw5X7oeMWPeNVt+2scywT988lLyqBdQCoUTuPWCBXF7jd6W2PKULoW7zNEFKJUnDs4pfWcfAY
SIEpJViSoLA/17k6IBN6POHrNr6pdQKXU5gAdNreT4mXf0ZtNNsuKggOEAaq6DVHdGleul3YIVtw
ILl+Jz5n7QDQUspQ6l18Hy0ybDV+pwl3151jelQJ5oz1hwKdWfLfjOvJS6l5mGgkEQkjq1md7Wbr
IeIYewbLG1TviQCk8zwgPTu/N9w9EjHhHx9Gv8gAjpNKy/iVLAtcvkyUtL8k1f8Tcas2riKYspFO
flmUG/vyvVJGKhKFJNyXxAx9QptJfkolN2DrfBHAoma2/+SVq3dqUo/r1ZJhAo4JGWj9c/FHXWT6
0i9D23POw5eq8J6E2TXRPC45vEixydyhLvdDaifjPQOL/aImXXoArCPLuFDc+/+kDPBWDwUrf32g
znxW1ES4tYGFrcec5Usv/FMeaPxYsO0r9qTrbm3QQqz3SAiOP0kp5HIPf+PrMIYdKG0OQp7gg5t6
uQZAaGy2xa/dexvvWBR+z/Ft/38+/bBRkiwlfYfMJUPY/GfoZ6DZLzC6nCbWuGHXMNJf98JbB81Z
XfosfiDFh+fnOu1Bwu62BBIcp9Ako4ov7VItXKwLtB+cluLdF9xp8ZXSp7l2L0umj0VJzAorJYXw
wqiVqM98bzbh9hhpehukAXuwXequvVQAwqu0uzjIkT+7CF0hhIlKKcvcey2w2yHfF1yOeAxF0dnB
xSo1YYb9bO/Jqn69YFnmVOoqMzxOjFUOAjiPZA4/LU8WaQo3JNR/TuDU7gq3DZevy9bXD0XIz7uf
Y6P6AZgSWJ/WHDSO2Ypk4Of23gs++SRfkpWv3+RmJYLLho3o2w1Uicg4QYlXXkr+gZB5qXnFnuab
MZyK0dkIo0vsgqxZjqs7jMZkbytK3e0V2FAgDUfqH22hlRAH2J9O9mlCpJnBjHZWwGCzFGm+8d1g
P6anARWAnMryZt07MjE1OteL1cMnXPaQ+rE+k4L6H2/tdnqP78jrKDlH1Pde3/vgBaHvMOfQ5WDM
DDok8DGY6mA0TS6kuw9RzfPHee5PeZaYJFw745Tg+xqKKZ/L+7M3/Pu6tCOuB0uuX0sntmAHeuMs
jsJ/xyoaZ0KD8DtE5ajkVIeMVko5F6i+C7JnNfu065bnm3m0TnKg2BWIYM5YBljOswiT0kgN4zRs
RkxFvJEKfgAX1gq3ulJfM3s36DEZ6XiMHTEcP+rYchhll4dtl2UiUIZIW+TJkZ2T42vw6rkkIQpM
vdzmBNvKIWoz7y0q4AF51bQw5g1Sjw+x4jcM1dloquVGCLOfkATFl2E/FXaeGkC9akgn2i/CzE0+
uEjtLaoJhGdPsTzgQAlrxxK3O97pvcndNHwvUpuAv8GL9Buly+8lY4US85CvkyOykOrK6XF4EqgZ
jlf0K4Fvctq840Th39j3GEOCu659twHoMpEdY5n56CiqAZweF9aWm4Q2trmwY8MG4ZU3Ve69PHs1
CJ6J56hJA9+bscBRLhUR1W9HKlxgTfJ54ZnKzMx3qGROU9awZg4VcrGJLE9BRtUxtELV4bqIukrI
RHH4fxfxVLwpSsA1XaMZr5KLTISd6Zy/cwR4dKRlyFv8QK2Iytc7b/GguaoXJKn8dGt4YATkOi22
HGveBURmDFp6zsEHO05nYiXBnoWVyVkgq6n2GTnMo8T0Eu3p5cT/4tWFuAkgXaxIuDUMtFsRyg2U
U/TGtE/RU8zKkpWQofVaHZwdsmlz7iiEpVFuehT4IUesxrVWbPlMX+GNA+DvBcg+CZNA1/Ld200S
bo9XZ8V/yqukycr/oz28aj15Rn1ejpR7U/CkhCQdUr0HVWkD/46itpVQQhKhnCcCYCWhyKllNQIL
a/cFJy6pqjnlFCCw92HkiZAriFG8i6xwH0dYe8N6dHZuuecF+5FqL1pKNHCkCZUXqD0+zkm7VoXf
4BwD33jMk/DH6ChqFn2CzQczIy9aan/undUrKku1oVmaSJndldkJOWhPOvJ3WeyjE9w8BWSqKzXW
fqsb74oOOBtjNDCJMA9GBvpgj3rfP73MF310xDuceJlKvuPFOBBh13k4jBDFjjMf+cEIU71c9m7q
Hm4yWXKiYDMe4b/amghGsduxCL/v2Gy065TX2O+Olywf2WiatuZQOOIIWKBkdLEw6buRHJS2OK9b
/RXjMrEhevazIHiPqA5Mzwt7Zd8gLYaAnFWIsD3zvFV701+9yCF8/R3YMIwOBMMscXBFQ58K8CyF
wDxSfRdk+P0POriBtjVIUizMlcuYF4PlXeAjtXbM9om0BTivouLGIFzXmpeBzxFEGwVdoCIQKA/A
kHT5OyQNnJF3DU28l7ip3whp5n7UvolRqWvAVY33CjGLHr1hbYw5nM1q3ZQmc2+vf//sVitYXyH5
UkBNrPVg3uqhz65TDt3M5sY3ohcLAq6c/oAx5MenmZZwBe5+WpWXTNwoILQVZEA5oPVLLolGBEfZ
zlpf/5hKvNIoBsY7yHfJhdSesI7CdddCsYhYioP18ObLhzY6HNa9uu9/2hCeiqf59LrFlTo0MaNv
NXwRhBInfqORWH2jinPf1EZna+f0mmw5qZriMZbJsoIV+RuUce4M+4IJ1efK/vMBTX9xbxkPmOrg
b0C2RqJdxMEbL+UKuNSlzkPmPlDHHQJv6y8iVuSFMHyb88NF6wIjaAxU+yaDAqJh4BEoWlyMFADk
Vl9suFYP47ZjzUG+bZNufr/sKdB/PbSDdwKz+H3jpR/kuBW8m28vBK9DTdtpKiGJZn5qMHPPJVmz
ZS/Gm9orlBOuP6mtQsYBp2SXmLOwf8nEuJtEDiwb0kD8Ms7AWptlAjXY4JyjF8dyX6XNVmm3ermk
9X1qb9jFlqHfkEgGuxcHmP198iC8LIUY7CECXsaCR6F/TGhuFT//idcoFVM+4Z/bVZ0Yd0Amr8yK
uR4Wm8aWKtC/2RjCAhFEkXg++18xhstaMs0qz5vgkhyHVwdX6vVF/Dn3v4wRcMe47wHWvAGt9vaz
u6zhgc7wIKQ1arcZu1wlQmPAKgc2pxDsxfj49w2GooiP2FJiHm6idQjzq9IQBI5uYu6psWPQWzQx
A8uHXSTbOy3mlTE9rdp47DNNDLac4dlzT2t/W/NxaeZOz2QtmGTIaMnDUAoDQZfKAeYCLENJNzOt
2vuML3lywGBu47mNVS3bZ2lVOdOhYoc2cTgkebKYR7A0XZ1M76y5DCtHSjIpg++9pnUPYQECgcMs
60e+YJenFIBiT4XFnmgQOi6jjPCV5qfx5S2d8Nw78wnHR0kveX6ETCKwk0UktGaN7wH47nxP0QLf
YMhmTE2Oh3je5WxiQGDaP9SwwDrvhCRBv0wzyIVlaZLXYZID044ikLzzJ8X9xov9w/bRJYHBKKG/
18ZZPO7edmj5eFmYMEzmWIz7Eu28a15v2eOSima5J2xekgn9FfecFtGsk4trjLWD+QkxUe4iBUFN
qixZ71oPbHb9SSwsyoIPz4u1FzXoAkqeEc6kCCZZvylLPkPrApndbgSKllfIJ49pTbFuYV1VdqF7
OEMWCizdxirYpzIZljGdYQEFW2VXZNoNJfspG42ilta4yK0a2Ick6HEf9BoTpQfvwBgOHwnsO6ne
l2Z/7aD+R+qsykZZlgehMi1EgzlHTNixTEEECizN1EpGKvg5O90idjLoJL6smfk9qr9nCgfUXLX1
uiRsWmUK+asMyrYU9nV7I4af39vE6zb19tgZA5Ud6oqbHDYybsvXG4c0vPnHpBlMGEJEqNdq1p6O
rOliQcS3C5Er+lPLmMrzX4dy1ly7lrTvli6QAsuUgBpMA/w9FiVfOjYzvd2PMlK3Mm/lRwukiime
peZvQltZzb5Pn70AgmZkNEfCWFHhx/tZDC1RcPcHrF/ZT8J5Kh9cbRk3NVbAoFzZ7jDKDGHmoq1+
oco1MSasnbRqQlHPnbjbBrl7XtXnlZIS2KFomq8A/doYtOI4kGYC1ROSaVW2xsCYnA/CiQdmFqdS
3KaE7olAb/5+eUp/waPOm4njtLzQnOpZAP9nAxj8TvXqXIdnb6a7EwLApctYl1M3Bfmnjw3ET6+k
SmmBYTnUEnMIr0a3lAkEGkOw8RxMy/pg6FShSoZrKJAXFYGzlobaZ3AdHnFIb94iDPg0L/5lSkhg
nGANNENQW4qx7nU0t3WGy30xtr4HjeTJz27oAQWE9W80vSZV2IlA3thw1/Y/yI2EOUWT2a6Pg8i2
GVzrjXZxKeqy4BU4RHMyyfPhFnrPBpr+5CpRBbDykhTqxTaHlapDgCeZt6oBbqV7N5Hx7+i+PiwE
YU0AKt4fJ/soakDQvAukgA/HYWufe19oNHfUv06VZNPg1ir3S2QH2SsKoylqZ3IuNApaevJTDTiB
hIvhBgN0DF+XpWUwRHaqvKHgYCDGjAjoPWPjWCRaMFVJqbsUSh3ON1iUuJSeLiAhZKOi9iacDJmm
clXozDzI+pov3qc4T6Hr/TjhS1ZVsEHXKY5MXPMDc/oHKRdRGo9oU90jqfXw62HACC3Tc8dqGG67
p9S+z+wddstlXJfcbjaCMSWa+p20xhbZPCXQVpdgxpFfKBWCobf4EXiDTbw2GemjCNyOhzJy9k5H
bNqfEUG1J31zwPtJtyCtf3nZXbtdLQbDJpmTGS8xoI/gbvBgyrbVXT+4GULzVTI4L2KIIbjl567I
4LdUwluKE5zV1IaPsb19My/FotTO0A3X3Zmxz3vRMdQ3Doj0yvvrrtleamUjQBQBQ/mw12OPcU2k
dQgHyCa/WlyVaOhmkuH5+CBIe9K2daRmlXMfWcR5xsoNWIVW2oi8LNNP2lG6MHBNcS9yXDujIgZi
tWkb/gfIU9rccme98TRzRsW9xE2I+HL/rKDYTWY7Q09ndTGpPSNDblrcXsQYxwnPwcQrqoajsmiJ
GWRsDf04uqHfAHSZBmEOSuvmYqNYApGAkY+q4bf53OEFYZwXqyhTdBuT4oO4PGC/LzBVvLX+kG+b
p5XP4WvgDrpc1LvC30wOMqj4SB5wBnV9SiCX2H1knWokVeBt8ZC1nevQHPbqdDbSyb2onO/XZ4hC
uez9m1mu7Z6mPaPGlKzlo1/8hbXH5O7kWMKGlVQFNqb8VsZ2ryCW6pKgo9QoG+pPUs+g1Sem3gks
e5cchg77K6Ut704ow5bfvD7rH/U9eZky6TpFld6wm5XuMIeUGXk980eNYgvSLg7uV8VKIJXYZ7FS
EuL56h5tKHXg1OKnPsqkDU6JoR2+imz6SlhbHZuL/EljHz/sk+mu+Z84yzUjYdWtCBeZr0BOu590
DPQzs59Txae5I9Xjph7MtpEFEJlj7bDsQ4glrycR39NBsMy9lwFR5w+c4JWlOC/uoJOPhq/rtRVb
w09EL8CY5cIuFTuuiVNc5RuGaHX7ncSGbfiUdEhMciCkXtPKL2vRxXFb2mVwzFdUOOkAAPStQ6KY
RDT/YVIjWTrZh27iVpNe9AU2WeN941humyiWx07UmUzVUYmUXI9eylUTQbr9akuCOz0QtjKz96pd
zeNWv82X5oep0Drp38Qs3iHgfmUrrR4R9nvwMuu4HZAGhFS61R7B9D2B4rMdQMDeXe02xOy13UV1
JyYunPZ8LgNGtVM6aydoD1XhdBPxeO7CJHj9PL0jAhSOBD3tLnHmu6Lf+BEoZyoQsBmHEGLSdW/O
BfWFp15SRRjU6o6qpT5GxAirhrpoj4ZH3hypAT+DyUJ2E5f3xNTd80+APIK6+Uhasyp9Edoc2MjD
zh/daydyIUSmnGUySZeXrmQm4Uge1NVk06eKBddeFrC+Vrrc63sGTHzwe6NnwIivdgEmB/y8DFuY
1DR7dGaQVvn9Z0r3jlfrUyHCJfk5tWCelJjcio+pf3DkJt9lkDXES3obL4uOQdhuq2MUh2PZA9ZY
qS3kiJI022JTbFGbq3ayoqFZWbHR3I0IcYU6hgQj/pqWHN7gvo81QyVFTiK41UvQvp3sm3qiKFjK
Sg/namnVMoKx5m1OymjkmlMMjOGTiyzUFBeUIeSV2+dMXjg+k7wVTlFFLsr/LkKn6QdoWj6YLmY/
P5vE2kPaOJKD+Q8uy8EmbrpYLX0PS87E30QiJextmY1v/c8We5vUN/EcnOa2c4gv1nqnrCMS9syU
c25eLcQtlfe0qwfiO8bl0cYhMVn2dZIONRWPBUf85N4OK62Ky1i8FYcHrixuzHHHmvZtbnZaV8+Z
qUC/aFl+DnP+2etwgzxXHXLMWM7RtO4+DITqTXjs7OSqXO/N5pxJCzfwP2ZUXZno0v9FXzUa5wqk
sH7ICnAlqDEFIwRPBWaWbJdRV6VoE/XdmeoJy+UIRu8ue0EOiS+XpuVdWXihpSD+tUbUOHAFg3Qm
GSHSCnl3pgak4cV3xxTyP8oflqgYnWIPObvJImW6lAYUjPvrClzpJRcNp85jNuye/DHrvVH+zxVq
iusXI+/UJK9yEORujttOldTQyv8jXhZ4DQHxi1yVnKyikmNTHnMgkotb/Y0DXUoE0C5/K7VGi3x/
ghitANnYQIN93TvGn+CPmEqfSihmEbswkuyagmlDaRUONwFpmSJDFJ4+tXdpiQ6+dmeAS+ALKamk
vvwiVPzl+e0OgFY8pKjf/UpPHwwDE4xSEQrvC0+fVaGqYDHjnP1sW5Avjgnb+Qg25ITLsNhiJBhm
DPyafinTzV+CKljqcGszaMsraO8M1Iq/PSl46B6uxBParMiT2DCm9j8z3ca+VerJi8MNnuteCwG1
iSphEtSxMByE+i5eWFEcshb707MkLvVMWuRGRjBr8Jlvd31/bKNYKuBzLINOFeJOERFq5n0s/Zca
+C1y9CGd8rpT5TYpcmEK6kzdhfVzoRcqfkjaTU8Xx6NDDyi6hFYmSHNIUZCSSOcy9qlBngmyr+QS
vmISG1eOjLTmNbsH5ipKBWL+8ETyGQsQ0yCWtKDRlEG/jK7x5Kslbv09ykpP7uwwOnjsOwV9mQxq
MlSuW2BqX0OiLY556bXx8p/2W/FUV6XzuPJnhSzvGFsi8Eoy4TM7a3f6bLuG6OFTk80aue95Ynf4
o0qARiVPDownFDTYp26Rxh3RGETPw6rQ7c9iQ+lJ0HWWNxve9w6t9sasOY0sBobE8VDg5BEmn1fI
M7pypO5y5/3e1k4irafoOX7AnDLOaACCAvqsL/b4zGQKNjs2RqG3ZVyBqcS9P6hBR5k3rWU2bE6z
IXkCChc3GaHQp5EPZG5TgTOjrKZbtum4SB7xShdBNDfIxvmOQ10pLIkoIs8pDupyAHErKdO1H/x/
q8INnjIDwjFq1sGIWOVf+i5fCVxNcjRO/6SzduFycTqs3T1sQr7I4cEsU3/udZENygxD+wOswgME
rnuBo5D4MoSn5G1jPOKI82gN6d5BzpgF9P/3KOyrMDrkqre9VCit6VMtARxgMWn8X9kpn8oFkka4
wy+l8zYwEeilDFfG3tMKpdNobR3SRKLSbK6W4V7hd8ytUwZfZoaRn7DZ8/SX8svKCXerYHq1ur3I
Chvd02vxKrEvrfDd0MXkES5o/gq8IbXYVypkp0LjZzGkDu6KMf8+56aI0htBL1nImOQTqcN9587Y
RjKDF92LyBNgKBW1TIPmxhUhqbzgd3444mSsknDwQXrzAmrHc1qKRRgS1gRLqZqg6eJnBX9mJu3h
yOnBUjyEgo89cIUkT+dKXsORtOV08dlV0UUhfoagdbI8DvhvBf4eLBz/zwlgT/ICp8PdLe53c91t
4d8C8Ks3Q6V36ieuAK6B0gsWulhuUPWCjfhDspJGl09K+ikYR0436Ac1CnG90KAnZbTQ4XnHZ+FH
zBUAVSaF1w0lUtuGZnZ33eil9Rl3v5xDChlUe5c+Yml74Jak6e6JvnqdhiTVX+nMrXBIHsPxKhYo
+f09pBt2cxizdHKrlokysbn17SEadZDYlL/zs40VJ163b6xgsOiKtrx+pCG/znADE+aWd7dZj6Ue
kUoZMY36ItxTx+u2L7Fqq0XshxXvlXUR19C4lRQZx4qX6wIDry4uy8b7KrBAgoTof3eY7lSXoF+j
D6TpgAmlo7GkfQPd2bHLg0wK9ZjPNH0zMcwSRGn8emEz1MY/IVhrbwL6JxDyINMbZMtevHDvslO6
3FzuG22u7VG/UYtv6p+b3oQst+A0P7NZt3tZJnYIywh6DoofYg2S2eh4DjhAyDuQbL4wiq/Jb3dj
bQqTtCX06lbQlqhxlai0Y4oVN+0ITTRMFxz7xu6lbygGzYS9SBmVVAWxBWuGEUzi6L3V9A6eX/ot
+PKkHelOLt+D974ixzFDZqbx4OeoJFNQjlsMS81WxWeF3yYXr7QVnBkBcHCso04HwHDLjPEHr4ZH
nUvWI8WUo8loD5t4OVg93vojiPlEdoLKBQvjkVhiqTrnPFqEj8OeHyaPlo0llBDSUslwIv2mlkub
AxFiePvZbqNHCw7KXbomZqiJwr5cPQPz9139PIrcA4VXrtsD6ZZTx4g/6yuzQ1KmG/lIXQwAXX0z
liUxUIq+CfJr0X26uCJGSUaCbPA7cpVQECixYqIIobniSjCv+NtVf3shEmeYLQfzNjEWS3rMlQKP
PD1n6r4ywpdpcDQSvG9twjsASA/2VsplzaJ902Fx3K7tTS79alYwaNB4SNHEN6L/32Olpuine4N1
SHHL9UH6H1bw7FgDriUYRNRRctTG1zzFtzHGF057TN9FbTRjgI8KISaf7Xi9RTJDx1AOcrz3AT32
EXE3/BkXDV50jJTc8C7RH+1LifiE0jMOqM1tLG+lw6quFETCUo+Q7iMmXBL/Pb3U4RFSIwE9aSnD
h3VaVF6mLtlaFgXcV4dA1IKhaVLNzIJkSUhZ2/Y5qvP2XseSlTadi2AGedtafNtafe76FFrr8odC
MiSrfBC/TsLXcDxCQoPHwZlNQebImOmZeiIkknjlsJ7Lw5vytVzZuElKfcr8duCrcSWYRkXnrX2z
PDG+xTLALTd9WpFfEuKrVksRQxvwwH6mV1IPn7fsY4ofhd1/BuDw9lQbkXk7bNLX2MKodK5VEi4i
iWQMsuIZaKY6HROzMefaviKWIX5PofAxY4QsP4BbcxEFeDWHiK1coaQ+nW+yxxFnmtd/DU2tvUvY
rLsxY3tgm2cWS0YkedCJAQH/3ww5Ku1qZxTCyzDiRcjxZcfPGSI/s4eNsDIEp4+4HyCHHaiFGYS8
UD8jTCZBGwxHTFKXm8I4Zm1oY0IoHF0dQBtwB0AIats5Ym5sw9RFUDzccMJcmWo2ln8bgXC+JHPh
KwwrBE+My1L8cVd35o8CjD7M2gDiKboD40qN1hYZGC/irDgFgHclROENtuHZ8OOOfF93LfXHNpOR
2xnyD4SxUGT7ydhgivBsN5y/pX6iS7UDyutDZtF9xVtkED8R1dwwwcrhNzcCa8EVI9ATNTB5Kacr
p5l+IZl9lo7HFi9tZ3hXMQO0ZFaOCyz3WnE4XhRh59bUXj8xcpYlxKT352F+X0BckHyu22WjaepX
xFKWm9fnS7hga+msJ91bjYqdtYbDGP5WqNnKcbt7UQ8k9X0oXf5YEyLoNfE02vhmdA3fhMyIvSj9
9Uubhgpc0vaYOS0o/YxSHBnLmOTfprlQTt2Bs+7kVSs8wSZR81vTWRQW53VUg2GA9KNOsWsabRw/
9EPutjIFfhYyFvvgT2o6MTcXbb7yQS6HoGa1iebg45NAMCVZ73fEN1+UaZSR3fyyu97apf6Jke2u
KzZaBFS2TnSqFqOTjy1NegycZYoNBHEgt2HT8ryOTOtl0fVmGG9cnOxvUE/+vz/xk306lGqlmOIW
7FRUt/y+zsAY9aR8rUwuGi8lIojth0RnVPEA0VGxDu03iFN5VgCoTChiDMJRbcrzv4h1oEbKHbxH
eh4hJEGoaM9uVQ5e2rir77jJ9wDXBsFBNeKURKMvcmsB6t+H3MY4HtGf3PXokNPBT7/6WxbvfVxf
7ccfQ2SHNr1n8ze70y8Lsbszleyuerh5N9ofb6PGNDTb67TJYKeh2sSP0Ixhf2ZU+ayG+LqYZPIU
6HhIlcsSw2UKN2VheQk5Mnbsdgya3qV/fq392Q5iXWYqTNCb2w4AIMAqQ37jxkdTbRQ5DzMd9LvF
Tgn+/6zw2EldQnvEsK16owVmkRt5p/olvVBkpUIFHxk8Pg/JVcBQkmB4WxwCPqm98Feo53Un/rkX
5I2+S9/LDhEMOOT4IMdEhJO4eSM7Lyp+GPH0r40HDMZDnAjNnYdGgeQF6HDSgtrFYsc+FjrmXRVB
PdkMBgy4mRMr1W/ktD34sf2OYwHD5DvvRlYfHXLl/XAYw+jr4oZ3DTDhXShEsioy4Yd8zYjIZUju
dSEGidro3ATEctYeO7F7AxjcE8AW/bqRntzwAjrFucwYcjnD6/43ItXeyFvkmjUe5nVW5BPj/doB
ovhtCJ7YaB8Eb6ovZY+owjkYobtRCrFQDZxmsUCunwrZ1WiKmMQ29JnS4r2gyWEiyu1zfYTVwfN7
BPT5fK9ak0a+6rRIUC6xJvcVkuT/TFVxJOX2NM4XVzC9in++MjBJSVCyEyTjkP2IYrWs5sHXIXRy
UJCarQC0Tmk1+EC3qJZ+AZ1iNNeURBJztfZqXKqcgtxVvbQu25Lw5yOJprElZc7HUgBHFGSsjxW/
0QlMAvcBczVBBCcqUYEcY4Xt6zc/kcOiC94w4o2PfSle3+6uhoW5oSzg764vIJR+YXJg6gNaiVe6
f0O35R6mrT4uFVjxT+Jzj5bpaOpDDJOGUc+Lg3rpi8Xy+RolKqApcGW2KxpYY7r0j2dh/MAcdSFp
QVKPJp31kYVY28CmmY81d83ADIBYcxwwPC27x0E+rRUUEGOUm5qaerQ7XMgqWYDSULK0XQc8STIE
RLlvjNTTdFytLDeJTbqPxXRuZIske7uppp2H/jCSQpGb+zzp2XOl57tB9PCU1gveP4w40thKqNAG
DhP8rtmwo+K59wmVjRfcK15b/eFaedzyx1ZIu2RIAgdnNdKUYBnYWO5q2s0dCGDDCmZ9VQcmxkxD
AT0CEogKLeuwKikZ3OL5sFKD9nE+bKu4N3ZSEiL9yqxwZxm9fQVWczpiDld7Fp0lNBhTTpZdVKlA
YJ+MlmhEI+ojIrg9lXyfEMB0CqhcWwpxYkzKDh8B+SyAPIh7Ge5kC3vnEV24zEpRiTDQMipF6ct7
DnUl2MenTZdGupuoUC/X80pkio8vuRnjFhMlYgC5WeNmsgoGJ1xF5aqHkSIO76LZLlloe72G2bSl
AQf+DgqyG/vqoDhGBV/5Y5RG/G9BgWlYnwIG6KD/ZY84GZxScWDNvhaieaxZmTF2kh/CrE2pYV0V
AY2m5RX967IfOImBfvfyDnGvAgnUu1uWWMY1ZCelQ9FShxK54rjRYkZJjPpMFVBu+1UZiHtNhWz8
j/UX0Y9zBDfGSEZ89rutc4srBDTDnnJFNGX0nvV5plRX1OPOTH48Xd9dhpKyOB1qOKwMtIZpw1p9
QbqnUb90v1NPP/A/9Wc13f8x8EHjivL5tgdQ4mjB4NqttTaZH6CYBFupyuswcBW3rc6SEiqg/v19
BrPIZc/Y/BtShOr2DdWNKbjresnRct51w/vNfTUiRDJoCwLkHqOLf8hnCHYuorqMHMccABOsBJ0B
7kzk/cKxN9/EG3+Zm6auOk1SY7gfnNWeB52L44nH3roPTugh9+i/Bf8W0s9eLCM1EuVJ6f5Spcgl
Z48oPvQXRvJdgKgqf0pIl5HT2+7IJRsjEqzX9ApBFbho0aqSARrnlwBUcTyi2wr6OYRk/DofCXg0
Cj+aHxfHx1TGI3Y0B8YkkdnP0slXC8SgSYmg3iNnm9C6sL5bEn0IQ9r9+p0zyZudxwl11Jj0C4W0
F83Oxq97TK24rErgQX3h9nLSmkt7bHvyXzfEwraez7h2F9XDu9BoNYB6yIEidH4Ya12GaR/yjRye
h0/yEwnmspJcXHlh3TP05p/snF9NDNVnKSydrzaO5LtEVHfds7VIVC91/9l6pcPvWCwHj631cabS
paXg3QjVQ8Fvr4wUrg/NHLDfo10BcHtAf/imiKEXqIGW6Eiw3WmmvML5ucL4qy+I/qZO7BibxbC9
P4fTpNudiTm3NZwiPOGoHay8IpIpSxpSJUaiE6y1yry5FSOsuw5eaV39EcNQiKIbD7BfJzTwX3H9
D8HyFClxJsci0vFO6qedkNFrP/LXuyfgVWnns0N62lD3dTVJKl/cFq1cysTW89x0YedfqyvfIzmC
a2BXkPM6lzGd+U0QMrh7NyZ8bOrwIWXvvJbKRDDMjx2rQih6BPGnzlxOMKaUHmZKoGvr0iW9UfNg
pAH0eWHcDmo6zN97cnVHbrZs2IJFpm0cG1iNv79Qdyrit527DHplVf/Ihb4LoAII++lMuMZYNsCN
OG/IhkKOm41gbEqIMtgroQ77oyD+cr86z5+Tiu5g5oRzSp+f9mhsA7okhiaX0EyGvjpI1KmdQiBx
GPOOMRAU4FTt4qz7giIw5I6WbKfRU/HMhRj5wEQ072wEQZ2cEFQJttwhK5tKbEfhwOPEbJyJaZR0
CwcJg7MPdfMdbnm6hv/lO0Ovx1FWMNVeaWiPmWKq8qGOHjPuYQl5NaZb+t3i6vQ2uTC7ZHcHkVlg
60il7VhSnUN86s1CM9SWFlKCFqoSahuDMiF0498lfixTHq/Z2p0TIFcFoKG4LxuWApxEoTHGyGwQ
TSvSPRG7VzHTSIyRIl3XhpM9BomKuXtK4rv7+nI20TNWFnOyz7fUGh9ar6vzlYd0S98EutDZPxD8
rYXhRrtNYZ6sC/oTNdhtx7n5SLi4Sner4pYMBdfjkJC1VgJC2+3ew2aOtg2OtUt0VvO9F4dXpydO
F1vCr02yDto+eRZR8JziVS70knbqmuMHVaMBLsvZJKSd/jbGvcu7vMo5+aS18ob8mNgl9GzoR8pM
7+VSGgMZU3dyuffsTL4PSyx0q3sGlbaQyB+QuIWNECyZdcJAxRvhHcQpHkP5/rh7e1LjUejoqDFQ
oiEFoS7NNz6itbc1fndnjJdzN1Y+7dAi1AEtTcZGTcHgME9BvrfJ5/FqcpFFnAzONyEG7z5SuK1A
d+PN6adMbxhmImUCfzvJrb8VhyxBYe8THxRpbUoohT5W6j4TkY7ff8R+ncQ4xJuJOskQslPTVEwe
PkD5sNtcWGBMzJ8Qw+TZ06st9BV2RSrdLGh8NAYJjkjQ4/EArX9njaE8YGOGCFCJ3yaoxj20x8o6
wZtydxkWPlQbtyFycUZHZUh2MxhKdjoHb49E/qIKKpzi+Euq+Wo8K632ANdC6btKQzEQe2fa1H69
iXcRrQ6SeBZCZa21Ex0uWXEAYUYcl4fd/hcB3P4k5W14wNPEvA4W4xX9stUdj8X5Ze+flhsL4o/z
Q+hzuJNjGvAN3Atoqfc1B5LBlKokoD/XNO17dPdKzi/DEdypeohlxVaqmnwIElsFp2FXjwjsYGyr
hcCm/Jnr52g+x+9Ph40VlOiG29xKlUcKqUPH5YlnfzenTIxTLSZu/gnfOW9dcbIWYdZqrDMVHEH3
s2DE9HSC3HCRxDRc3reGOIvGbSbZNxO1xFfQtVjyfb2AekXBZn/RV0bLlF4gYyaDkpDkJ8ybeiIn
1Ak1gQ3D+7i+S/LI5Xs4bMDJ6AXyvcnP1rmu5+1Ed6aV8Ct/y4oQSMNzzt6gVQ7LAX6L2AO0fopG
pIV+JuITrM6v54M1H6bNik3Y753xJp9C1uRmLTOndbIC+9ud1wvoR51vCxdZQjjSqCpZzlDuW9J7
/f0NX9vrN8B/gxM6Hbj3eKjuvhYrS+VjGCXxG6WlQCy6Ziexl4yBPIaJ/DfKhDsRbXeFsNrCrey9
BOFfvaUD1ZDmWDNr3/4CirFcO0qgBSO+tJ2DwIsfJ6kU5H8Y9dHqNZ/ZcAY7Aa3OTs5LiO4Zp8Mh
2i5+9Z2QLZhgPsGu+LHgkRBjZcEBhilSns+HOjkDJwxc33YJE1n0ws9Ulir8XPyiB8sNfcti5f4P
wN0G2K1kn3/Cb2JPc9i1MjdlyPYJcbpcs6hIcY+TJPnAAtEMut5WG60FWUhFLyJiq9gcyXzw56X7
VYRLwn3WphDdiz4gDDYJei2SnPO0peTEGDnktVr/ZIefPSmivOXWpmdDjaNbDwtO88+UQ8CSDaL7
Pm8Q2Ev0plGMHwxaf/PEVnrhgMZgPDNvCMYs0zpKKfkPIbHdWs3bUwAEyaJ62SfxtN3rbqiJeACx
ZLW38tvcUVP6ngVKfZx0VUU+cERCBCP+hHsgFh/6h4dxMBCeT7gwRl9wl2l4sN6gtVjp7oWUs72n
oQGw5oPThlARf8PQVnnIO0WmB6MDwytXQkIpFfjJqEKT7MoO1P8XDK3UzwiMC92ZaBBn6BahYmPY
JnK4inH/qKu1T82C63TdHKA/0cAE+0C11Z6IOUSzvonQYLcJ8LtNb1SwS2ueLykn1Bk9ZuMMQg7w
OkGPrl/0TqeTJZZFCoszgM1tBMosbLLUq7pZaILtL/MIH/s5sLsXdy62cpdUhzwIGMLRDnI9CxgG
tMPhgqFNalPPgDoayQrgc9KvP2d0mbKq2MMa6sROSOyqIi81c7Cw3cRsVLuSS9fXGgxIU1v9olTB
AVbUwHxmKfvx6uJpOhskgoD3wXJ7CvjjnO7iuUdQWK42/WTGky2yR91cVsqxp2Sv/Io4DoyhOLyZ
w0DxHxpQMmRikz0+UJSyjHo6JIKnCmivARGT4Z6zKtb6E4dPyi9gM73zHwXWs5gmCnTgaNEj7WCH
/ViQXc5fwFgFP89cy/qndOluunc6ro6rdQD9L0wqV4MbWhhylIcbs/ILYiQcYIbTdWDTO0hXtLnP
0KnRr4Cay2Lje3XLTPcUap1QGYQ0o+v7XT77TrhCy3djOtx3AMNT1mGzdeIp0g6RBYy6/xjCPcj9
ay5eBpuC6HhD7hMv7fwgTnS5vwqvEu+Q4NCGMWifGXcbhAqI2QKjuAWqSLTojfc9v9KLQ6sOcSF0
K3AUFe9nIGwgjX9dhxLgm9bHc0pMoBYbSZ4/XHL+57ximnF2XEyvpL1eXbo6S5XO9SaqmlskyLcE
kSwZJPzYlhhkGHcxvsMETbEUwB/mxcifY7VwYVTdLfqQmY7g4NGjtL++oC2i5nZ9QH515/rdT4tB
uLkpsQdtelne5xLmEkGhCKhz54ZYZS5SzPverxy7a7S0aK1UrP0sN6jsPr4jlueMfFr5jaGg7uW7
/L7wYaPOAc4Q1q51bXqfaRKDiccdopI94WTcODAKcA8VVNrhDS5FDhj/5UxvVEhgcZjoYBowWCn4
CNP3sCW2zJUSyu1XZ4b35aht04zcmga0Par3X01RN+HBbfx9giUaf24JdDrLPvYoGbn9fMf4HxP1
qNfvvgVWnc64+d0pgYprBprAm9Ubo+5M3Ra2Y2Z4RkOkqLGxrKzCI//s6G6K4hgpQB6qLRJQLVsV
/rOmHzZ8IRcrGSvoJhOtLMfh645ywJd2llldLwBH4GUfnUTEcMo3if0PZAqcZiGcq5WIw3igF6Ce
4iJ5Bb9Dwh0R0MAuLZoeBIHBsnoFloJq3+FsTq0CQvop4hLXJo2nvTOJofXxY1bbCrd5G/NDD5hv
3lvwymu9TGzLtpFyHlwvba+4V7yf0R8sJfoEZZpgEwEKa103eidegQqVbV9yiYjrFL2zu37C5efm
4TWWDTS7RAnTBjzWd517wJ5QlkZt812tgOH/ZEO8VwPWcn6w1oLv6mnn01m0jtm/ffHGRXv5QHm/
DSjBfvFirVG1mwSqzP7NM1QdLg9whzq8bqREOLRqRqWcwsixVhLbMq1MzJ0/86tGxw9zspVSyH1z
USqr89dJJB79OCGIzO7e/MhviwbtcGeU6QMIe+6G41nzaZksF42vTufPJF59/Bs3OiMd9OAGalzw
RphVhRM+9HFnltF0ge+af5ditpMAX7dWbKKt84b7Eqxd5TbBPleTFEhbOa1AIjXapR6uYLERwAfj
TpuKPreT3Ge/pgr3+BMhqs0EJgd9Qs1ydoVMXbZ9csFNoNnz9hlJjVCbdyiv23kxntJUlMb5BKlj
RH83YVDrhE3anZYv3UMa4d+0eYknxvUjilkcU8wpSm4zci8YdTYEE1rm83HooV4EXop5o3aL8HP6
L9Sd3g1tZNmrWwpay5A0D+nXta2rbbqdPuCh9i7d5Tzt2gKbT3ysYHzWXnVDevr4HUib8t5SGFnL
jLNpFKJ62HKga+f4UpT6IDEXYOrjW6YNoVSKH3FAZgEIp3GiULqv/SF+0R7VJMyxuS+8rAqFHBf8
gom1CdQz+glqm8rL9jySiFXGIn38cMIvH0SuhBeAhCQ2w5BOU9ey7qtbr1Ov6t2M75N+osNfhVcL
hJ3RFVmBWRmGiDMCItHSL17knMF3FQX6+KC+o1Osv2EkNaAj7kPutRYDrxvK4FIa/jZYMCLnCqiw
LzvovUSEne/ZTTmwuUoao9sD5HVqmVSFFe29Ebw6GF/0LUpy3tyoTHdxEVzL3M4AheGNuja/hmQW
Ol073QXtgpgylG1dMXLcomY9PWMBFYe1JmhxcvNNFnlhES+8QymhtUCINgUDfNed4fXmmqDZsv85
t4avEUeMSWInEdIqNfclvPM3kXuE8GkWyiKv3CypkNnc7DfwitayDFHhhnwNah5GpW+oadyjXFAl
0L6GgSrjt/2jMu2u9cHHgxgUoMO4vkuQoOBuuWY/xnVFnRVUGgoSwWK5YxpBwazZfp9Wb6Fo2Z7J
MTUg0dL/uMBak9BK7RgQMtlloRbX52dwDeztLANx/sY2NxOzkPbtnEN9YMvsFIfiT0HcaYle5y1g
mFo6L1bU3jJi9Du/BOAjK/J3K+N35rKSymoE3zhV/yNguS1IPUC65dD1cAnSNrxYKJVjND/xO3Cr
GHIS8EjOeQa/Ri1UpX5S9DIza0Zlb5BMdwsp4MjhJioLpRee1XQB4Wbgta/yKiq7PDjzfAX3SQ6E
+cl/QLeU1s1wPv500hnyE6+9GjWNT8JUnD6cPWEfRUMlMrVzAEpqCRRjXoxihtivKoIpWQVYWjes
Vez8EZNwTSjA79/V21quQNbA+FzrWsz52glWjv+5N8AQxbqVOv9JAAff4QYB9+C5flRX6sWqV3p1
jNrMB5+2YYtx7l30fvUHyo84sZj5KNADWQmFbQCKr/vJpRCof4fnS5xw4HixHOlpE9Nbj/sKkqEh
Vd/McPUmA0ciaOC0i/6Gxa6BVIM604EEZd8TYpU2p2r+a4w6MvvsdJKaBTIMuwtkYJ9nLz9prHbN
D/BO9lQOK9HP9jXneUOjPtKKnvyrGaRnBVKUZy/bcZGLn7g89EMJtmUaweQEY4vpRla2ABJA0Zuw
gRXFWd46KKCRgfw+k4pf1H+Sx0MYxYnwJFSZUcqwRj5mul3GNQehf6ObVCMUnMu/RrJarHfDjpez
ZZAwfmJAvfKehBMYHXvPHo2KV1BdkIZxsOe+4fECaQFXhAOMRYSMFQCEvgG5b3XgdJ5pnl8qVdEW
oOHy6MWl/LMVNB4ur249S75wyFlKROPa87HB+DoY5oC7fDRnXyQ3sRXK96khjqFn/KiNHuqow3xK
lZciYjSadbwAh5Z9OweBlIZuNTmOypgMWQsgLRxr1YSeqnAcLN33edLW6Rd3RShrJ26aDm8X6EuV
IVPs9OX+dmCIp9pjexDA9LQOS7VXGiSOWUno1XUMDEpfD8c1YuAwUFXj4EgEEMKiesu2gG6DPtzY
eDdpeCFk2MjxzV/DZ4D8A4ZiapDOXfj+MobZUIGj8UWNKCo/3D3UkPESMd1qbwBM/InWMx29+QfS
WF41GBJnC/u80kL6knV4gQW1uIhF5tNjdrMTDkccxeJneB5eOOaNPt39fdFHTOY7XGFLbielQ2vp
OCr0agnSijJasuvqHVsbIXJa5UMwPw4aUdGvsbKHOTOEIVZ3vlSQnqrOpcHRm5kkZsOMuHrl+28M
i/ayD9EfH6N+PGWObRhfkVe1FZSHAkGlX04QgFhjyMQbkJT85IhszPJf3tV2P7cMsdAIzXPmy+0T
CqAycSO8ikijM20W+xc0jCXiA2REH3WEuW+RHGM/5JjNSBRxhnSI6Zuyw4xtUNQb6tHieCVDRGFo
pUdLfTwF4VANFZruG+bwxY4xztzV6sQGDohtmNNs1yEgfk62V9ehM1CuPCkjNAwn4pAKviZ6jICF
G9hAj+IdiMBNMIGYYmyxfeGYVmm7wEqCH78vVGLo3UDaYyuAKdfP6RHApCQGnkbp026Yk+bXxZI3
NEY8Y+opgRcgP/h7SaKtWm2DENkAAvzgQGJCfDlpG4b9Iprh1Way/d5GzPeQxPwxeXdS39OqC2Kl
48aswSxEDbdUbN8QAL3ycp77668+9M/gQ7K6nHLvBv8e0M9ARwFoRIEyNnTk2z/4y/ErFlMuVoKe
bUtojHiBEWKMA3v5cIqgIHX+si2h/PLGiGmak49rYcotLz4g+Exc0YgFniwd81llDYr/skNzGNAH
S+7cX9WT8ol1/pxdrXYrYsNriuKApYz828RT79Me+j8SltGt6vGN5F8pYjYwfK5aYdZxPGQVRmvY
4DBcw9LdD+dDKPgW4ogX60w5SDykpNB4qQFZ/0OLgn7Qg88OzZAIEIcdeDjXqalWnF6YeOvGWH8h
ERtIZR530WNxEWmCik4RVjFdMiTFP61RGDMCV4VydZxKchD3ui8/AHfha/kxTx3oB51aAKVIg29I
MbSkDQi0l4Fc3m9ilVIODzUa7UDii6oOUMnn65ABcKQYshLOEEyNS4achpNH0hvrvOTo9fqhsCL3
8r4hDnjiiJQwdIhNVCIIxMcVa/5CJCTSuWPL//xGwHxojjnepohZveW4MQfSrcGA43wBschxYzdD
efdn9FRLHGsrrzIZl6YLXNZXJXu03E28GlU++AGaRK4Ai0s93wsxrMzW4a34lBZpx8YwZQcpfHnd
SeYGF8ij9IQGh1fD56YLavv9fxqw2alYDQq3jsrIV+ZuKEP7WgVh4SxKXkbUIRHC+jMcycUZrKzk
x/chqZ/dl9q4Jb/Q21lb03fy0LLrc0Z9MIRqRVjlEqlZLjvejL2WlqX64WRGaO+yoJR41crS7/BL
a7BoQaBS5IfIByiawIi99JnKyOp8BKK3RZZN/HHyfBoePN0yJOP9fk8E/Ar5Csr9J0SyB43a06bi
/9qhOYzH04pcVRSZIcdKGRNfepr1eZ0X+KJZXGLPvN9Q1fJlSYMKE5tPVecr//pqi8s7P0KcU7iB
sqWj6O5cQpRCynR3BaKVY7/BrUn+sHd6PmPhsnYZccMCwLHTaHPbpfJ11f/5MgX3SMhURLliHflk
Pqpmoh3Qw5CZNIcp6/0Vr0Sszm85E62rrENKHHXkGB5dyo0KfrRr3nIMSdPBPW4mAE46rJd+Kiw2
vdQzPeEWOkbZNluaHK4LLKZ0DQOeB19ZEwOClhd+JrFYJIo+i632EneHc53gt8AdOyCanXluz3f1
URqxIp9WsZRfMKczCFrD8eqmKkGhMYVpXaPyQ1gnnia80ufJ1e7zm/xjTuTG6mOYrykq7XEgyReY
TZBctPef9KvrL7hG8TYBLlxN3cutRmpphiylZrRZDzSkGqDDQpFM4LttGO+N+747klr6qvsKHMZS
3Eb2pZpMIfdKCL1SxDbXK5bX6vlUsWngdyQCD3J7Sob9OUsxBB4Ui62LZykKpe6Vbbzq7ZblndQD
Rkery2QfiG18ywE6RjKXIs4v5qFHIbf/Al3z1xVk/HBK0NYc0/JhU+XU0f3CytBslAWLJWiuQAZj
xNHZzrdC/3AFS9ecZ3xqSJGPmfE7IH6KFiMWr5hrvYXDNX0/WSlVdNvxAwHopJclyep4EcRyOzsh
+l7ijpIMJRxBS7fdn0HVz0JKT/QG+ASZqnBC3OlX5/eUbpAjTrI80RzWx2wRilSk3BmiuwZxyTFQ
6P2cWaAKet2XqgKjpmlszSi+lLh6kXQW2YA/8Dsom2vkXb6ArVHiSoa9XQ6nSyBJRguXhK7GLlqH
17mc4EJvGIu4AKfiuLm3yT1ZgWNWQfATHd+JbeGLpUm0HidOu2Z+k0O4lKjAExZbioBXh9bygjW5
Vuf3WzxeXP/Rxrmo53WH99Xkvb49CRdAnP6N7o37F+sy98LR88mPdVrZVWGn1qb6rARX84CqmZZm
AHzPdOy2QeRi6UZGOoG+yTQ3863t9pJeIQp6O4vQYXZc7DBQ9hRVgIK7R2wda1r6AkeU4hB/q+Z4
KkUziIDP7ZEmyhqZlXiUrjPJGmQrqooWmUmnr1fLs/jY31UyYvWWuJK9XpkkTMAQyKMpqQqX7bkT
HGVWdNhJ11QOYb01PU1qIrExMydWWD97jQFN8V7LiKQ6h7die8nlk+NGRBm3ak6QePKvEqTve5N/
bDE93Ge7okPboyxKVIRtHu6cbwxx3mlg93e+zOsnWU1MCe9BCZ8vVSff7LFtkXrqa6N55QtksfRL
eJlzvFXoXNSJf/turqZYlHy5DO8R0By95rAuXXQ/C42zaQUtR0afthSnOi2tkmGzn4RFi8hpuksG
qke4YAMF5H/jvpxNrAsA0iHIYXpafR3nZ5iEHz8VeT5UPHDqw348JTFV9G2mReSUDn8YTGq+JSc+
EI27IrPg/1UVQTBeCVX6pj08ssgnRC3geuLibJ4AWknhUNVO/BvEwffBJWK4pixeKN64ZnA8SlFr
Bel0x3pMBXz9xO77Pm361+XamCjvMuyS+D50ltchNaMMK/fJAhECr2v2e920bWgdb5JvHJdRD50s
AeOk3pIIIiL5DpXNb/m9zEWds8k7wwyRyxjxXd02dMxm7KwrhJWFGb/uUDvvabCzlngg4LSM9+yT
1N7AGalY1cA5gNMVp9Oo2BLDj5HQFfRMqm6sQz6sQ3ZQuwj2gMncbzPK/bpIVQh4Ie6kdNNdqT03
l4ImfdVcnFwxbfXtmVB8oCcOy/1LxvKHpodNaDqKirTKFCxHYZMqd63nErmC+mgj996x8pvlmPge
3A/Us13T2AvlZxibT3/ppM1bBVngS/ZGhKF6d47+LKA6ZGHjbotS5anz/HS0wjFpFu8k8PAwvZdu
Rg2Nqopt6mtzlcEnzw7fwWms3VLCVfQ1AADRRXTBnzQRoZGc04i/GDNWkOhdywMUBPXA3uruPxWu
2TyfmMkcCzU/r7oPZCSrgacm8fySwb8Z9iSTwQQZMXd0eJhlGC6zkOJNWchkoFJwyzOsLj6SyWxj
peibzQ/lqjmMaKjoqiH5ZPiOhmyClnw8Plz5wHDbxLxJ8Md71nMGipN0ekf/4nEH5/r3dHDqXNLy
iccD7o2jUdSYoacgR4gU1+4cn83tbwVLBbApIM8Mc7y6R+qKXlsSwfPtPT8LFEHBD/QGKpU20zSu
tDo2Jp9vqI882a0BWkeJujxeM4MvrIOxafiNHHqSNdXaXXWWXwNIQm5aFzuHY74lfri3u8AvVapV
O3zELrem5XW8VMINr4brU4J5t7rr0vcdlqKXJsxLSLjLsHs16ALjNQImFjVlyvZBHAO4pi1gnPsQ
S5x5TqmBkMHUKj/qioIIECKPopk2+eDupXyMdXiaIHbS4RFtuWMg3tmyAXyP+ScLRbG71JcnHH/U
8PRQUrJc5mlFKROWUPY+GpPlxYgx+2SGjufdtNkLkrCkBQIVDNEbt39XohknlhIfN51m58ATyPiL
5EchRuw917DxtKpNFx6lDqPwLkM62gQM0LfarLiaitUprsAYfIJ2a17B1CWwmKO6qLOm/uasSRCy
sAv85nEmcbvJXuIwfcvFJDqlMwpWvH+E8oDv8gZpu+e1cFBumtRMHtxJ71OTvWsEjhYONxA3+VBW
g/NcJ6L1VkHAUAW71rz2KV44s0QioeAohvUZNfN6wjgDvhnxMBnDR5KsbW7KbZf7vzZwRsHc6qZo
wydQfsrj5Q7OTU3tDU+OgDh0QISNkclpcag6PGWL+iSyhAEbsRWHVz4npak2c7RWLK3p0BWRii7P
pdBGK4XhPyMMgKSsOhF5oaJ0jO+QSdepSkPKKQdcK+xj2racYNdRanJ52RQZsFOcAvLFEMTEbBu5
vpEgj+beS+zK9dH2enCDnmBKL63RHR8E1K8uSQC3UjkFWbBqusnpb3H1/9JkZeXHXvaNgw7CFLfA
7TreN9TirGODOoY9ArU+5SLAzn4M2vbU1EWExPLrfPNkcTmgbVRxiHvuKfZkckDtupCnSDtmCJ7x
H+AybHXM/55gkE2zmvcKGRidGW/vLjSqbQ88hsMeAoyjjR/ARGpbmdY6s2srJaStZzIJPg6o0gDU
y8yCCS1eqm8m3Ar1qT0j9FtCtJBzTNLw5399Fq6q4QE3iubSlX6JJh+bdzBG5wyscX33/Ov0psus
e5alxp0GGfANr+VLBsnyVS3Vh9wrTri9jbk5OAHOlBFggAQfBwhVL7+wMXDRKWODEvnCf3G/kwm4
XS7fl+IjwAj9aDeUc501iOD+2odfpRGbJIvGiUK9NMShrE52hyj+JjeOmslg/wSsVVUnE5i4nA4u
shuyabCDHCg+LFPpu7zHxgWN8BGtyEHs4V0QmTqdKUzxhJXQc4fmeuxNDueIhmT1R3e2ZDjdil5S
vRL3ulHfBit50PA0LM/QBAH06cZvDW7VI6pXHp4QZ2DaFgJH2flDQJBj+lJY8P+5+p5fADFnT2LS
o+uDr7blH+CPJgTJOVoHL/1J5KpAXT4YF9UIzTUCRzCFsGiRt3CBkF58GSyxh3JrIBtsJRvh87FG
I4gqW2iE1Lj/fr/BTXLvhIIDboIkYawo6X1NU/niqlnZ2QFa7hwJUEva59jKdQZst/uWBO3bdy7N
rbi+/3XVahohWbil99L7MmiwgHELGqgUimmt1lgJoyPJZJMqKfnpZgyzKGizYY/38zxi64StWnPv
rX2HtVsB+v0nJKIo1udrVFzGOhSrpDDfX4RB1lnGKF1Sl9xK1zdwWidlcsznZfNzLcGlfKO7Cpee
uTOQjPgzCG8Qvxl7WDB+Yb0gSIS0wY8VUi8mde3x3I5vBEVfLOlSYHcEdZtQeMR9BiuMCeZc4uuI
EiVIUlYtOHb4lj2qBP3V5jZFU3UAOKsi1BTbTaJ3cO8WReaxYbxOA1b5WUm8usIMx/ZdbD48a5ZB
drdYq7J2ctBK5JvdXCLi9w9Oi/+RAgU6LC6K71eLp2UpOP+7Qc8lHbnOPKmtx1xi5eRe26rRV6Kc
RIo5kQJ36nb0qWkhdlE1hPhWYoJy6y4sXyk9G2xmJUGt2fvt4oXDL7zzyWIukQD7qtBdiIB8Dtls
fAOWAXfTJII2o/9Iwh/qhMb8DkF/1b/CxbSJWPUQrkP1aS2f3u1qDWgyTjR1WVv1hlVonYVeERgZ
KQiPi04/NYNVDYoFd3ri9Vvyz0FpLYmYdlIUpNeo6OY+gFoNnBWSD3eFYNqCcSB3xyipG/R+rPrp
QFMylnUw4IaaTV2U54Myi0hE1coJwa9p3S2VCUYfNd6zsWVJO9a7Wsb6qV91HMghxx5PBcrECAdt
+l/jYNszLGfNjlM6N7ao2gRzTzg9UTNf3vHCIEg4VkQXuEWa/RImVYN08Cr1VVy29ig4tcbx8brZ
wV/+WvYhY2x90vyZ94o9jVxVlYhiIli8sC6ieTJQ+BnmpWord9+jEa+WHQVOTK5iXwye6YJE8vnD
DnF35773otAULx107bKtL/hid6yI1V/nzn4a5sAvH5tb8AOmdApnBQ42gDIMRjU6IvOzX7pGeBs0
p6xL1cn7SxT0OlwKLH39RIMLprTIR0RS6jEII8E7BVzaeTsScqvW+CY1gqep/34I9vtfW74viyU9
mulX8HRzrj5ipf++kp+ED1D879P0dD8jCvGFHZZfR+vTl4hOIp32FQOOPVAF/oLXfpwLaOJyQWXC
NkXB20NMGpE1pxWAaAqyOHUyb2s1BvDv6YCVTmfM/75ODSLWD1kSfOBLT0jw1HiGyTd1h3jplDyp
XJh7FlzZZD1j5CVasluWEzv5lVAUxsqvk1V2kw2GhJKMli5X6k0UQx9pLcU1uJX790algQFaGoZU
wXU3fg1y8Dr2O3bvkqt6drCrJ+YcwHJZC0P5KcvXRxetHwEusrvEfuWxFNn0/4FSzLDrw359GKdn
8FSbgYtBPryrr02Jds8uM6qhHvpDXY3bCIuPL0tsVNuZGYMunp0p7CwHCZf2YSo283kA3RLpkL9l
geS0Ux7+LwKNn1jY5RRwvyydvVCh0CKllZiawc28zW9mg66ARGN6DyleHvvhMDDzKGxVfd491Wq+
/SoegqinnIDXE11LUI4rEr46FoFp37YJPwpWlNLwkjJNmkQCq/0MlHbu0ItjSOGzenOBtRAkJd9V
LvszhNAxzohTvDpjX7VlyOfSViS3PMyeS6zkpgXUlDutMAMSP5fBBTMixpZiYqBjiRrinutdxCZ7
nDsaLflJKKV7LlcTMlFDjVzsy5C83+d4ig/kXLyWfUlXGTYFhHin/5X5zR2Nrgyct5LV5o3VT8Qy
Xw2yKR/n6Oqn0k6YjvXNTWBHHidlJuGOPRqujrWCmUEezskOmZ6NxvHbaDUCOT9GbxXNRdO5h+6Q
c+Vi8I33lJ+JUO19HYX5rn1lbeo85hPe84/1vXcGVIRdHCaiFgn6ql5bWLbGAUhfiQ4EwAn3cWJz
Pq086kY93NGOWoXk/7c2arriqgYu2lhxgAvhbOJt7CjvBl/S/mb2n6CMskPaz28vTGUnX0M/Z/nc
3wpn9KWKn0Zn19/+TPzT+preErZHS9id4zQa+xV5RUdHKbuEGUqr6lkmbUOkzJ0TThV2zBFUvq3T
2I+PNbppLzhGNXALxet66J38QnWJJQzILXRt74uPrg3CdGZ85fRBe1RQiXY+EeJS4dsPLlC6mpfe
+7oH+7n/KYstsD+3Otm1pgVfMQE9/5buQkD7bFCq+D4eo5OJcXDj3YxVPrqluPIM0DT5kW2+bFb8
MSWN2XFuMjaR0s9sZRXZM27XricDII0ywlORUct+4IQUaUA1SedkfwTKqoNHhmOFsO/bYIKk/xOC
qK8k0Bx4+XiR8P60SYJICrTDwxFEz97mBKbZlrJIbbKfZ2WXbq2LduWDq/ZOBwg5swIzEuJaDe5E
UgMdwqCDiKUufmRneLchbIuJfxJ+X+spxeAZvviIoFkWx1iAMgZhmKmuKAIaNkXJHo8VCviaUhHu
cgkgkRoZUfvzACazCSU/7ctGxm4FZeP4PnIeDACP6fRSS8TV72ehXG8jGuK7M4AgpZiVzs91mU7K
Bghtn+xNPeRjEjpABd1SazCVs3CYoKU9kXuHEgVCtR0Erhfhx4aoeFIwSRwbi0jDbEcSBk3LusPg
t9N3Awep4+FaBsRjWp+hZxpt54TE+zXkIZ1fEeVvSu0DgM4NUcYo6oW9SA49E96FK3ZZmfnpJZBz
f5wzbUsHHUqEtSCd4sbfR7JkdWw4hQeKDVAT31zby/yzfU31TIcZxF3wZrkxZAyHGx0DdRs4RYTp
J9BcR1+2xLyoFoqvR6shOMvfQ9gxdS9xyHeAzTeMCDmvJLHIXf/+O8AtUSB4vJsiN/442uDuf52Z
AV9UUxtlwRjv2xYWh0OiMYFoE40ufJoHm74NDkXppvnFMjDftPs6FhZM4mVb9e7COfEssmW1mNyB
Z+ca6fgTKKAzkdjOILgLX2ZMY9TN9SnXdnkC6bmUZmzoP6DYfGYRjJqKMxaS7g2iZmUSIt5Hloyj
aOXPOOdbT4eQgXw6IPwA8aPte8W+cSDz3bHBNuRPJ6Rjtz64us66ZxlDwFaXtkGqt4nI0oPWiOBQ
f/pqWDCwIRno2cc2XYEIateX0GAVIN2kxUQSYuIpVQsGK/EVG6Pf0kGhk805CiO6hfOJaYgVTxCR
A1sBpSZX7Bm/oRX98uIZq4AfP9LXJg5MsK5fdIwFi/3TEJCMYsmu2J9vbqUxWCI4fxBty6fuaHl9
sqndVF3Egi/dIze/BUK6gCLJFnmqoo6ucRTYujCTtLUsfLHnMP1WTVmtHHW0lUkS5T6Gi1jOzWiQ
HD1jULz81nYrVHdRCx5hSym95goHikM+hiQytR8I0EW/6fyROJa6oKQOR5PDUGTVoLmzMloN4984
5m/SAg8inkj1RgND9NP/ebXYJiwxJzhmO1EH6113QU5gcZfHt1ve2HGLbxwCUvAPX68qZaZqZXKM
DcRKlzrxF4aJZGPcoNLXGwtSsoYKt8B9tS0laxpTt+cl0GwxYrDaI1l89TtGHBXj4bPC/PT6scIV
8lMAei9tMlhMV4eaD1W7Pc/JP1oNgXJ+kQXjVUr75nFBttMP8ShOPaboTHZnEuP6oeCpKWRBG5k0
yYDTKPJyqd5ScZYzGlGw6ppCbqNCIKZgRaLvUvBICzpVRmm0GzP6fReKQKbjb4x4PZKfnungFIfD
6tydveacMomSmpSvpri69Uj+OT50DScE0wDMrv09R5/slHqBj2Mdn1i9JEbDTDS3DyVBAtNkEm1H
FDNclrge1WF9NmxG73+g91QU/DBcNoVbIx9vS77VBQjIeBzmqHNL30TC0I9+D6DbTZWFH2IUYgM7
HExuZVxPpsgfh3YYclnK2kgYZ8dBaNRkPIfktl3hqW3EbzW2rWQeiioGfTvT7pjhfJXmhpMEv87i
oyikA1g3Jkt8oIi10BKHuR7IIaPNrG5bmOxmJlHII5MPyu56tdYNhK9hJb0Nu+jBbmvt7TBJhZ+U
Y/sqOR7y3NNJbmaLm5e1z8o3qsQed8Kf2llXeZHr3649ShfdglbjEBGGn1YnSjEBHQ2AgmWNPe3E
mkr51yDnP3SbvN+xQqCIih30tfXkNhQORPJpPPuc8d0xh0ngRBWrgpaxVRvTm+4DCogNSc1URq8y
34QYWoSGmKJMBIhrpkHJ6xPz6Ponkpbm1LTuFtDSAKB31KfcDkwJh1YBebW/bCPiy7Ayg+VAy8cd
BjCvR94SjgUT200g2WBwsFvbg/xP2EddSpM7IfJcO5dr3OqZj1yF9EhP5f+pgqyUGmOmnlZpfPgH
neu7RcLXzg4DqedK6lNBREmHrpGfJezEimmOsk5//6X/hz+e14Wg6XEchjEJYALUQOlWDEm9fpln
ioI8P7gXEi4j1i0x4cETwgZzAj+NTamLrquns/FbCTYymGB3Vkb3dEUxHs1VfnZphl+/C6U98YBP
h6OiqPp3QlFoIXeZ1DwK8Ya1mYg1RUvRFMZ8+abVy6hleSrXRob723gzmDvsF/DhR8vvK4WTXAFD
wpf1FFZ74wChRP2M9GRqlcYd1IvL47VCuW9v8BEDfBMKQ4/O0UDOd8Pv9wSivuDqJUCOIGQake1H
KbfWYOm1PhUmtt5rF0lJjhJry2DnfFflt2yqqvxks/Z2dPdiaMGPn1xPIZpCgnts+z/yIbRM81NR
1J0J21w4yOXW4klPK5ViLgd+Oh63/jnRuqC7u2met45xSQGMdDwRHbMFPChvIZSTcz+xoJ4ZLq3m
gjJqrgL+0egK10qCjB4uKVwQw49GkPYxG/jI7FONbhoxFHPUSa8/edrVyF0ytj3rgm7VuF/HGq1z
yn5BIbnzK6Oyj7BN3ZDpdVxf0e3jJCAl/cnvhJNWygNyrd/QhL5RCLPIhsF4T0sAPPD++JO5VBEM
/Xy8CODvC+4XvG6CVViwwrJQCXDfnfSKWHTmxOoAb5m/5wbUCAypTQF2XvCJoPA+jALfNweZ1yXW
gRK+D5ghOyYoYWvymCx5UW18Lopa3axnFSjBjQNARZ0CHmCx35NqP7sh5vZBuVuxg9NG1w5m9s3k
dgomEZTYC0laghYUb8FfcH9GdKPg40KaUnvBSZtZj1SpJkFgqEFB/EDlAde6FtljGWyONOiCErro
0THFz0uteShqZM5bNJ7hlw8E7Z/vB1py7qoabnNcHLEWn8AmSKkHDd1G5rIC9SDMaOjQ8kn8GMFo
8vsSkd1GdUJPfI1B10KR/IIVZq+YvalVea39mdAlkxGmXwUB6v7hWqRRQIobQSXEtFIrWw65gT1a
txX+6spYx5XjsWNmYXXKkkqljW621VdCmSBNT835qGm+DShwIxw22cA56uwxCaDcxGeZVwJ5xWPd
3OQOXvmgBAq0gEdQty3MN43dQArNTJrAfeHVDmuuLwRoTKX1aIS45ReIHtTVMnSYNYWFFb6xthKe
zY5usdYkjpMiUS8QsWBGx4+y+BdYkKXpCOWu4ZPUk4+xy9M59KiU5WIMVdc+VmjDADmAajzOryqy
Na8+L6th8V8Atie/GMlOV/Dm0JG6jUdU8ZpC7d894xM4awdZrDQFyhvukmFNy0DOeyPD8/LcrrRp
zhp0ldHv03g1nHUQFTIbs49qVWKlXd+iEKsesuZwpZYW0Ro3q7bBV1XHmO9Z2+bZQT9sQI7GzqQs
F+4zpiAvYPx0QbedE9La1jEIU/1cbjIJdp6TLP4juSMskeKqLupX8nw90EMdT5zY94m5aQcqvG/l
GgBDclHJzGjO3wvUaO1w1HHcWpGOjJtWGkH2OQ2UU7HKL2W5dvsoy29leXiwSs8lZ/3BuXIzeD6z
cgCQcY8qXD9n06FvrQC9OCImwZFKUMvhAdRdYybGbFzIW02G/M9KdaaGC7tJPryKnbq0W0VzBb40
C7AajhEHzawJh/TzjIIg7jKulv2ifzILZ+uZZ+rwHgy8k49oHx6a9m0zkWAmYHVupsJl2pqjWGkr
iIyau1h1y4WcIWak1Bm/AUs/Xzn890WXUTAhKpdlBPSdBPDVFGUOxNJRTTOuSCpP3uxx9ix9j3vZ
y0ZkbnDmudHuREXqQjwiyXjkSa/3wkujdvYI47hoIbXKGXhp/A6PcF9lVEN/wBdToqqDytz3JrpK
9lY821vnBiUAxa/SaUpD9kJ0MXOAnd6e4ed6pOVaI4tPZDVjqGi5sn0wX+tA+AF2CuZs9En/Ou6H
BaQOvjVzloP69MdwPFm0Na/I1Jt1WK7wlaq4BQY9vGrbV42xhiCYFSVhNY+Dqelu7HHkFckzV1MY
JcbboYWjrqT0GcsTRrboABqyNKrWicObUVERZxCxr/osmGNuuuTaSAvFh8U6oR5P4zxuVSRG7rMJ
x9v42lS52KH9u9YV8CsiagdkKOiv1Swpuyv98FXlAVrzLlGuPQFYLmChcx2xGs+rYcDian3ZDhJ7
LvcicBY7cizrLnXdBA/fkFH/wA/K3c8rEJwmc6aL08lwXCvNq9Z0IY28ZzVquUODons1BSVo05Sk
iUGQ6LEEZ7/tMpDJZ2ryY2W+DeMYZI/Ge0hbEMhTrB2pMLjTYmK5TCcQzEHYyvDTdwo9efEN1Bk6
/JsCT7ztkg0MqLZHrxsutBhEfuqpF+h3zlqiPMy8bOnLwogaK1oWNbZGNRTCMwCzAFUUwC/qGwzH
iZ85onGL6aI8prK9P+0KP8/dtAN8CZLBzGtldkrYJB1GnmWP5+mOAR8bf5StXoO3mpRxeCQ9cCKR
XZdxmFh/S3tFkqVLDXmD/KVZq/0vq0nYaRzS2G+sEmUibmFeclEcjgrXDLnFUwEJMxilBaTzSmD7
fGvo3f0mTTf3YsyhUE/pxo9D0QlXQp6KgwAeMHyxraLOa4kfU2gsPt1opfRt3A+0pZMVXNyCIw1M
OSp1Va/AX9dSQkeKOuHDvne1iUShiNaGZP4XvzIQXT9R46mku81o0YWNZRo3irMofz+n7IyYhY60
bOYRX4FNR32qeco9yvl3NtzVc0R0cYLV02fvISLjcG775ALgROqnoUPEhAdxpO3xlMOmr0C2yZ4O
LVR3Edjt2lpoqFu8glrbhqIRMMC5UfvEA/fRZozGWGDRRrLUCDAA2h7GKjbjLOyVKZYV54+Ykcv9
27zGAcEdLp8kbaIUcc43Q+7uZZeu0DqZGsEyYqMIFaxWEN6IIsjwNUYknJhzRc5PwWEagZPXm4yk
U0Ec43dEx0wosjqtaIWuGmzTVmaOI0qMxMPpgk7NP4lrn0QXcZFoa7DkQQyHhgpLv4s6lsAYE8D+
HTdjRugi4xm31S19gepUgLqNl3HzlRtjT6pIme5dTLEAUY+cv9B5lEIyCr6zyvjarZvqEI+2/t2P
85MQOkJMwJRjptfnocckCKRUmCdG0fs9/fnTM6Yo4oPwhyQ7WSWVYX/8oIR6hHNETb6gxK4ytV+a
YmYSC4FGX8iIeAoHvLXzk7lNZY6BvJdJicgnYtepzfd9Z6mfaL8wvWENwG9ZPQu/Sq/fSMtNYzwR
IxG/xTIdbza7ILbhRttpo5xsYGufz82hRwgetPq2UFyMf6OYxNSKWT0Kgs+1ydcQWxtV295ydUnA
dd34vkozUTUFTr51Ms4CGAM+I7VEgmGJnBkhBlxLkrUZCBeIK0Rl3IpiHQX1Ct8dD51vGO0WCtyJ
M+A3qLYzb2OXxDcZ/lzS8sEivip8WHuFu1vojDrKG9Brr1vIdgRWgQIsbTZJCcItb6i+G/BAZZJn
C0MBVrcbS223tUshvi25BuO2ljA0YrgByLR3vu5pibSacj1xIq0d5TbkOF/TU0kRNPsPSGBnLGdY
nanFTPWDmir4efXWMDKCvQzOqJTrVVeUg6zNKVormwxcuuoM+gAH/+T2C3DVZpsoX+v839XzptHs
jqa81mS1FCbI8PLbEYXSBC+2QlhRWeLXj45+zAoHtL7l+9w0d7BtDYIXbu1phr4C+piv1S1AEOLW
Gu5H8pSBPoj2C/Rq4xch3aKaEO/ugYRKUhiM9kLELRUYqncBP8kubxaNFdMbOs5MhLwfofps5zm/
TmLkoyPJWUu6WkoMUwRB+Y3lvdjsUe1G8gbK6FfRFFwbcaizSJRH61jrGmGRCaJmBVHdOJlEyAaa
xTdnIKxx7g2E9hQWuQFZ6oruuu2H0qLdhABaj5UdTn4ojzHzLQT41Un5WPBqmJbwtzV3aAlqVJ3j
yv0dADIGDptK0QU5/igF8bGd1ey3g50xiI479UszbGaksaPce8bRN3piqEltcasX2X9b1hEvSHGY
dxCrRETcrTJxkPhO5CtEJeVQH92+sQYWj+Fr9jq8qQXSbn0lV3cxRILDkXfCD4Z7hLIEVVrScrBE
fzncgbB5XZUIGRUa8Y11KnEYAR7rOvIYZdcf+6eUdcpNyU8vej4fsLNb1M2zZwC87lY5ImkYrcPA
0iRcyeG+/QPJh7t5XZH7nWCST9H+b8BcwcvCUBui1Y2Lu0Ae0v6R2pL8ZMViRt/d0TJwfrglFFX7
4epZc1aIXDbggrlRHUY0HUu82x00EHNcJEdq3RwqeqOz4ipdkiSjNw4Fbh4PRUe+1DrLePZXYNpZ
qc58G+ic013yzljbPhoMPaUMiUu4gQFhKyuogSbN4fFvHz4Axm5/HQCXIjOIPt1wDODMfp3dChbY
9v8TqW6eHN2SHI3KH4W6I44zbuLqeO9DnWliEwKPBoTsk7TxAw+mxYagodGAPzSwSneGh+T5HpTs
V4LujNZ0QRUvKEJHYtbzw3nHEizmTQ9e/rACmUNa3DAAJa4W2CgDyehWcQnyIBIE1Zk2vH+c3NuN
9BzNsiX6jG+GctXzUBdroREfJ9grmmRXk05TjeKXHAj2frp/oCW6+vTYVAl+tdKb6mhbsSAKcrW+
F+DvsgW4JAwhZutigNZpDnmkLIHf5Dsv4KeX8qBGhTVItvP3+eBjSkG4Hi24v5ligWAoHKbzi5it
5Ch5lNmC/OdeWApLaAiIIKs86kUyE5v0+lSytUVo0I4FdqjHCD+rAP83S4tL0X1JI7VnUNEPbj2r
yazJxJoZs62pm1iVSh2LxDyMnZWMF6INgGbPgN96sCJ5HYDug/ZpV14xa42KnhOMV5L1QJDgB8ID
5zBIrfEAiWYHONZcRcBepb5Cej1B09aHThSdfngphIiSqrZp/unerMPpkvE+z6RD2VbverDeXlWc
AAuQxFCef/4n7ESbK7YZa7Rucrzae1wFamwHn3EryHNnKQ28uquzTj9JJlcKqkPCQJpBthfXjq2m
7Ln6sZxpBS4u9DiXsVe7h4fD904VStaI+1jlFCZ9hYs2Fvcqc59ygm3QbnDtmpylEWC4rmtVe4dC
96H0RhEpbfzDZot5dEvgH2FfpTtwunX+uQoxaZWzMw9OKulXD9L77UXK2fn2wVF50u7ZkKovJdFW
IXmLpzP65QiwR5UYGYjmLTB+oxdD8IqG2zIYhjfgUs6uWM9n8FPGX7YI3S97I25VGIEKADfa9oU/
v6a4YwCr9Jx88DY3uYFSUXi7bfqpKwGOrse63YV//xCwkcg87d36pHc2NvhH8b2OKrbgf2R1GnQd
4NYoEloaoP3UAbSTK5Ts/8gmvf0kEzE01BXPZQisQlQejwp5jCr0syq3w6Xiz3RD1ZuJ4Yf62rrj
k/6hfvG4lMz02HDt5hOKZee+f9kskmnYp5ZVkq110vdJ2buJ34H48bztGmgO8ATgcuAZgFOSCneG
56yVJ0DE80LYNsXTPD4qMRs6NnX5AkbMDqNW726+M5ifKCesb7oFjyVn6ZxwAm6mXY9TlNM719UB
3nSSLSK1YDbBuBAX8kNCDpGSwNGYn9P1PD4C5S0kaxzb1oE/jbtHXSF+oAxGp9lPUw/wAS9Hk0HR
xCBc4XZAFB8jzH4VsRNSbIET+7c+4GNbA5xgEjzCdsX+JKXhz6TPIJ8RtEIdid7iE7au5JONHRmq
YiRN36LTXSGXuQkJBjhi4uiKSbj0KS1cQdvOLXf3M4suizVGxtpjWVlCK9PwziWUWCdYbYgSxAQr
aolgAZN35Shk5uGT6XyCEBoRWhavX32DXoIjSgZo9I8T1QhQeB7frNK2m38SkY2pdOc9SRQInnbY
ctM1MvISEA0+vY1dHOHzwbk3zLcjvdFdtpO3YtbFNJ6/g22c3jPZWyq6UHNqfY+ro4pzgLnmfOG3
dONXelbnaYLDFvp/iOQwujsHPibCwb2pM6c6JBQnOAffIxwf6hjA8Ny3p0c1LoVzNpE+0TSqyw7J
+ICaf4PfG+fENLneC+RwDRBX2bf0qFdB0zbVNnlZwkCz1jUP5i1SVzKEs+3sRSiVVLlZXhSmuF1V
nJuY0Yao0H1fvI/pFWxp5YuT+bIA8clvYV4hJYHguI90W5/sEk3mNfVQ4nl/5/AW2o2ths6Y1gxp
sb0WjQiJmGJuPZmW6Ov8d/dcZo6qAM/eU7mQ+StqEj/lDPsS6alQjD2WdHTE8mN87W/T24mOWu70
HJStRxUE0tcLBeoAZiRfr6orP4MF0LRVg9OeNlmMpTop6XH3kyeh8lZrJ8+xDRwfQyvnteUJIjoT
ilYvOmTUa/o90o7PQ8gp4OYePUPI7XuzISvirD2LAg76zqGs/p6vax1BYc6z7y+2nv86lmKrfiOS
eSu2gRD0+ZE7+4Z41pvKk7WY1DSciEGejpCNPlbvjbb7fqm7lcsAyzx3oZb3aNm/rLt8whSO0xfP
YNo2QI759oqnGDMHI9F4QZ8IFJMVTtpxOes1ko3wdJS5vEzyBaBdJnJZUfa2vPj+nM8MWJdRwM+Z
E0CAyremfGqM8q3w/SpqATkIfZCG9xpvbFTsjCt/1f952bWKEE8KH6YuLy8MxRHPCrizcmbPwsvc
bmEG26DXj23x6HG/OCqgK8BCl7s+c6hLYyVjbq3Z8VS4gePB4iH6BRi2mJbigszSdWlFu4tbKaLQ
+GtzrJEnbkDowxNF2tKJoQ3Bs/Zy7kvMFstjthQ4oSaJ6Yi9ZtXPEKNC9vFYK3meExWTs2unAWyV
j6ldW0z/Eqyfy+BJxBeX8EiER4xDiwAk2YU20lDCXjJ9l/ztZz0BWnSeAAPSHjJJZGFmnkX9jlVP
XygS8TnqLuy0rIdrb3MhHrmEQe7ul3DNvafQrsQ6Oier9Ft00TlooEvSK4YWYSg7XZI7f11hcxDO
yh3aKYVAaudrGeObO2/ChMsuEYrQmMM9GaoSUHlui8HZ9Q8O0x8JOQHjSgWTdtZatFPG4dkVQChf
p2bo/Ux+Lc2SZpQ4jA9RDt8cT1iN3OhtvvNGF1vmakLAa7Sb96504t+QqstXFNqF6SzljV051sJO
48eYKRrwZwdHEjMyqi2gtY90jXjblYMfmjSmPxOhJaWZtOua2xIoS5kzrrHvlp3dHFykv9n2S/u5
WtW9scSARmMYIyIIkBTea0PW5f8wsQG3gd+bVnc7eF5Bf6ag6P3nPWBSgkSDeCWTSCfWdFzJxYxU
dfM57IWxTTSOsXUAmjiD4vif23Kccp+8ajWE/BjT4v4RTQ7KYfz3SBvwEXnIrk/JLTKaDaEFhJcx
Fh0euN2nhPUQmSXDtlHsXZchl8sEFCYfvEdBWqr4d0z8IBy59mjcZvujEtg6D071JcPAEckelpus
GgtIKsbospBQMFQL5wsRbKjQdIbiolcgp3UKVSm453TWi4Eye0OdyGv+MYNsz0tuKhTWISSf8SKD
8mtCV54BZECgDXgs7ck3UlPHNk0VDcMCI8bUgtayX6kr6avnFLZlELGMDnM/bfISC8EdZseNB4h/
ykXx7WQcgIekrbExrvyHbScq5MtnluGceIl0Ot/N31hdMgks4TdYEnkPECu2liZkQ0P1/rlHZTNt
oYPeGnVWlCUGxxu2Fi/1Zyse2B7MIm9HzEsztxLLUYg4Lc23QoO+aJLQV0bVZs9LMcJQQ7ZGUJHy
uz1KMvWkNjz+hxHYlyDe35KMsDlDLi2LNsyI72IY9BLqRwNcBPw+KCzSZbwb7etSKoogAQiJ7TMJ
nXKrNSYioCaye8QI16T/8sKlgWB+T/Qpw/uJ6OZ/ro39Z+MKSVEoHurI3yBoDEhQmLDQdFxuc06X
iRyOPhK1/1mu6W5Azgjoc+qhu4WxS7T+0zYRNPHzJRdAAsUbF+oSBYiClktxG/JcW+e+8kRkUBug
bGBzy372bMymYTX6w9+J5pthm8DqG1ACffRRzKNjuNE6lllTUtUOY0fbbFjq6X77Ap24wLw2OO6H
wfVKdL23tcMtIy9YjSgz8Dmd0jbbJDCMJSUB13FCJo5uuk8M/qD8oxTUUiVmECrY7BIrBNBlUFIE
yrzBO/cCVfQTEAMg+jUPcoy4UuEN2hMhj8XopyzQtJ11FTvjHCExgeJ7vZCeoozlnqQrkboI+vj5
npbIdC+pNLsNaaWHI1BDwk/3WCinVbk+Ry8rq58EqDhdJI3FSM4sTl7C7gm5hP3hUZSTcy9ZxqNG
EpG05k1iIeuijQt3ZIX4rrf9Vzj0dB7pXkQzv6kpSJjCNNwK2Ku3g8E/nq9hagrtWJy4PMcrq9/M
K26TkcFO/8XTGavst/uZo+CKixh0hxA9/SJw5535m4RpQiPeDDab+/5+5qDSwy2MUFIiLG63GC4U
WD3QKbhTZ5OOfN5Cdmm3I00OlRdnATqCRVwQdk18eAWwWWx3WcmfuF2iOLn3U+GEsKKStVy/UXql
yqz8DYZKaZbvGnpzWky7ZkDnzt5qVxywJen8vlFOc+xB9Zh36/Z/bG2fUG5jScqieMSkD+xkYVF9
cPc8LJsEptdor7i5uD2sSeOhbSniarjCeSXK+Ytq5znrZFQNC33var/jM+lk2xHvL08JBUoOXJ/0
r5lSBOLrGI9Sa5iW6a3vKIyrcffiLO9yAbCWlSVyOhD+QtYB5w3XfIb7LqQmwdxsoTdmgbl3/MUQ
NPUg97Lb5MMjuZYf09PL0Y++TRW8Al6NdGBNB40AsSrvgRCnrl/plxHPHrqofx+7V4wIUSLb4C2b
Jj5Sp8spi5atbqS8+Cw2FRoiK/raDlgrhQecU/LIVNRqWPBIvEaluuqk587EuzfGWpgXQiNzNBTf
AayXnpxwLNd6cl66o0WoplBJnFKPdFiDx3jPN9SDAgcU1xElX6Xzamm9RP+q/msnrYJpjAeO/vkt
5jZjA2DNbcUDb4B2kWiimLzMKc4eAj6eE/u1RZwyBEUsGb1ausJdqOFkz/V/6g8WBpkp9XHDj0AF
SyKwiU3CWTXVp4ejotYwSrnMNyyiTiNHuKZyR7zNJLpJ0GPFAkVddc74lmI4P+eDWgSc64hIQRQW
R1ut1Eol6dduIxRoQ0x7YpEcaX17AFBCWNhHNN9+Qjaq1VOzD42W+XnPVBNzFXTKXzFcIDPZdGrF
HPvjCA27BZgmb3lj2scZk1eQ1gyjmhnRa2H8VG8X3ieZtqZWRmfW9wupaM5kcoNaD1ijA8+DGYfp
vwRm+QBetoS70Jt3KIP67Vjhqa1Mx3onKq6pJMANq4Zw4U3jbbcoQt23D1p3qNe8jFFmf4YrqI4Y
eJb4gjEy/5dGJ8ANZm6fCRZMdOxiHroHZy1rnTWYCP9mU+TlKmy7/EHy75cdP0wQj3qUIlWfYccl
tE+9D7QJDO+hb5tKx1R4D4jVuK580XuLNw6P9CJAJ28M7Q18zGuPjx/KqF97Pt6Xhlq0zh4TfVLD
nSCPMSF8sFUbZHtynyUSl1cNUPXldMAOZNmi2+wtj5XBnLjkrxOaO9OrVIxJ77avePa4qUrrnmUo
YITw9CeZ7l6IJRwAXcMaV5BzHNzQUMu7vsA9RrrK5YrOuuOUcceNnXd3A/ZdCmuhF+64mAYJAiHj
l/ZWYPiGSkBb33xMhvRZQjmEGIdTiL8rOt1J9FEEQ9pHEneC6SS9B36bUA+2Nn9LLG0Epy/kuLhL
hoN0CcClb9OfhsfYYGFj5Hg/XZ6W3qN/qqCZGZy15Q6qGWTjZuP2c8wWZnr+BiNnryCWuDHgOCHv
2Ciy0spWmXnVvwSRK4tJ8BiXRW2C/QEGQLtm7NCmJ8rwlm6F6lmo0pDQ3ZyIskEJED/d7VmM5WuU
2wQtpv93O66xnmEBv379qiGfjf7nn1+u8LfLjT9CIhnC3EcTvva/tgN1qLGGTIcbv5cLIHd77P4F
jy+JtCbv9czu5bOqsALQk1FypBMIxcS9v9oEXnKx56IQH/GrOiJ5dvb830NZIE2yvgp3EXX1jUAI
hCU6h3m9fQFYkF0fOAcDNsiowzCqpXoKIQr7mQIf2DEKIqaxuWz07u8tkiHMFHUIrcXJMydIP9sx
Zp/Xa+u31pytag2+iBU/bVh02Y47D3wEclK+vXCzOouDQfBG/V6lVgFU6WLPF+uE02g/JVi2LrIW
cGglax9bAX3+tOgCfJuwdNLICJPvQj+j8adDfayhF9JHaNVP954wnSydubm2DHr4sEnWDCjRrncn
5RJBaoFGYgPy90MwNYutz7sPIBOpUYjJPAHUWPmxY6IgIYoQodVOZwt8vzNttwseHR6qo1wdhcYt
4rz+Jrc1EQyEK2obnIGq3fbxS5vMKSVAxWNCfeaswUkRw04LyONdWLPrqiXgkZXpnxbAcpq+ZKu4
8Cs2SUPQSdoel1f3EPI43RP82AKvESDJE8pQu8kdXE7Sv7r6Wl/LBVQQ55zT7coOcfTZJfehuz+o
gnsVxzIG9pEgQ+U9GcY+PdjxO6hD6AkaCwIxBuX9rmPOZrgDDO5Zeamop6XqfD3M/yW648ryhh86
iV7LTKJgw6Dl7gaRQR1Uj4Zl/5munGSmvBf0CJpSezd5KXiBG8h3J+qM/4/55ixhKDHXTp0i69/B
QdDMUQ+QxDCmz/GwiFqqEFIPBUjpgdVRyL5SZ3M9WawpowQr34dlXmkLlsEb0KYtCEl4Wsq3N7iM
zwDN84Roumsk5S/0Gu/Q+Ulqc3SN+YqzmJI2O6iJmL2PRkPK2QhTtU1iA724ex81csv+lVORUbbX
KHOgEQ1Me9hmLgCmAG4oyjq/ori5OGDoxjm5b+1S/UOy8xVv/Xm7z+nO7oRJZkYjdGUAXtN/3xs9
oGKgLY0Kx+dFwy3NCUWUz3UDpQEAMig4UhxU80tED242S7sY6/l7RI/ilMxYE/qbW0q/rHLs3tk7
+xjV6fuj6cjhFFWq3QIwfe1ZYdA0rSJHDjohMzQXA6VcpVuwwrVqwYo+GuD0tV6ObhcvaOiVEGlw
1qDRFiG/XWO3/FWk+CRRgZk/jyDqlbgQLXAh+ey/gz4izabidvQie1/OjoJoRASGe0m6p7xpmNOx
torsDV3maqUck6d9/PXpk2cO3j1lR46iBmROj1YT0DcsABuhsqz+yly2MsbicPGJNxhBw33d+K9Z
96NZr1v8n0b+j40Cw/3Lc2zAFtYyxZCRkVJEp0sQwiz7tZVO/dHDyWCa+6rnZX6YPMTPmw2WGMyB
+a/S4hd/p8NL6bQmXN8Lv/Nd6vEYpsl2CufjblbnjntMN+bvLd70qkWVaT4EBYtEJBAcygccOUJ9
wEEpNUQWTFMddA6zk+qOGUddENUE2XpBKSF6Y8DKbnjklxQAFU3L5t409FePbxm6a//jyzJ+snLu
h5Pcss10xRNUWPELHsjWJeuL2CGcBkSwcgsqXqbfh0vBkjpxgDJLiitD/bGJkQM2+PdsrJM65TsF
H97/ZujxX//DTIFr1RZevggoKfRXgkvEeN0TCY2B92z5uU7e/lxM5IqUJfyK1BqI7XzQtV+qOraI
8J58UHDa6uujw38XOMRcIT23v2ZC6HUvJ8GwsNP34uDxSiuQJuzxvoWWfHDN8u2RT/5obs1oIEvF
K4nmFLgs/yl5OWO8Zhhh+iWIwAQk+Iv3is76ix1WTMOgO3zm2rRhlnz5pWsXfwk0wkrnjZQJOxjx
vAI9nRT6YMyhCZHnfclOXN7K9afdsy5baI08hNisUpcmYYrar6FQp6KLY4avoGtB+B4qivMpKG4S
bQ7U9qrB/HM76y3ojVW2aERKXrLh0oWcBOfQ0Fkzia6FXgMgZEsRui7Nv/DZxdDg+ZIh1QjooFXd
dUYhnxA2JuC+dTczhCSjIkacJRqtElTVfVy0RT2HDrhUllVtNp0+9lPR/iBNC0v72pQMbeUQTvGZ
zX9UOfrnshoNMAOLyfa25XzgMm27fEyskv1IuUMT0IVZflQ+vKWpjQXbogcYD9xby/HSgLtlYgmS
H3/1BPoMhnjKqfcG6Kp2A/DxB/F+5uFjX1Vi5d3cLgLZjbmcTtoFcWIyo1KUtWt+WR4fRhfAOZ4v
PIebHeD/CtkG0bqXPfi/kLLsb/svzU5x/xPxcP3872izFgTxaR498FHfj6JIa3i22c0hVraFPLOC
0O5eQXKPIEvRagCIElVwRleWAoiw1ZkpC4gL49wmGkrXBjq5tldc8DdhP7pFCe9Pghi+aEOaXj0K
+q3Wd4hlRdcp5hobH1PBqZMiyItJ8OYLW5hJ9LEdYHOMiRuQ01JOS2/TndRiHUykkIO0BkVvvAFc
L11FSHfelAiXADZ8gwaO+WKOzQRIKM2Hd5VRYpQXeZdeLL+L/NN0lCYaS3xR9F4wCxxElfGKbDka
pL4t0ZHjmkggm6CpF1VeQnqboLgCZj1RIvKkVOeIpohej1fiK3ASrBzC3ZobFhw+kLM3QoJVt1ip
gkf1gIGeIJSOlEdYm7ubxghil7xBc4LGA6SkxfLUdQPiimZ1YaYmxd0XwafnJBA/wGycCc3/zKxa
nzu7Dl75h7Yc7Uh680ix7RAk2K8iNocmSkJMNAjshkSl6uPB5wK8WjO+Vkiksc+70YZX4IHzIgJE
xWUaFjv4ifrVm5FzxNU/i0lUidL1i3FlaUP3Vmay50/kkiPhkKu6fNt2DplJDts2U8QgkYyiEsNQ
HxUg4SOlUy3H5vvcRc3HQm6apFUeL9sa7SdH536PucrhRqwp3f8bt5t7bePacs/fX54fRcfp+bdI
+7AI643KDMfcBl6p9l+byV+MZg6xhjbDPE8CrFpTNuyl9Or/t7LGmIrjNiksJSEJd3S/ru8FQK52
OMppNPUA5V2PmBbAOYTXMv3Zs843HWwJaScke6+koO0G0Wtl/R463pfw7oX7+qt452UcyM+j7bXG
5P5+z7VLFpMlWOiYXkrCq5X4y9n6uO5dD+oERGlpA+lnyNQoJhLiHGPa96xUtma1WgyswrlAz51Z
SZ0mmimY6FEQGBs+f1KDYfUd6G00XKMfIfWWK0Xy9UqRUGly/KilWuNIdN3kenxlOOSZFZZqiRSR
QWwrg5OdM8kKgSylePSGE0uFcwZyZIH0ABUcaJH/N3qwZAQL+12S8I98JKiU6cIgaVkMWE6fSMS2
Hw/B+KM1Ur7nVuq6OAYPdy2Jgl1FXm7Cqkg/MlegVgbr2yOc64SYx+27n54mkO/rTO14eiceurrf
VwFvW73o6GY9BlpjWPWjkGj6s/vNHfkeEXsJ3E59fwCKKOnf1SkeNmnQBj56B5wc6CuP0k1c7MPk
ae4KQvzTzO/eHI6Jz1kzQcXdkwzBrs/7T1V4r8rKpdGX+0S6mt+3IxDCfnhWGCVrKCyBZC5CaTU4
l3fo400YYidQlGr+IgP5V2Sb9QhVr8TsuU4jHxPW150qqWLPV9sJDE76eOl8hbg879GUJ9+HvJTK
qoIWdPnGe1ENcB3hepL+6tJOh0Bw6oqZerQfQcB7oF47gmTtX1cduWT2SLVXeDIH9/A/kT7ch5k9
5VHVT/si9cwUUeTGQ3XtbuG8J0eA0mS5UDJcSg1qW24G6oBsA47jVUdlxUgyDv5OzJJ1gEqwLMUT
rh4TXG2tB2s/pHNdRtfTDpACqRmmQxGjs7lIcfAIdtmy2m3Qutbck4KmWMBBgAp2dFto2ANQK+TD
SqsVukEwN2+4U9LZKQeP/MOBHUzFCrRMi2dOVP9P0nKvrMgv6tCWfBOk2MqnIpKM23Qt3ti9QdmU
Pb+t68IcK07Bw4g6TpzYYAU9QTRZdNyNX+JLzG8aOqm1IA/HArAqIkE//2ioadaJJVnmV37Ls76T
o+xvb6QcIgZ6fQwdvaS4GczhsccH0mO3b7ICSNnqSvsDTMS8IqIQSDsJ+eXN3pxZA7CYreOaR6Ti
DBGu6szUfRDUCY/ouO/dyKPOOG4Nm7dBnYSpi7IBTBMkkvDCcWndfpNN9Txq9J2j1I0WjAe6OTv1
TfYi+AY3HDKNRfkdB1zOzJFih5tcXhz4StQqqc7D3D9/5ZlL2bct9XIW/C/NC0D4+D9ZvRFThLsI
yEc+VB0crziwl/nwtFe/zjScjuurAGQQ8HNUJFPp/MJbI7pnPJ9wmmhCSJ1bUp56aDkr/S2eImKc
nPhyBZLDzcVblZuDJlVw0t/imWZwVRSspadiPvjmOS1U5fvdYWAdZy0JsEgKHmSCLhGKDeyEx6qi
iTPq8fEoh5xs92zoHS/1OLmJg54rd2cZ9mal99y38a5NT1ciSSB5mv2BPOirdEsjo/bsuT3mPF4F
nIeUGNq+8lYfGT6sVwnnah6DjLE02SnjHLiFUhc7+NF40MZgG6u+6LYJE/scYk5NlruMEK9PL9jj
Hab+fvdBrMMwzYG2Gdz23dgdO5gbNdNRgHNnN+wFvBe4H4HTXaWpThsqOvapidXCsC4pba5WZDZi
FqIWDxmxg1ugthQc/HLdrDFfT4XLhiCpI6lKo8g7+FR+YGl2UZKRD4HdMV3DPkvT6SepevgXjHT5
Cc9gm8CJiGYhX0RPpmFUv8ZvMPE72R7U3hBXt95pvGCiuqYbt3mc9WOlD3pHeLwu5fgcjNEwZzxB
1VjHKGgXoY383xue5yAJdoyAKBjD3ECkt2o8LqlfJcKKvDrV2UcXcKwxnuocZj2nfIxuiegoNkV1
9EfjovD3yIkmRR6JeRVjufaBtBkcGGNcsJpLWVFrijlBwRxo47uabK7VTyzU7XxUMuZ6Decy6JbJ
b9CIUlI7+Fc6//MqLvwdX/x3FZhuW6Xtr3qVW9mcZxvW5OZI/B6F/GtRccoy6XW+yrGZWqnW7gK9
H85hXyRRdFHS5N8jZCi04w1MPvjjhnenc8y9NKGcv+ualQMyXCn3EFBgdsJNMDPHP9YPMF6gEANa
3dlPolwKDK5oFJJibUCgLXf+kY33/cqAhJhjpC0mO6jTIgy31+TsEkX5BXt2vYJD9OrAKDjrE6Yk
17OGdMjyOUh71D+o3DSRnZiY4A1r0f70I+nkW2FVPhntPDWoieoRxUjDIEnznBqHomfZUGEKCb0+
4NUSaD4c/+LXqdf8UhzO/2/dy5BaHk54OLFgLlCCBu1UNF5kWM3Ukc9UKF2PmAsx7giU1HhNw+sv
Io1YNL8qetpNHsOZ/GoE2RlJk2pAUn/OjkKMaDGDpKPK82oV7/EbVFVzVxv+V9YBOGwb9P88Z8yG
lkYrUWsMQNH06ngExWQC1m4WPNWON8LZY3+9XqH776IuJKINxCyJKU1cSrGecuOO7tDMVg+2uFT3
SL0R3dAbhQh9VGowhp4WcjkOrS4zYTY5usiwY4FrbbJcAf+sZ6bWLYXxuUMYGs+BmeQ71v/TBxdv
x2z0hQRExbOfEZrC45gkrhlkG/cjAM0RgxTbNkIx6qMvomfLqoro1oDbAUez03Lt/gMzvIPU0aJK
OyUomepoGFpKNtbK6zP4FjQPizK0dFdGGUlUu3WrJ5ikWlmgOb51Pd7TwG9JPmuBSIoqzO3/Pckr
vYtRYTs+9CnUc57FXvfHAHGBDFkMHCHkrT4fXg/tF/0K8rOJnGKFsNh2piXStYJDYWYLh1P8FFgg
ij5nsG+7KjZhcXLHIDQDMtIDsnDlcjJGc/Iu/HXk2oQT77qFRX/Pf19uCmvHEiO8mnHmYGz+BPXh
XaXAEc+I+EX1XEK7MkmMndWMLsygOylDTbyYy7+soR6OWqhytv2w+LFauaeimXHeAzXMk3Z4p9fk
SJ0408m1hvfMlddQlXLi02q1hVkHimdtotB1JQ/RULCSEvjwui7bZEfepZQPsNrRTp9QzWTZSELu
kKOFaG57bn/MruU2k1qNtpZxzvyfuqRsxpI11qa243TuMJ6V350zLsql5MtgbUsf6SSfv4Zs++al
3FT3WKtF3EbKkwOOrECEaEkMpLLikWsVcBNvD5rXT5YH0c2LqHpvKv2PNrqFNjci1EFJXh3hcQw/
t6KrjWwCnnOHy9fHBd1vE7aW/vuNfE3FF+eKt9Rj11VQ6hKLx4KcG1bnZqyXWo0uoAJkuviafSkb
/Od83sPuielp6tJKNFcY6Wi01HGGsu0r02l8HIclQFy0B4COnMJDu4YVnYmktKfLDTfFBRGplkki
AQJIwNdverPFpf2kONmQizFe10XPQ89MdilxGI5xfgnoiz54gWwT4jMq5JW56DehSvaGeUi110wA
friDQapxRlDUXz4DlITJb2DCCubjj8Y4zZPg09JfXoQ1QplSOwWLTfQMNjdPFc/PjACAxkGVQirc
WfpAV/8akBNbdg4BVLuBy0kO/Rzm+yQE5uOGwx6/0yGGgSrvLX08DaTKZKa/gCLL4cFJrPffoB8K
CVTfaJbnO9yfBxAdiQLRzX33XNXc4saKmyJmSq/UgV7Nw4M8ya62fZsyf7up3hFnFkG8Xv1paq4O
g1nB5Uf/jq+8wNpR0+pwxBJPLRUrgYdI04BBJDlSyd9Pv7Lk8dx2VRvvuYc2/zTHQUQC+HVJ8rFL
iLWj7aNmJZgShyf63n695eG84VBcg4gXBubR3RkxFKlVylDuMdavtXr1/Xl5ZTEcH1dDvJROlPzx
9SUOo3s7c1c52KQ4iBaU6XhNc6GChzn2mCmrkEpYhsu+gNrrlE6xuExWdqFNQA12GLz9E3R6zbj7
MsOCZtrPPqAzM//D/BNeDKXeYOEFs2UITGkoevzmN+quAGJ7TPRp+JgrrTuETcrLqYWJkb9sAC8P
9x0RRlQSxcgcl9GlaclWZB6RPxNm6/LNzHnrHcmE3XqKiT2tgmFtSYnutKEArmkAXoEUxnFVHq8z
wPVu5ynM5fQnZxGc10b2QNuC5JfrFRSErvx+PCLNsjAAah2VW0HviLibQ2IIfFeLnmbJnc4RfkVx
9oXcHWE71ulZn2qQIyMgNtIoLaV/P8xNYzmsUsYNNfNc1v9daqSZPXv908olkTtzk6Lz9m1MrtxN
XxNM2KNkenUGsWIqM2wZAeMx0Sfqmpx88pra0H9p0NwnKQaTbNNZI4qav5INKtZ/uOiaeecOkDDh
NKLamTDyNHkmr8AIxh5Mf7E5wi05lezhvsjSLR/h6tRXZ/H/Ql2KayGurHUKmpOSsxqGRWUQvyui
Q239kVpDmYyfzkGaTWVAidG6TMnGUB7+VK4bY1koY0lrYYI3mfPuwQgrBXM8pZvwnNuaz1kb2piD
rCGWg/pPdIZ+qRUWLTUbNVbdDuqkSk1wBB2ZurGs/PP8bYw8j3S8blzez2qdnJu0yryuTZ6gHVw7
uyYLegQZv7lSVXfAAbl/e3B49GCl4ey/F6r+arxHlcFNvAP76qDIQLtnZUIkSsJ3kD3SEpNyLniw
iYm/JIHvr4DmjpuXtMWCaUk/aycUeAm2Bckm7oSjI9P6BXQknHhWSSUZd6LL/KxjBCgOeQgFK/K9
jPM+gOaQjWei1ADZ26VLYTFBRxXtwP2+H+RKanxsH/huJgs3M4js6FuJzaYrSOYtLe5XqOCZuhcj
+DjatfMirb1TyEOgURQk2OI8wSQIiD/RSJAQml5/sF8WaLCdXn13NyFAEkda5W/ItSe3jrdU2YLG
khbUMbk2aiUIg4AC3AnuAcqJJ2Lkr1rueB4FKVZEErcWiEIVwGhbHOJIxmfFvkhbqfwm1X5FGRr+
ej1Kk+jSa3Km0gtL8xY8uboLZCVTh8npthDWVKxCMn8vfhcQ1J+PqBvK1y8t7WNuAGK7xszEZma+
xa5KkBT2PeiTOq5hZ34O9Zm8X5F48FJT+KI5r0H865Fz59S/8w9Xm7v0YoCpUI0trFcDXYNP0B9x
CH7qCCM+NYBnVN9sq2+y0J/kJMtmGz8CwO+vvWWutCTcO1RzvCM0sQZ0VQIFgWV6SY0THQuv7gzz
EvUibDlgtnUSBMdUDgyMhjPAinWZvx3hfueMTpPUuQQYak+z4otUHO4I6N/JUAvJIfwtfSauDKSl
VHiSsw6+I3LjuaU9x4pd/3+svZ5BiHVagQCfPa4XIF1M6lDaY8VeEMLZVscxFXC4lUJNCi+bQ4Ui
UsjSKex66ckXKZuxGMTe2jcHDfeFBheyFyaHRXa65Ln8TEdXQ1ShABLuDjmSNlT1RlayPXfXABri
e2pXuCAZW/RpwZ8luaRJxnoDB7SOw2WYbvfJUapT1nx/gAUXG5L1GrkVGb+guiwWDP3DrDJ2mtML
F2ajNzQgoTBpEBl2wENsV/eUMwdHkaOBwwWfQ8/Rct/M9zsVvTkTo5w1YYRnUVc8Ni0IP5hruMMy
ophIardQWnnNWlcfWUqkkKY/4E8i5hF1qRDdE8hgdc6tcXoptUXC0JQW0YVvc0H+Ns2Pxn+KXk4r
uo19soR9rQNkfIog22WUCG9EK7zgQRK2eJwSKCSId3r5UMcK5ud7BuDI1oCstRF7cYXEhfzO1ZAW
xdbWCRIv2S54RSGWw4o/aWVvl7pUlwLyW307Uv62wGQcJkrUP+vjTX6o05SHuVAA21KzNFv5Zu2F
Cuy2zBqPT3tWylJKE+iaVJAGHGhFbKRrgMgYP8fh9rnrOSwSnD+Q54SDxc+nzoafwr2oL8yjls5x
2ArAVKJq+B0GXZlcJUwOiEUs75ysUVVTgZII6z5yGD8nYckDbupmPzNV5S+i3K6FuBC40Lw9UgDb
ZcPLDdkfdgcVop3of++4od3hYowUCJd8ZLNYvfT55fi0+V26RT52a9DciFYRgfh0H0iw3SsEkLpO
0Vkhp4YVHm9WYh4RKjmxHXTukmn6FvMWbs3RexdR86M9IJniOiMx9bj90hhLPSL4Wr/Zp0HZndF9
LrC7SW3u0wTpQ/UC8bquN4/Ne30c/e6Ueddz7n41FHpjvIRy8p5Tp8crnzf3bYKrzMk4Y8GdoBtC
GOmkpEFM2ZKlYyclImVWpXC3EWzPS9w687rfrrpc1BEzZeQC2Adzs8mZ7K7xNvFmU+vXYqNS5TY2
AzwUQwxe5B6xljQIhFOOb5ri7FJMbY3YFUiP7VohshxDoGA+5jjHKJzdsFO04UJHdyQFKN6nhZD4
qaXbn9mKvL0FcNcrQTEvOIxyLnUqDED1gyuhizPOTiU8vx49U1w1Kq9xYO9jfsEOYha2Kzg+Dcoi
rJAbe46sQv4kvqTQ8vzsedkrB1rQgXZWDTdWun2sXXPTCwRUq2S3ovY4q8Ks36HtWO55EDqMe8NF
48yz79XD6ZuzJyxmeoC3w6IZTY217feDiwSZIJpDKFoLxwrdJ99gpNQ1sSMFT0FUk2SiTZKwT404
om13nRn2ZGoz5Mnt3wR6z9wYsnW4Eris0q0PTHCSo/vhUx6Vi36Exy6jFRv1fMc6uHHyvGEAYiqf
IpRqMsYkJ5uNvNKoJrDcG2Tamil0ZOKAAao87yRMBkEzQB9lmzyAYZ3uKLnbtN5cFjassaCF8nQW
QFgoReyURg29gVUI0i6UH7rtA9HEMxUFSci0A/CjZkj5yN9NRq9qOZ+67YBJ47Jd7XIOQlD1nCfL
4aO5heDT0sTzEk28Ad5v7nBI9RrdT+NFjVm9qczihb3SFRlUk6fXOrfNWjOy+taSEpXjP0pXSVWb
PIOZWmAaafLfiTjGh5nCEBPjCQj8EpzJfWly625aUWWAzL8gLN/ZA7vguoZ5ykGeLWY/h+uIA673
wB9N2V91a3l3plf4CK1nuHlg71ziv9crnjSzlMXAsPws60OGE9PXSwjLNUUCYJLpySdirEVn9jmz
PsJlR6dXtUtsdrQqLq3ynSlotFSeBV46mdi8XMHC405I5/QTjBK8v68ExS3DTB6vKxYpo8BoOsuf
TVg1NaM19oCSKwJQe/2yHiiVh7BWOI8TMmeaa8UveloE1kLdsUzzPbkhT+Qf4ZEOI1Rj01gelwkj
j7Cc3SC8qhN0Wr4C9YYUprTj7+xOYO3cjTolYnmsPEvdN3LqkceXNWz7LovbCYgqIVbSNN9QlYBs
gb/I5b3MtzRNW0APZsJ/JamEow/csPfNOh7cAvSej9/lYXgLZstKW3Uw59EfdX3aNLM6Fen42D2q
z8fy5lUkTojaUPkIv7iApAZN26Iq4B/JQ61UiKJLBLa1mZDbzP92IlYFueUhQOWL2lnzt3HG37vS
5CnU9qf2yenMOdgj4hr+Oy9cVGGMTPuF/5uTsO5XfJ9Lk+xwpjWSyASPHb7LpXWCAt43i4QoWl6h
RXUSy/WyglLSEtTVZVZA4aJGDXONbi3R9wKo2eMjIi+dMtevatd1GTYAPNn1IbEHRl3nKWiK29li
hs4jqIIpR3Lfsyu3OKzd7SFVFqKYw/QJQ+fAAtMyFtJLPlfV+rR5I+2AsWgGGX7+ZdxzLpZvwS/z
iVsTVtIqW7fdErEdROwIzJw03JUCprOWLVrQ46wvuUMnbNk/hNgc+oTlYKI+qlf1348vrZ4wu9Xf
v2vMHuN1wNEAyW4KfcZvy0YqQD7oKruagxpL6kf8ie+ZLd81lyb2Jn2gRwnQCbnSGid61aI/e88V
Ka/P0dP7Uz+LP8fhch2fojX4C7MuVd50OaSdMd0PQE5+hW3jAWzxpXXNW2Q9BMk/op27U6ku4re8
77RALmjVaELApRMrl23Tg92NDK5cGEt1Fe2V47GDrD6K9s3oDXxmcv1A+Dm9JGQ7BKyZGgCGvrmU
RrVqCbM/W0rUJFfsSPhHqbLrE/hobSS3CaC4qOPzTzWuMUwgVGv1pZmncaEpLtUsiE/iplD78OHs
GMQZqi0jDx6604GY+85FPmUhfgWmpzDs7UW03oJC0R94/qQG18JPYqLhj4P4/J3Hhaus3gIZmNks
PR20woFmYFZNsyd4bnRRZfKKcbWEg1Clkos0gG0AzCh5HSKhdHhKW4zwGiXnA+Atpjp9Urg/lNlt
WHcvZHssYhFF1S1VaQIqZZzmvha7HaPy6Clva0NSxhcEHEM7o35/u2VsVTRiCETpg/1n8m5jRj1R
3//c8TZuLHYmwTyg8G65+bDB9PMm1yp6x0NMrYYNB/KMWx6b6KaeeNR84e/bXJkDRzMJ+jiu9H8c
yiT+kl8XtfFWtLqGqp0w3uRkYZ/45qtHjGPW1dnZ8lvUm6RoUDq7XAZ1XOOry2XHFGrZ07mO/O5I
0i9UYSoXPI5ZczNbUGaRsz7nQsXXbzF/uyiwYRVrO3Wr+umSIZIPU3rzmTq+MVodb27zu3JILIhj
oE+KegEuMPPmrvD+8xcWZ+o31J0ya8psTJOmm8yIIUKRfOAp79YHkQEh++kVoU6nlzHFSqMce5mZ
uCSoynTNAj9EmwInnTRwJewMkfJljyh6zSfJBPxMHGk33bhryJR/VrioXLkKWf3IDhQJqREnZ7dc
4IuCug6uEv/N6nisLivI+rKywzELejT+8eYgHAt01kJfHeM39Q/Uq8KqpBa+YzvVvcmYZtMzrEdk
tGuo32VlE1B1Fq+O8Jw91yYplQ8VK+tKHQKgZxgvJ6hmVVCg17ekHDnFJ/KUhqZwyQPSzPCLnZ6R
W/9mf9ZNt5nE4L91nPqaFUMBvkJ0cqcOgIlQTjWEIQHrWp6lWofIHAn52LPPm42zcKNe6aEo4XU/
N20CtWbAR9kTvT5PRNt3tP7f6/MDQRbuxGgld3lazWU22SJukjITXCNJfPEniA23PMbzKykS1BH5
DD16/1S9FGkNGqmpae7kOWqrYKQuST9N0GW4NKGc7IDESeolSwdIFX1zBL1gJP4yEyK9OmozbrZy
aPFzJHjcPDksHcaVZF/pf8ZF8pGIIFjMu35uwabFrbc6y+Gy9nFCwiYxQAQKVvWLXCcNhG27LL/T
ueCwHRewSLgqWjj0k1yJ5WTB23Z+IEDYJtI+mH9ZFT5DpRSE5TQIv6/KyfPyW8vdy7rnMb45P744
ZVFBzJJffvoYicei40W144DdN2D2SboyDgDUuSu2OdqkRm7TvS4Ftm5Rs6Alfi+Xu7QKV/Ud9DB1
32vbYp3s/oWL9m6wAm28fr69DB9lGU7unqMiR7T0PdAjtGXwl4W8ldaefWISYZ8vI9+rUMDf5hJq
zmu+ZURVSeU25e4HkQcr3mbtje9kP0fQZci1lVQOYmt/Ufv/xWjmaJJ4SoOxmOIh4DJ6LAeCvygm
VJW7OFORm3zPvfRutiq6BzELPdH/wJBELm3xJFHFC8tQHRrjfH6lf6VSKz8diUA6OLmMYHw+GlS9
peMVzH7sou79VbyjUo0gehuAEm70kzMQYJ6eP6i7gmPZbp8AIpH4dwt6JwlCg6MGxVgTT6oMBcB9
kPlqX2h2/pJyjc8sS2G/nvciT9uphW4CeTYRAW/uHc81IH1A0GPlpOcNMn2UDbz8WYacrh7DBxIO
/96MK69UYw/3HWP1eftIF+5XMw3EfnFJ1BLfuJe7YovihYANAF1D272ps7yFAXXn4T9jtDf+r79w
+X6VS+H9HsTUporpT7tOPps+Em4F5Yz3U5TcLw1LdXzSZYXcBj2jEmTB8qkBwWRldgwn8zT9/DEC
QqX34mheNrz5/4rjjUS057j5BYwFtVdG6IIoefmuAhYysz03bqdWQmQVFC/i5r8OTU0ammHzYCQl
IT2bZxooBbR9kNPSwhavn9BHUNN7J5kU92FAtxnD0Evmsrm17JHIWCchJeQlC4dSiBmRqG3F1LNx
c3GMGet2FUTLq+i8Y79ETpQuaSq8xHjVEm4lxhQeT/PrV350kG6uQtsMW7DYZ2gu7TBhPXr0mo93
GnpXYXtlo9lln4rwdNPHwsGFeY2rC88pgSAJd92PqYT2rEPTes2cZHTrDVabJjgRnrUCOFAuywSR
8/M9tZPyyM0ayz0etSn1TW4Ot7upQbVYKrHlWrhQXTeuRxjJvFIMP/dGnoQ4tdFEnN3kIBpl+1K2
SULH6YdGiVQJ9KvyQEsr9yAiv7H9HyhGTvrcXjcni4z9cO7LtP9Rk9vqMedLrVih7GAQQW5f4+up
bdFMi69ELTprcGuxl9JrlFvLk4Bwi5E9WGeFu6X2HxQuzIOmwDUw8pOJHu4qmOB/XNk62olyxP9C
Z51A+oa3DVW+SwytHIjVu8RaXlL6Z1iYMiQajY4T9l8WGJurWUx3ShArzvt80daQJnNDiQl5rK2o
o5yBDYq4t7+coIaEMvLtah6XxEET8G9PqvbfSS773V/rG/JD2Drt/JOTbeFC3q6B3FPef68RIwIE
BTy5tBt+QyshMAKPq6FhQEii6PG8ZjM479YkwnFE3Gw9cp/Fjqm8ryZTxaw1rCbwhIsqfcKerD6d
1AYZmfUd33AqSvOm7CcWMbEpVH/8N7Bf/pnQO/2Kv4U2e3K7yTLClR3YZv6+JmqoHa/QINMGgqWt
hxAQaLlyhhmc3Er+9JZh4csX8IgyYYHp12aOgUwC4AIjjQ0X0svIvQZHdPOUOhmKHjHSO3iMIlS2
IZ5SBDRO06wrV7FNniCi50D4q6IUz3V5cntuOQmrBrJXTFUtdgLK8s/IGIqCdaET1s789k1g+jAL
iQv5gqp8JBY3jrhAnmwgfKG/t0SU1J2lgRnB6rMKvbbRfd+Qs0KRDUSLKqAuYUka5O7xHJ/p3DPZ
h2pKGxPQpRSu6YOc3qMuKgxczV0lIceDJ92aSJb60g1U9EzvJ4c2TSth9gOOq9ox8eLUQ9EH+VUy
fXpupgP1qtQrynQJ7UfkP8XIdhsgt+12asHYxKxnet8QKZLJ05m4nkX9/UQB82XY4oIFEYBh3Kmz
g2YFZJK4uX77N3U1RUNOriHL67uwGMMo+O+6o2kghkjbowYqULQwzTESMq+F2h0mH5jmRM04avsN
Z09hH3d9/ezLJpck/frZQraz/vxfzIKbblFXvV84vZim8KfSq4RFlLLIv1y08xZnfikYFmnu98cb
81ERijOUw/gZabu0uC9WC04j5u+fO7VowHrpabRlqgt7Ndh20nHZChc4508roxAob/QXIVXMlGw3
+Bcfz5yBp9aaQwiBhz9qbLg68SUUCWSSGNcWSqYlE8dSokKeCU8AtpVBywAVmGEFAaMp2VrtpkTo
1DAUCARlXklD70XodNHU48X1w+WrvLTJMTcJoY34hJsWMgoAxtNjkd/A2bg56K4xJiPCfqNheGDZ
EgRJe9/R+9TZwgg0JU5CdEqbZT0A8Ok1BE72wydNyRNo/5RninHXJAfUu5Y7F/fx9q1P28FPMQn4
HryUhJKbXNAVP+pGZNITGWABgkxbDLfwWA+GW++6sud1ZghBWPUJG/3khPJgD6IgOelgMevdPfnk
+xYRsksHgbMJuBuV5EP55K0n1aFFFue6N2y4b+009SG6OzvzgAU0igz41sbnFiqMEoTPcEnWi6gu
IyZqtsRt0zSQNYh0N0Gk1mu2ePcUzRzZeqPExhXR3pnu4CAHXG241GucRSi2tz8UmfZQowWu9XHz
qfL+FnSFWLr3lcsIOCliKD+vR2UL1hFPT6SozgdvfX6F/kjo5TJjv7uXqm5F96CZTb0wzzztLTNK
3R5KrlipmPYKCPD7pZqHgri3leq+v5KFYoBI29s6VRsk0QgMHbspXWiyz/VwD62k6+f6Vu7BRD3O
9ZsV4Y3t/HugN1XukvZClfdchDG9djLMvC6+c+i9dLJi1mSy7PyMfO56w/eflt62qCTaAVnMlJNH
0yXcOG5x37/3/FVAQucf/D7O6ttOpMigtEKAmkajUiH1AMbh7qO7Dz9yCB9qkJtBMnExCwNBpgu1
Acr1g0w64Uh7Qfz11OjMhkcR/A6ManfEPWymJC6xFFub9KeurTVfbhkZHR6QodKef9//4pWHd/rA
tD+Q3Bfp+O5cYFIseGkebmrnzfUktyJKEQvnBbcGHGrQ6PdvBGvvSq0sptG/maez8BowoLbjF7zg
osWU89c8CFBljmwG2S6ji8XNBpRprEKQeMncG2wtPLm47kjwgxEcF62/3sOru/9JfMVz7X5r0qgk
UxMDZ46XXK+wGa72lqOgwLfAH/4wqePji4lp5Za/XeiN4+9EfBM/BpiS79+ufLYwbq9ImAEcdaNF
TafLVQ0+Q6qQz0xW79F9gu0CVoDnCFxGTJ6prA950Y15FHos6FctQbhg5kuCG0pV9T83LpqmfyyU
JHkbdUaPcXrRoFEFS+gjAdFSTop5rs3sxTlLN2HhQomhetE9AEHLcNuWrRGi1yRgAfboyJhQu79j
IU3ovfkBYsJ+463VSFyyVK0PEd+HxtOwGKreAqY1Nd2nXxGaHJzbpS3eOVLk7E8UI8lKB6xTHNLc
hc3yQCt9CYnId7QOqi/3lSMAW1eGbzUBTntURh16i3BBTVgt1SCySMzVco3kodg1Jmb/11Kjryu1
y1jqJpZ8cfxkhscFbEm29W94djITuRBMZTxj7NBFX4uNoa72mmCx2PRG5Yj7k7mNC8iPs666SHJw
mIwxpEIU5pWMIg3TPnPLRZr1f4WSUmPL7sC/VwIzqsmDAwsw+58R824zrPjXZ/4CK0FFLjZNV9za
uSDb1bEd/YCMhZtmwZL1PrwDZCSJhc6OksffYk8sJ6+KHkyRIRyeSh2f1Sqsy5ldFvuP9PhfhpMe
vNISqH08Caw9RT6rgxnjiWIudFrbvVnnuRNLJYFdzSnagYrSw9LpNaw9y5dyFQMZCV2TFzeB8Ywm
jnZcci75bki64Fs6qG5WlcOItZ99qyzOkVDg7fXT+3wflA7tizklEl5TEbCWniT0MHBnz1vaqmut
DjQ+2Ydq9uWx5YdRYw69D5JPPa5HdQ69ZGhLmj8V92YExXU3sWsvDJlZHJaiWPZt4pRFJeI2PsCO
NhrjjSpa1RNFBuUtWnuiia85mymwHvI4KOtuIQVCbXDUlfAk1HLv5dIos89+OKe8j+Fw+4AgHeyt
3xXcq47HfuMQocG7nlma8TPsdeKOauOIcqgwinlbW/zsqWb/LFTmCyCOXPOfQHDz608sv2m6L1tf
/Ml+tB4O0MgUZxI8qiC1coz0rbskcdhRMucIS9XWcUIrcbA5m0ovA6PhDoujALBRYzeReQ8+nNlw
9lDkYJ9zeigbOU//04PUFCmv4+uOIkNCueN4l9TLn5SXet/taRAZX2WEhcqWeDTm88viDFlAO/uu
pODF25+oplS8sf8pQfOwVPtlI6XfyeQ8QwlziiNAZAhXTTP/pUe6nGirjqP5yqlOKghbqSXdBaPq
P0x7QeIn9C2B6S3uIzc+1FsunhlpHChE78I9AEQuwaRA+1eSd21mfxq6isVHI0ZfwrIG8ej5/4Gq
XRxq70+taMnXh8qYnCDTOC68XRuhPQ1F07jaHM2UklvMcmY/XmwJvrptVZwIA/ht6OLEIxkVtWH5
Kv1PxW+f16gY9LEzvGBoapItt0qQW9p6Ek+sLABC88Td2v9AeXVKEvrrjXiO5mScnVcDQFBYcZkO
zxA4eOKL+c+Q1CcKdHvwVeONsN5fnsO3CwKqyy5RjyQSO9GY5L2KxnNrNoV7klrrZkuRqaZGfrmN
/V7mmkFqh84yZAhrO2pzJyNoJLID6B0zHCfWudtVUm8461MN2+WSFGT7m+9+j1cw2dx1uZAO93s4
hZsVGRTbl7TT6Br+kZo9r3N1h1pS/z2NA756BOBteaW8Ey7S4Nqpd6o+SIX8vwtnDPW61bOyojoo
gcElcKlW2utDOG9PSce4bAS4XDx8LbqsAXcU9G3iD4xab4CTJPyTbj3B0UFrFLMZ/ehNdNeKovm+
es6w1f2XajKXoZ+Rwm/7jACKSPPq2pnxQd0H98P6rRvtGaAz+m20DPutq4o2z9otopGSE9k8mANi
9mAxWg+PCtXYuPM3XwjSDudVF1hqVktM31ywoqN6ktFnoosNKdgyNTgLNdTgFrn3yRJP1LnmY6+3
SvRrn43Pt76yJ/bcd83lc/MBajf8ZauFapca47ZPzkHiAV4igpLti200JxQlNTl3kag17XNA7bu7
2xeLdn8QkhbS/lKFzrXMHmE50Y7E3aSF61+pkchRW8Y6Pms4p6DLgrpZrUgZNBRuCBmUMN1YDhYF
G32I9VtD4sFV3ITzZgLn9xtfPqLIj9HRHvEUPfmYYKnWadTXsjC3asL70HXkQ13/iYC3lb5JmM0D
ETGYm7d7xHgR7QZAIADDmC/a4e5najPv3crsrAm4xvBETnxDmHFB6vDHxgI65qcD6pBpYy0IoYBu
HSyE5bqCPQPm2g1nOZyp05nzQ0N42WNQ9OcRXRHL/TuT7dPnr3Fcf/MoNXBMLQKBbkI/hI6klZbP
qVbxDgrMbA59SmbahMqBjSHEMVY+k1HeEWbF60eP9PeAljk/DinFKydSYBU9/UjYH9d73+7tKzX+
Qya/vDX1ZvOYX08x5fkUIeR9XxpS78Ju6fgtODWGtAiaEVvH6Qhy9p+1hUFlA86QaT2WY8ORVl29
lhTzBJdZNR7tftPrQCJWW7StK+MmEGCJ359bmoU0+EHqsvz1qrU8AEzBYFhlA+q9Frie5wEKEIEX
HoV9UaAmKeIGDduTpDi6OPHO0z6f9L6U2WT1dokebmNCoH1syDh4LC68NTqkfgR5msgxJome/AA1
MtXATwSMmg3hCxgckR0tY13d/eSjV7O2vYGJmDpMf9OnNxL+QJKsWWaRM5mtbu5EWpqbbfxpbSyJ
+ijN5XNGqsiS7xxrWxKHF8fxfVeM1NAuMxSvmMQ4tDHdeSE7uS9MkCu5rZL4rXap1sacpMoC2qMW
CgyapwjArwBWaJJ6HknTmRZjINGYunvMrnEdRIORq4YxJgBkpiQLeo6puXVFoaHBa84CRL0WQXFh
W/ytwv8EO2Qp+nWErt50gdb12bVKQklpXCOfARxvEVpDlHeiEG8hVix0nJdyhcSrn/GyHPDzaW0I
EeNQlzdQaIl3EiYfkx5OTWDO0Jgf5/Onkk17kVan1I/zabADi2kNWWgSqugo9QFhNXrdYRQxuOFx
JPXyuGDjh0EC5Uvn4MF4xGielsZYz3lzzN5t6tZnY6NyiXyA++kU8kkI/onNaoHNzLGJlDl7QsMF
zQRIZgjwza3hiT5SatqsGCQ3DNQgtDFnrLgpSkeZRCSAG9vCMa82jAC6+xlITp/rijfuRaUppq4t
/dd+e8G9sIWg1blO+g3bDOJWQjs6nbaZFYNORMSE26WZesdl/v5cBCmtQjCTSmXqh+c4qRpyqOtK
EHtBfM5ny5ACknakMp+dq2XNB5NJiH2R1mD60HcDvIXV8d32BAM8KZWnQwXFURErXPYUejggxTIN
MGAcpqlXYdq8vT04ama7rPsK3vrv8PYFX/o6NjqlpyTju0eNFJ78s7Tdq4LC+WyJFXCvZH+iTz3e
+jk98CASYoGWD+gxWKRoswZJ/AWILkkRT+NhbUkvTSHwGJyMZoDt7BBbASydM3LwlkRpZhEnmAW+
FqcbgAWhIdAEozedMnh8MqbqU/e544QfY1syCVkEyRDbxra1UBgRdL+q/1TT9H6ofxh52i4UX5Gu
rvvmDccd5OjAZsBZKnZd1uKcjhfuLblp7EDDVuIbC69mP34zRVXpmEDKL6nlo/pXrGFXeZlIxsLr
K8hY9Cp/8oMMFXddFD7uozrbQ/Z9rkxmYhkHa6hlCNCYxQRXmwGGvmOKu6nVezAenn1rIH2Zhluh
dZxNL1wRpZVY/SN+XCZeUSN/JslbliATXhjQF8zq3hlMQr/fV5IYYvhpg4QrX6GNXaRzi8E5vNeK
cUN2G0poSse8V+UBgwkhhP9PkzwBzmTllD5AKFp9HxPLjxxiDMf+v122DqUpCa0doAFvWnxgQzTB
xMRi7rCJmvvsnbYg43370vAyb2IYero+rlIAGIYsh3VLa+D9+YHDq2iMHYWl3G3mmWVBiVYD06qh
AJa5ZQFGMw7i2GOn348ehZwE5934e0G8nbUAcjns2InQt6TCqjG6latxMIyytC3phi+zwb0xz5op
diG8B2xtXcX2yQbF7uG4YL6hBeMqRjbboQchSrq7AEfJTD4AuK8JHzEhxXb+1SSXFxxD9Fz2v292
tdrkrjbOwPXVCqrJ56Lmz6xUNmgX31BSEPQj/l3TUuUyL5GqiGag2USekimwoB6vX9qeIUwTgbnd
BDjpEBfS+ox0H9d6vPa23AqJuQacuqc7K1ICYidAIh5GyCC5eK2GExAYbWlcWbFrmO0iBqMc0eh/
qKY3f2uSHUX7nuGmsdnxlvT8wcpiWXRjoEbkNdIbuYV1js0efqjEE+J4tuvwiJkRGjcxJIxeX6z0
R29Udlethg+WODnT7tra2mE5UgR1pMsRtcjdq/aSvwTN8XTOrHJRNZVlM3cg8m+zJc0NRR9A5O0l
whSzx23BdRWdY/Wl2p8wlbAaFBFQrhV+oiWMAZ71gZ5OfimF3UBtpGlhzbsyj704RnWgoBjMW5LY
0ayOSNO+7n5NmpoNix2BVeV5LsmR+9orjAJijcPz4BL6N5lhVfGi4jQmZi0gmzu36jTfeYHn0UnK
soIyQMO3VK+D4Y5KXXYmXC44ycyO7M+DC/kBWvkQKPmfv50gSqSBOmA2w6LuT3CaoVr8+0w1dD+C
d8Hw5mTnvXm6DUixMAvdvqaNU6fR3I/8dLlA5XDLri4JDdd1Gr4HQgKjxi9anSYKOEKjFQHtUMeL
I6T+/+jSYu2EgDF02RxOh9dBJnDwippaBhZSLEsu/vswEYgWA654nQttWAaEc1VOLLzTqIOqFmUS
DeEafe0XdK3eWvros8EeIIY2+cAHTIRTqiFlWZnEi057cb2cYWquJydW11dl6P4ltZmhyLGQZ3FK
WJK9cNApJefEYcLNMupu/RBoW5obU8Oc/ssq6UBUIAcseo0dQErkCtzmzD8qNUPtZl+iEd1QBtkr
7BLDUKwBIX5tAZqKnjNk87dHqfFuKkREeA/tllYbXjlBxxDxAABRJ3gn/srI4n/rXhgP6eREfttV
bOElE0/Oykp7/YbH7xRIF8Y+aUkOLf/1hJtBNwTpzCc+FM7p1JWOKlkuIezK199oKNYOGLqP2y/T
V+yODdCxL2aDJCt6tNcUfK71EdFGdcvyVnDicQIt9i9TaSPGFVMp4rwxq05zjB1aTYLGLi8WpSQU
vS686rIKh0oharBD6+f2s6Rx5uFBfyEe01ENpbujO2N6ejz3+nGNuVRNAggEEsqEmCFdh+LTECBE
xroilgXu3gPbh+2eBS4KBY5BkXpINe1+tCH5O7ZDeGH2ADaApxC9o6nbXMIbTLXPzGrx5YvmN8A4
lk4eFzCD+qx/NYXwivo5nahiAVT4lnUBueDavQqA76YSkNEgTKNu0Q8jzhCzxjn65U/mYsYgnFPP
vlZFLyFmdTZw6U6fRDcHUeTMnesY3yF1uvttA99vKeoH/urvpHthUGqu8r/qO8uLFZCAi4+zGQpa
qe1lMgIghKdj/PhHXs7fQfHpEAeotLrXUGKMXPIPgiYe7vJxOLC+EjD2+xkr3wpXl/vzJNjIz0Dk
p0++vlaxeZgl3oDGHG8oXmJOMmle2iFyeGQeJVqdWbWX7QsAXdjy35DXMNvc3tXpK5p7cP5Y3cv9
X7t67Exi9sPtJuEX/O5xWsYhCJUxQGn1uYr7uj7+tHbPOyMQN995dR1nuzhVJByeMox36BKABypd
RDIIpgTRgp+N0cmnJWJo3sjPfjdDZhyenm9tOGj3IOBqqS1meXSQ/cAWXDnWPw8OJymPN8YJZNdm
BfMYnjwy0WeHpHfM9i63eU3HatwBVy7/CHep2y2zynkV/ZsLd7pSVQ73kakiyLCf/N2rytV3tByG
zmhUTZIDxdVpCTnWmPZnkIssHU/Qqo9HPeJjoVFh/g5LCpsbTea7oLbTfAUIIAVKYFGMkOEOfMK1
b3xVKRvd55H1UKidUHStAQaSvO7EzxsTlYRjfDvedAe/VGaJUke/8cARlgMc35ptRz7wGPq1vctG
w//C6sZSHkNDZzwG6suiyoPfymma5xkZAyF+dcStrKjhMn7fd6mz4rUa4fDlgWfjeOlB2fc3CANV
I9LQP49vgwRiK8CFvh2H9krKeFe/o9P2VyhUBcIhQgML08rZ8uYmOUfGSs2GO6GvsKNOYgP59x2r
uiD9CZ2c0YAGF/Xh44pGHX12ABiInLUNPmmn8iJcJhdPth1wm30kH8GA6FUVmklYAoF1lXq2Y7zs
6CpwEWJ2XzoTY2BXA0myBUX9eSoFeGJhKgmq6WCnTsH+AW9V5zMO2C+s7yap8mQMRySLbfhp9oAJ
J6EeR9/At1rrhN/S0ZrYSKJxkO6ssuy+YAU/ZZ20Uyv/Td224BxcsC6ElNEdjoM17oURJWv+CP65
5Y+sm1wCFRE0ysffHmYXQRgD9H2h8b0/sXIKPUJRz1FfgZbs0swscoyuNlMTjjz6cTN6QGxt3p/n
vqobUlEfa08ftJ31iw3P4W1yVBLd4Gy+DNbcGVhfXVsV0BOOIGj0GINP5Ue6St/PYDrClRjdzGbl
tzuozpDC4m8dUC6nyRMpNqAYn/fNkNoGJNvPurCc/hy5DLQgA8NhF+imzQ8946HHDcox0VJ57q1d
+ZPRlLF/V3gZSjd34jK1K2pAuDc7vzbdEbqoN/OSYERSMFIdTC2hH8Bqna1wvtWLJLtUCI3SRQ4/
L9iT1ZnUI0Pie1y60xgXjR5gDWhb2GqFACvpjzcSuPYBNwD74zf5+Cz4qgWsO5Fb9Y4e/Iu7pdDR
amj/oWGPd67/iVZquwXFx9mw4VHr2a7cXynv166Ja+LjznufSqBAII4NeeSze4EcY+Cw4p3CHPTD
CTfFT0SHtW0M7x4q4BYbqEQWMf04UWK5YuJbn849HBj/1uKQ0/oWAafXyE4qKyVAiuMcgxa0CCpu
2+Ml5mGhsQ8T8FwXxlCHNFXzU6vGngZQCNnVUGqqiwlo7YjGYIhqZxXjad9B5d/pLoUq6ymmBfJB
IUiyJXznYNWlNYDDmJZhqYtH5kDMY7V4nofx93OmFWUhQdRGeydP9yjfARyrWB28t90/MRUuyOg1
tH2wFLOUnvAJtjrZ0rtbq7EK7e172cDTA2Zv67Yxd6liFu4X951cH24IvQEIPkqcKtYLu95UkXwc
wuf0lFwE7EsgivdsiJ2QRRjHoKu+a/s6al5SCG+xpsGmUd3NxpShVG/c63Tg619p7Hur/Wt3LtEV
prI6sIGUY44/dTJ0taZAvjkk+rWs2EJ8Zjg4GBx3lcZ5ukGJQeSK/ydOuSnJLdYlNVsMDF94rARy
S8rO0j8x2JHqv93LFcu26A2+fYc/RjEKv3gUdmCUgw6CY0q8yj7SDsxqvT/+u0kcAORArE794sK8
uZcPXfyuuKyXpvn+iX5xtNkG+75cFnq7hBdaWmOjNAPjRjDiGWypT+u944Y5j8ldc/rC9Zkk8ujJ
sGKTEqdFAFX5a4bOYAjxWil29kCXOlG4GE2glBE9KjvWn5ILoaNbh2GCuoT2ojPWvAJI7EWKgLIo
JTDy5AozwTZCOPG8WJO+gHVNyGne4ZxivE5Bk9GvxcCp+4yqYpnhaIlHfmklviNzZPmsbeX3eIHK
X0DhE56k7SF954ixNXi/M+u3z39Nfjaq8+CniH8W7ospBnZ22Lu6NLcce6C4nnyGBCtprkARWfNJ
vwzWAfc9EpXFg/VSTurlzjbm6RUOJdrkzYyE1OIpj14tt72OeldFPH5rVgC8Kz/chJ0fdvcuC0vK
E+PbrwQIiD9VrIqCegrDp5V4D4EG+r1B+WZ948lHkMS8xdw6UxGRnEDVto5S2lTPfPOY2YLUC4sL
IqIZXGdJd878PqsvAthwKb2mkpyezEZMA3PXnVAQl5RhqegMyhOibhI7+HqhYNngOLLIn+JFbyqK
LP72KIZOOio7ysk7SXckBXCdI0nGpiDE7APuPkNzgH62VNGGURdRZARVCpFUnQuiHpWtWYlou7De
6ZKokJKP9OnTllbL0xgw19xQU/iF7Pbgm8zmVa8KaGXBmd5RRW7sCUfpmZgm19vWCkU1jOLsRKUL
VAuATpO8L6mUopIJN3m6xwhoBsui9hExdWHnXtMOvrvCgTVBSPq8wtaVY+QZvMFlqg8crtQH8/OS
lsxPKrqgpvIQk7ZIfVa+i+qsXEVRo3Wn9YoZWs3BA6gUo35QF1aNxug9mZkEZbd2vCJqyMQuxhkn
nxMs8Mj2VgmHfClCtvRxOglRRv61WRgYtoY6uIR+guE7NNi22yFSiM8RwHsJxpazosjkD3blGxD5
mTTgkAUETmYLiEDHofOkLQbRi4Jwklt8ERhRJfUTvav8qKqv8of7UgE36ao5vp4ezvUAYKDGn2Lb
3myBIe+Esg7ikNym0l8Z41j62iJ3IodDdE8V0BsZgqEnwBXdbyLzF6H/voRRtgtxw2k+s26QeXh2
A2LJCke+ETms72vR8Ay+m4VqqJwTDafmA2+adRJz+d/dqXwyk193flfxPOgSQ+fMGubW242IEs1t
TVM9IEAazbk5mjY6O6Rz4NmKTNvRIHtiCa/Ymj/6IfWeOQaZyNRRe7TlDJuMfAm6s0zprrX0GmRY
O11obQwt0WSNfKydPbelKWX9XU4Hk6xVzHqJg15I3zkl8q99kNw3v26f+7wkBuRDXqbArJ0wIo5W
CAf8H7KcakJToFWIBgXRyI0f+uNSJzn5K8mJ5CZuDP8yYWIIlljgElA0xCFcwHyOutxiCWKZ5zDP
8o5dRVFzWbmHrZjDZthWTPWLl62q8Rm1B7HO7I1iE1LFW+IrOk9d/kdqulSkQD6gD+qBSdCWlwgK
pUZvLFrRg8bohn2YA0yU2ss7QlkAT2Ko9DSKwjpPs2DbHlT6al2qjny41vw/NZAqHO/wDjWupQtr
P9EHW4MOuQaWKLgg5IndW9o8myIUf7oH67iW5LpuTlCi3s6iNt7E3fe09bLO1ap8TvGo0ShiL6T4
p3KDHc67DpFJsY+1vRUCoKSOz83nYUpHoO4zZa2MZBEePM7/ii6x4VAcbMjQmPKKVTgR7BF2o1oS
mSzQdJxjgyd1uthjcm1nGG8iBzjMteybzODMJG8pNk1BBWlGU+g1PzBNALxFeL4EHabbAxGU+l2e
smK8keNVKphBCCgVs3lhg/ZhAf1f363UPfcSSnXwna6Bc1V9I4uYwG/HoirYDtU9Ysy5Pn1KS+JO
QqFFmS/dbwqaGQ8kef4MZgeAjqLS5zPptN/+uzckyThyRV/fOFCV4P6bQ78mwE1ReppilgL2N3I2
sw++9j71Zk8L30Yx9Z8VQQUhjT8TX4QBuWcSGSXgLMX4KVwfN/k31Y5p1InCSkJs2P1M2sSkV650
6+P73H/ENYoZa+OQn/RKigcetEE8AvUpZGNpRYZqPNlQrhv0AtZ2xxc1mRkmnlU2HaexWr8MdFAj
QTKlkNVpMXBo/S1NIEZudB2QNSgqzBnF+Wk5t+hksruegYX8/2P7FTj9AuKh+GYIwwYQ92q1fn9t
Vl+iQLNas3JWrSZwpnj0O79RFELUYN5jkQa3+Giok67x4ojumCCU4d+X/gOQHHSkWRpiruMhyIzh
Gs4ZwwFLxbza/b1flcYby6ehUa0lKWK9KAYxXVNUSnqNyVhiIVNWbzV7kdmAey8TeHnpE150UB8j
NJDav1hW8UpH8DTZGDrh4sd9J98cuiK+ZNvIEYsBU01/EiQLXPQgJrEwT88sBMr70TiuZOjaBx3T
KjjASmci3HbSRZD5vy9yDlx2yQR0ndENFL9gAMMGFaZl2x6XS2CTRrP1xnIrT+hKuNHGUUznolDk
N5Z5V+z2iw7JTJmPq+eiik+s2qlPQRlOaB8MWVw9Fcabq1diXofdVlYYNmpVjCu8gYD4MRHeLb53
aQdS/0T5iq6Sr5/2EE8razI0KvPNddRday+A3n2KAT5KUTO43LH30+jiM02sdoiXLzK/qSVOYEZe
uYVkykPehDXBQAxyyntT2kqRXHGyn/HCrMdvnslj8VYdjWzpowfiVuahnAz1YZcYQYQHAMc78LmO
VBMtUM9o8E5wGlKihSbIpCWwzv3XF6WBSCPF9bNz4lSA54DMufFcI6CViBZ93rM9+VIalicNqioF
Y/Ok1db4ewBnTv7qmZ1/7pmS/TjSfgFYBZX6+z8b3cuKxiro+NQDq3iHDppeNvl5gzYhPOsnolgf
6OxaCLxbvwkmLh6SS+8KebOUcWFSJkIEauZwBxN+E2GK0mVOIRJGg+gEbpOsf4gH8+bboK2PjHQ6
ISkf7O/OzXLiLWwIcOA2u4db0nzIF+/AmZ3w7b4cS53zd4gLyDxTuihyaeZvGKDK+3EOUeRbDKgb
KkZWRegmF75IxTRt6Ryujv6InmwLwjRFLYhOLamUfDU8vM2apZ5QuG/1nAqqygGVThZzorvIh1tO
nCjEHb0TAhHU2T9KwPB4BBt2q+24MYXqd3lpgsvp/nQUBAa40H5sWn3S0LfAv55kMnxwoCsOexLF
SPpMOso0jj6U4NPfbubw4meOJTI5WuMB02qX8RGb4eWCEsOP5NqH/L5hLku85tzgggBx++302eox
tK+3905B4orUFrjBxq5wPdH/Ktpc7y5fqSTlRLCQMtnldkmd9Hb7mcBbBzpZqrNDlRo/AkUQq/Hv
zS7Kn/ir9xgl8EZU+V/1T/q+L5APkDpYtHZG9dS0uGpFDRt4uZKqUcjfX4y2VCMrpsYkwoslVwta
CNIV/Wn/vrHW0N1YK3pfR2cnPCjvYzHLp+VVD9fVf+mQEwCD4TaUW9vlN361vr7VUBxvybQI1imz
Enw5HeTXpGZsPz/BIM3vyglspJeWV2rVNjeReUByrKlhaeq1SofGkzC4FaFZK7Kjx1413iizrujG
PNyOmGfh1SBJdKmo92SeEGofOzznZ8Oi2uQMipEvd9AuoPc0R6DIMFHmDqso2HnxJ7Npq1mLYbgh
5wypfXlMeHhRSF98XhzNukdt+BL+scnVxAmKDksHV9pjDlcXwmI5qL/Hw7mzWWK6VIEQIkRhXvmJ
kvrUzjk/7qb9nyAs7mn5cAigmj76iSWS/Hw4EW3Lg40Wem/EyAtbVmGqnxI5hdKEF+bfMfLj5ese
HXqOKT3XSFCVpGC+B6dpFwm7xVoHipFxdwK4viCJYiycjO/V1fZQePXG6g/99+NNBngyJjiOfbTv
DuXUMGCHUl1ciIQml7HAsKo50forUQKYKqWbooRPZ5vBftvCbGChpL31FDDMPvdDl3GnXia4SX0W
2DtzGshDq6jTwSWbK1yqVdRhoUWN1FVMKeoWRIQlwhoKwi+owp3AxsI/8pFGyiN/CpyHpxD+H01+
UkYndmycDF7k3k6jyYSgB0Xm+Qgu0NKVSqTMzi/DfLWu20FETkXQKAk64kW6JtizvN3T2/ca03ka
RftqhKTQ07aHbPuHpG+SgPaSmzCCO+r1ZeLzbPYTYTEImajwGs3caLM6XISPEwmhUIRDKEMOBFal
t+/qxFYtYP6uv/z8M/VxYVNfq36J4NkVDlS/5sjXT8Zqmybw3PXfMm1R8j99a9rsJjYfiK8nvHVA
Nk9swuzXMZbiIaXfOIwxqDaXRKqozCKw8BQzavN0wczP7nUYVx+Mr4t2hJqCbtRXz6I1ltiEcO5d
vVkleb/BDw/ptGBP/IFI+nS281kCmIrF4YBOx/ZIpl3r5JlNszqtAIs2/GpwB342/oeYrpSrg7yO
+ZaxwxLcPFGd7axNEA+amTLGEP0ZngqJZofKP68A0EahdL+TAPhf8RYygZ2da5chxFWolzBJ6jqs
MZJnOBMiqRZgG4oYgPcz7EZ2Dyg3Vn70fAYIsZTYUHkQi+Iv6Wxj6mU2bC4zw8WfMgqYF6rXl4Ie
pC8A9Sa8X6ooPZn3Ubaxm3O8mwNVsc+lqUKg/3DCplQ7DzDV76P1qAJjWCF17hDNeQ6kYLZCdIeQ
avtFIYW53nFGT0XkeQ8c8Wtj85V8OrtLl4yvrOJOncciUQNtHatakdFVHaSnQiNg/4DniK1puJve
6vNPpeHrE3/M3beTjAjbsHYfM4xgbMNrWRrquBW1tCwICmA8G8Iw2Zvo9GZ4WazXnwuNsQEHnb7G
7+78qMOg382yPNJ9O+KmWHV2jEa1aU1fXoYH7uO8KrxJhOUWTLfSJV8i8NdpLzJTGlsTR8Bz/8kR
XAWqTzKSm61TZ5TAhWdnPAsbV9BA+q0FTIERPr0DxggdtW3ayynwBYZn/sOQo4u/YsdRkSGeXTwv
/uh3ElLPJ+FPgLL0Xhy7FU7VDoA1XJLaYLvI9vTe4GDaW2TafiwfCQbyL1dJSfdNowt090vmsSsx
G/edD8EJwNec+4pws+DaWgOVT/WIYqf48ANgX2wxwPj7bjmhCuYm41ZTLApm7nbwfUx0YS1FKc/0
fO7VzUSaSqgreA9QIPhCT+yLr1zdn+yHt/aPoFdUJPaqs44CblF5t7FLgGdQXpYOQtoFuaMwZSwM
cFotsxmbsYMmnSUID9b45QoHc5pCwY0/cFFBopqe9A5ky0MKEUkYnf+rxUabo2pFOc5MQv1F1Tw0
n5ARjMtRXFy91ZEiThUByu6M2KTs1TlGabHBNgDHzlQP368nbSurnvz+HDVXPnKyUeg/r7HHDfEv
bqynxb+qHg1i57tiSheUZI5HCJJN2BxcntBuxMzx0hKA9X74tu14iDEQdkbQR7NhbzfojIxzQSJJ
4NkDcpcj/6JJ20apdhxgpImC8rdB3UsA4kKYfpTyNqf/XHEMXdwh0HDEYXxXAICttB5P9nUwUBsC
08xVyF1S89KAo4Rg3alr82F3VNFGypSECjBet30zZH3guT7bWof1UkxdiLg2s1HU71ZstJKkLjXC
qzq17ALzAVDzoeLdN1t9pOtzDu0+86JIKxej3J4/OWyxY0dPbGNkobWaUqHj4zoyQD37KexHkl5b
Bxaww0Bi8e2SMQXg4AZMOyUp98D2X/5gO5inaw0JVBXBaQu+2hsHl59sle8YsSUU6mukb/Rhq5eD
glNi+ngONgpkLRhw8o8rCcTle1mozP8KYmwLA6QJI9fNLL/V26jjtd8voGebk4KB3oDOZkKTL5ju
vMwC/1JawmV5qSPhNRPVvev1LXihGMl28ahJzQPQN2XwfdjHbqJPMPH4qJlcFlI/lHNMs22zdJoX
TneoloyHdhmQ97Duxr+XPiK2rxZz3itraOrdMnAKRBzPR6ZRP6+ix5sDvAFTgyKb2xGJR5GJ57cw
M4XGNahPlhwSWHsfORvWuFaqj9uuN9QFc9sBNwwDDeeWePrbUUpiZCMHLE2Hvfoo1PiISO62Rhu5
fyjeCO5Y5sXkDJTUKd/D0nC8lAHFugRsK8BKyEeRjmbuZijRopbwL3KjQb7bcBX2XSnsBY+N2h+r
T0ErmBLSZRwrmP5c1yY7hNbYGsmkm+lW2hZ3qkMO4CeonLPjB55aLqOCHQWcF0W3BwKYH5gqOxEP
FlT210/T0QJM6MXaMHmw28NTN53QtWuUuBfi6f/jy/H7BUMWvsKSCGqGC0X2yiB+DpGA+ubXbZUB
3eVoUhbZeoH+cRJkBmkyxvFWg8VihE9JEK0T3BCzvShHZg9OQdK+4a9RolrMHkUVyc5AvTUw4uO6
5iQx9+Jjg1xdxbaNMi1dAWQukq0O3dmNMaPQh74ooiZTWs96mWLj0t+mg4m5mnSY+s0t7OddiPyb
gW5HsOP2v0Qk4SsX+qhD/tAVcX6w2B3Ywrv8gaPqgIULIz/BoKee1CxOTUiRt8vkFQbLaoLm4eAx
7axEHsL3Yb/GyO5Bd157fbO+a1KfPPBprE3++veS8rk77eF6xvsT98wWo3OO+dGalEWnHDPujr61
7XXtcYWh9ELY1pCisYkQdGy/OP/xq0++tPWrST49eUEPnD9SrY8GtHTEhioP3PrtEziQFYohYW3q
+J/84LYhSvNl3t50y3pNgYr0c9RBheQTJqp9XCF2FJ6IIqiwuyKQtPXjl/pJClvGYAdRQOi8KNc0
mbp8OGqyCazjhlyVsKdaScCvMu0A6tsTps8z6S4GvXSvIuWDgfJWeq+a1kaJcDLAgNmIFCgmIS4y
DR/Hnxz7Jd20qwUQQjb7uGpM+bJunw4Mq8i4KBudjdkec8Ei7cR1a/JzNCF0kk1/D/YW4WumB+VE
SGM2iyi/dNyrHbz67CQEC+5rWzhbmCer757fbwEcGYy1EJle58CIrK8rXYxoIrhVQtBXupvddhL/
pNvzQEUemouiGoPbII8r+Ka2Sibxkc8RLRMn93ZJKP68NnYxl13ZuChhwaMR2F5OoA10dBGlegHx
zrLKP8ddnDmc8GZ01HZvwKSsatSYpIuU69krVv2jyVR2Xcl80BFzUIkgMXbdm1AzcnXnk2H+JTob
that43HtI8ppWL/k3PwnMYggpqQRS5xRbtse+dsPGI1naGHY6kjiTfYrhnZv9nDbX4RNJ+qF/wGB
TEVEVg5m5PGUoXwuL/Owb29HyfHtrmtTNQtrjzgT1q06DlyZ1tQQgkSshfLG++UAGrUM52wttLjf
HoDD3sNUtOtceiDd49p3NtvnrpkPfkmxfZQ0uh13BsgovmZ/F2xwtn3VQE2qEgrcZulVZ+VW4E7X
862y7gLgVHtifk1BPf7J6fPiEBKWdvoAC5LiJFYWnGa5Q9JhglMbQrO1Ek4kIonFeXj/t6ffPZhB
kG1c96OaBnFvB+qCqrGJkFiwz9O1mNkpyKPSqc/+AxOtyzHCofU0HSC27/M7W3BO4YLIshegqUWp
mi1PwXI9ZLoNtjke4WGdxYlO+eWKGlKpCC0oXm8GZnwbezHEESNpPL22HdycmPhCyppVtLzXnuSL
5H/0dgcBNKCR2+ceczBckh9R9y8vnRNfUAA4yJ5uUcUvKUJnERfmtWVYePbH93c6T309jLS6+iy5
bp6agBV3qImNDGe+YnawR8ngg89b5PA7rB3FLbn1oYMc3OWfnCXGUPym/tncHISP3PVDJQWjPsBf
NIGsYQc/IWwWh5VaJ8P+cFLcWHA+sVLuZIAKtEo5f9XP9Qfs/MPU8f2JQm/dwNQm0PrjmgDZoLgW
1WPUwBPXzxCKdPJ7mXEe6LmcOI1MDikPExp5dpP70QP2IuZt6mqDVBxxrVL+6ZZH8ZFyP+Tx5aTw
t6RBZup32DhAlDNnQZsn+1i/CP+juOGn1KZLeREapd0QIGx8FO2OWgA2JmYy4bCvL0tHl7jVPOLz
xjGYU6cTkDJEjL8Ow8GtajgrOFJxYiWbAFo8Gb4IWtgjsve+YSC9h9RAIyRDrQQYtBD1z9tOpl4p
XIiDCu0Me3r4tALh76VWEd+g7E0dALaaR0Fp64zK76vrBAwyY3ff0tGV/Rn2886HXRrYSCFhG813
wOqroeAVgYNEyQ2cHR3PzkFwNHSuo91pIUB1fwK9oZTJETuLvyFALvEnoNkjjHu5G3lxBoxxl0Sl
6q44spbRs3cNchdx69C25qLNauMtvk8xKJ7kW9hxV8KUzdU+nETXMjznbpJNaZZDp/c6T/exbefi
xsovC2uG6zyTKyxtUvb3AoOrzn2Ulxe1/q4x8xVps4DUmgqpd5pEYgwIJOmziyWwMzrTijwsuxso
HIdBjhwCPvni6PwqQ0ro+2D7wJ8/656VkX/GyrBx0WlWZjC2pyhQdhlaMkrnDw00JoCSsMl/4HRN
+1ABTTLijPjwY0MxRnryeEIiIr/nCiZZRstOsUNtgltYVPpQdOeO0gWfeGcjld1SToCuVY6dh9Z5
uctPNxmRcOw2Aw8G1Mf8wyerGqQsk0idF+MYbsHgbPMz15GjBSbt4NJzhDh1HB/U/cOznKeb1iHf
U3yC9WoQDBqLnb3sY4d5EKXp5J7u4AWVwi2/H6HB6p6O4+RNQzcLQevLNseIy0Ma8kln3+r6yv99
uXpHV8ZVFeXw5tm2Qc4AO/HOwcFbzUVxqLxkmmkFuNeQbqDQTOe3RFcS4Sg4eAVajIOZVjNSe8Hb
CAclfh2RQn5FRYz2kxKbWVXiYShQBaGBB4AdV9QvZLyJMZ2icthvcFGJ4LWCYpanWINPPhqbONYZ
79VopUjweicSDRjk9/R6tt8rMyb6Y17aM7Dj9d3OtBpXdWK2jFS+F1V48W7hO/LGl61DJM+C5CCt
SeVJBu4Axc3BsVKefk2D05drQaIoox1Eh+cPCr2paxI3vwBYqjdKSaNY75iYindMxnRHLWYRmBrl
TrIUatRka139dWTuXXpE6lXUVbudxJiJTLJz4mS8uhYaWuiWAqS9sR+Z2JdudjOisidZ3a+B+zGt
EXtC89trRMghyHR0z2qbPJvGv8CgpqjHN3hms5xv/FxWokp7fHcfMFzzQRrNaIZJTbc3xfuwLFn5
E97S9DzGXQYTF/jU0sYoenAsZI0/kIrxWYLi+IPZS6K6n7RZjImuVnIz4j3OAW6okVD/4zbePUUX
mKRPyeJBeSDrz6dnQRAfn9kEls5pQBpDA6qFT4xxcFR+OLgzOEiQXFeUmEc3MKpiQU5u3M05gwle
JpVJTb10MOo5qaHhO7aQyf/a4bmW33G/aLqxRsAvNaXq4gthg45m3PzK0Gopgc40/Uc/rSU5xFwO
dm/Rb56Us8Gx3vB62EUw4oibIqtbkNvXrl/rIWl9nEgnr8ap2p3gXxEbyumWn+o0PIjxtbPKgtd3
zRmEgH83FSNI6ECkhdAUXIBLaPQL3spAbWtp+N/79/4k3+0hkAgV90YTtd43xmXFdnvZhsVULUKT
SIfnpX3GNwt5+XVtiiJE6ZEOzpUCWmZwi+XqlSgfMxz0+agQK/J/9CRMrRnO5MvfpHkw+hPlss8B
EjlK/a7AvxHKqqhXk1cQhGwhjI6uDXg5ABKlwzGo4gLkiGsRAyEDvqFge7O1dCd1Zdq4bykVQNU/
Nyx+ehT8mFETDVAqqWt5VTm/g6iqYru7IK6odisQwSGu8X2Gcfw2f2z+AoMtNctjLEv6RMnYFEhT
psBT5iC4FnALVvwtQsdntttEBmj0kXg0PkoU2r82YXPoJ1fYaSfg2LZSfXeuszbeypnKQtPLtz08
HEHUys6T3hxlpQfOIKoewMvpDKEIglslgjBllPtF7VD3dGlUiawzXggCQRQgCOJB2w1mG2caAf2B
ByGGyfpAHunPYdBFZvg54nOxD0Z3rnPD7tyOHXPjtaTGBqEd9HwZpMcVCx/ZBoShLvzF+aG7VSXD
5pUomfcBX9A/DErmn6EdqBxitUmf2kXQE1ekDVkk0a+XBwpqbLEN9tPDtWtVI140e5zOgRC2C7DT
BcSB8Rft7QOaxgan6i62fTeX0qFxeICIxwUW90X2kF/UCX25iJw8GjkUKquM+OcdG196eQLs8Foh
seWRhBo/nzy6vyX9BDTXzQ6okXtivaln2YEHLPoBSUEssK0t6k6Zt/PcF1rRVfzEHAhw9bPxG6La
jc8KPCaB5GajCdPopCg4/B4YP30CQaBlSA0I8LO2JDw/VdFAeBQ9oW2G3x5KnhtDsHmxHARSPQst
G2iBDftsSj1s2CdMmQT/jT48dB/6VkaroeyCGnvuZdVWiNa8XYqvpYHCVIrBFrss2u7CLgpfxv5O
oft0gAyNusnNZvNPqwFq8KKwp+6ld+Pe4JFpBbZafMyFohgPXub+20yCixSkgYLKNohaonjsvQ5K
vVNK61jUvEV1awxLmFoiw3hkdPYrvKtg5cZW5Y7/QGllhIguT+ly74ueq+nBgkZ5spRO2ngQXqi7
EJR6oFRIkxzrJHHpFD5F4+dTeVDKxizMWO6TGVpatrMhsYl7VxJSk7V3r+SnInA96OYieJqIFuMS
qp2gwmwgxcf0q4EL9nl+LRJhn1CSnIjiZtWOBu8fK4E+Z0ZIEO/krsSassAt+qmTeZtBZSk7fyaU
lvG7g40E1s3aO8JY/zVugOjex6hunEjuYIz4JYsKE9rpgUTnCGCnQnr6XXgq0Fexe/Jxz34Ivl1j
c04tmJe17EYZJX+0/uh4BS96RokuHiX+DGzhRPs5/HyhdvjXa8C55tss0y78sLde9YfYU6SFwoIR
B2B0k3gR0f6NywRtQOwPCDdMbYszdGD6JP/ZpAxPr+06yyQdx4ajVynefhdVw3/0scpNHiKjELdL
dXVGIfF6crQV8vSJpY9VCHj/qLR21C8Asf9vwRwLwwpuxoe9VFanP2p7oF2MHYTbldCG1faKzFLu
4p6A8PC1N8JVch4HwONYDvlFk5J1toKFm6kWsLlUi13LB0mx48sxGsiQMOqbltQ0riBQsHOSPeYP
LEh6IhQXoc35MZpF0e2SjK52pgz7drO8F1N9JvuUXh5CQ7FYTpbzb96D7a6uT29peBpk78hGh9FB
8GK32pZ8kO9L8QZmLstfSNb3kwc1+KmkMAMg/8ADYNiPCXDVYS9iuMltLaNe94W7ucJn2mgQ7aEU
uGqNBEYO0EPcy7FnWtWLX0drC+b82/arQ8z4bNAzem+gr1mMRdH2mtw8uL+Sd5P2ucEakzWstb8Z
0+nJeXpa3y00jOq27uzenrgkZr7bL555/W1ZwWitj6iH4dCfiUn8EkZK5VPWh9VBivzpfm2MiBSu
F+B6ovHo6VNh3mpOAPe8kNfKje9OMRfu+RNrlq7lpiHL8Z0XUSaleRAnvc/OOh7XROt1vO5ghHem
7Vl3MGykFrpZ60zQ+8EqY8c/9Q0CUX2H3OulK1ONfEdrdZYtIgOS2egkD0yRcZSwqhS/nGrPn6yc
KI9Zqz8rb3+fZVvehr5te6tF+lOYVTYr8K6B45WE90cyC8sRDH/tlxi45ESV9Sy6+Ojg5lMo6ATh
uSzCD36pzhu9QjXZsOSma6gjXF1F8e1UCWVyldm5RsW+OCE3xCLYvsxp8x4dTPUjcHQSoBDTtgRe
Ot7SV+xliHsSe34hHVrXMKfaiHvOibPQ31Yqt5mJQ8Fn9M3odjKIMC5mmwiBkosJIJEPAAkBXLsu
D6+MyxTq8/tfwXylCQ2dhBb36Vzn1UvSTQCWx0Qw5Q/Sgr1lm9jqoxD8Jshct0z/+R8QyuDfTIkj
9p5mr/oU0NPM5FFwCBb49Yyzcsfad8SkEz9xdGK8rY1qS7BBZiXLJ+jX/znHeXvZVxbgZHH7aY9b
aIjMolfLeEP8UoW4TXr+jzSOvymVMHtJkc3RG4DG1xNDpa1RtblZ7MnV23p+9yJAwqGvuAnemHu8
+hYSFlufmmtVBl0+6zPaEW8RGm4+CtLLiLz0S1oectYaGsill1QW1FcKN3uhS7MK9pL6STznf4Zk
uvoI2PSBAlshCR/CNzbWadgKAdW1kHt5He++b0AfTUTAhCmCzurKf9Q03CMhW4fl6wg8F4W3qc4Z
mhQr6VsZVHRElsS6hutKZ33M/6JkHRzNyYWsc9jO+Blsv5Iu+Yi4PkHE3ynkUkPIrEfllAVaKbjU
Vm+3/0ybn8rz0vYWxbBLA7PQzDVQS1Q5I7pZAsMgE5h/rQbZ6/RufRRJv+xX5Miz+tAxfD+vGfiQ
NnyYXIksDVsmw0gf3Maf2LtV5VG8sCIRWV+FsIoCvB94CmW/RwpMlLNgzALZTQcPKcVUtOwAiy7e
CH9IScbfaZRQvoYEslpljFzHExJmXVrZ1bgoAZBGSAlT9ttzNM69WsqphLv5qG8vIIT2b1yBk7RX
BW++gseSwyguhTWNH9fxj8D3qYkZ7PhsINCkQTrccpYjLOxKxENXzofWkgbeJAwePN5bGKuntfBI
8kyr5UdedxDSkVCD44H/K5MaLKOPB7vuFNVZIeS7gF+NkYzowaSWxlOtbfn0C/8LsH5XGRYHQHcY
Zf4DW90vuCuKEIxGka2dSpgov9jD8N6DVUHEgokMQrOfgNRo1vHljs7xWinZAp23RrTR5sh8/mnG
JZoJuFoqZR7/3NFupCCCR6dltYBZdq50t8pQKMcvYB2Gag3pK8d7YcY5/RIt1xm3ev4Yv9KuR4n5
P0P31qcaz6M2T5GFHkFvJUos41N61QHxxJVRHweQdGOFhTr7wEAGodXQ/Oz9s//+T4e91NqXzgOn
pIsX2Ko/MFniR7VJCaJ/p0t077cO40pNYOPWP+mb6U8k4vEHDWf696OL21iB/onskm/p1b9PiUnX
QgWezZmHcn2Ex+AnhxFirAyGbblhdBR7a/6EJT7OA3/DlXicEHcoJWl4w9S+27Sk3+nQjs2aeB2t
xy3+K4XbMsUaVFitXepzlH6HQEuiGofOElO12CJzkMHMgaaqp4FXAL9RBqWz4xlUva7V3qoRIe/O
Y3Kb9jgXc0F37bwxmBCVTa6BXtbgXT3VzgG+ij0AlDnlr1Ulaus4kNV19Q7qiwP0u/JibxaRkE93
z5YVP0KbZnpgfFVrgEYqH2hNOrNFQQl95CTD3h+6depfsqS1qckV6aYl5g+ju8ooa+OjXxRPcevA
Bh1TjsxbCOL1NzEXLa3tdad++cL860F5eG4PxKCxKjS65GiHHNTohxnX7yPDasGgnVb1/R5DwvbV
hcqcVtc3/OOUDfjPLf5sWGoTIllcSWjrhOUc4g+g1rKjbdFpeqwuqhVt43ntjrJBmxtaIcf2uA1D
lPoqrZ3aIojXTlz+/xbOeLIENzW7RIumP2IOoni5i4dvcKTqUzoN99TJn+sk9gmebWwmnS1GucW/
8Kp8Ex1jwQYs1Hy5uYmg3suvWsHP98c0fnOapi71bH20XapRHQgrantQAbi295SKulppUA3cB892
nEG7HRDwQY8tpEkNIux8+MvWrx0yKYy0U79XGp+bgB+9URjlJI5FXvbCHExb4huA4FM+C8mdkzBb
YxJA/fYNb/eqzyg3d0KjmubOvlG8dL9cMsx0sv2vsJ09CP+0jirXY3g8mfD5nRPyKD8EUcnJguWd
hScvJUyiRD/J2ckucGFj71QhkvjGzcWY2N96Qt5El2AdLKrWyXYt8Vxphj81ZXDWRecfmGb0MZrE
FqHNH0S5R6OPFP9sEpAGhNGzlSPUUxyyN1ydaA65jNSIt9TL5ELDkuyTecPjbpr8i9VZmYVTKisJ
HZrrCfkIaKBy17J98qBaxkvJ7mf8XnZMb3yjlFUpJcVx/nWLI02x+QGlf60JAZR1MsZFMUfIFkRI
jcx+wo3qLnuq23EwfGPuN/5oaPGZ8Hnr1NEbhNLrCexsxbbfvL1PyTfs81baGoFgC+B1htfyQBBo
s6vyVc3BRPqX+Wbrtv1adcM4pwJoU4OT3/h9RGn/HarqeT58STNbZwgEt4kW0Rh54E46tCZkxorQ
Ass0+9/SU9+UhPCY6kUrLAxBTMLYIICXvYlzHvm98jwhMAN9vRzLSqe/RY4t3SWQuKkGtx9eC0zU
TooZ+oWwkkmRRfHdTa5T9snpz14Mr0ZG9JEsrAscVLpMtwrcvycFYwAGI28Oq737fqKrDhHJTqNG
9055hVhopUHeEiGX0BgXfeTTELuftncXSGzSh62WD/6Wc47NDoZ3Lunte+Gih/JrCDS3S4MLZP0S
ImOQ/o78beTduoWaN/wu9mfSDmSnSu/9W9tyDLsjTEFv1/RnE7iQ2EMpUYpZsxixUItM69VOvj7g
EkM5jnjcakxpUiYAJLdVHCaJEu35W/RIuD75Kc00KLODsDRLQ1WRppSo5dxZzcEBrTQOoL/VGfHp
URgqdHoOoxzIILPa6IkopmrFTFKyORUkSBpoJSSk9G4jZgCbwo6imZr8Y8LbXE0IOIkiHdfdcmoo
P2M412PeHBq2Qfd5fBYyp2Vr4D8u92inYsh4jxzOYijVakoXY4pC1Dqhan1uYpXBVp5+xaC47usS
+qNalV1Lt3zgu+Q76HNr1mJlKIIJ6FoytTo/8Ens4gOZwU6bCP4bbU6dfmpPBKmYBYbb7YEfNBJ1
dm7fo3mBM+tfD0SthmSwJ7fT3UNzb8nOSjaujqvaFHDKXkNicnWfnpB8+J5lsKxVe6eRZZYzv45U
8mjrU5weUVjfS+vGTX3oQlpzI2ZBmuSrRvUg2BX9Nl1tyOUcBd0qRwGYi+B51B99nxZGWo+eGvyu
mgmJeH276NUPwnparKuoNqbwEvr+922qPXA51k4+vDq8sO+44QAIGO/s7Ff1QM+RO0QVLL6wRK2E
KZT7WfjPaMowFCTeOJshKN2MO9O9QyP9PgOfmlSqWA7LnvJLGICJTj2pxqL94m2AxsO1/NvoWNdT
gfNps6YRgmF9awqKduZ8KNv1dmDWi2lNHkQ3x/uNYj/JNl9H8T+y7EL7zMk5JRCYNHAec3txtR50
VKpqXJj78hQ7Q5miVHeiqT5nRHuC8Dj0Ze4vWHJROHqsWWRm5UB9REMhu/4C5rriS94okuNkDUtd
5nZG/w0hBiAaIh//6mDhBppqeX0cvg8KE3XiSUR7iW+Sh1/ZFqTMYLcRnq3HgE3zmPdKfRS/uwhZ
4uvCFDDZyixJ2Botk4a/Yd8rgLu72M4mv/RFIddKHUCXOI6uJJeaO4GhLEv6kaGcI8DhZuvEyppH
0MM4Ju3DNTcTGadULseJiT2pGPhrvowpyR9ogCEaQHnf4HIFQp5FEQo8p7kV3JtbIY41BRhDVQ2t
C8jckprSQAJH/CkN+AtsrXr4MARnrIs/JTU6qTkQgOVuI2rICcUsjzgIXxlX1/1MmtQP1gpYJ++W
hU3UgKvwD4NJtEOBjDStC7MFeYpopfQ5SrLJ8zBeGNxYT8BBNlp28aF0rUCSJE6jnV0UGZH0CzWD
DFQ5+ThhbxOjYGqxMPg+6ekwkzWqTudz7aflm6E5hAwI999dqwIx4nBhl8XIEAvT4XJB1bxuyvyi
Eh3BQC3f61Ki2wH3uzR56ZNQAROwQ8xKqUNZ3bxhCstZQEkpRtv8FbJlUyGyPb+BjjN7Vb25t9EA
hlOr9LuIJmlQMlVmso11ia7qpQirW8JNCfHvFCx6o7j/dbuDSTzjxlQZpWECgevUwj/2v4ccIy71
g3Pz8rbOOubRbuTvMnByZqxYfd3noHq6mz/zkXRdK+IbLPTjjoMAEwB1Nmi78jKfzLkdyWOYBrwl
OGqacsa5yUy3R4kM9fftuwmLCdaelnYlExgowSdonktp66tGffmzC4hj2borXzSZiMrXDuOsIzrf
Ke+p2DyKAJioKyB2CNBdzvVhFC/Gy2v9/1ooYQfjZrf8dHvTJeanXkzy6c+io8aFBZv9awm1f7XU
fcw6QtND53PYDFFdVCUhhutaYgAvfOQeIbChpdtyZXIec/TLiTKlRx0Xkcvdoqc810ZvfZ7SqQN3
BIqLIVwizZEmpug9FISW25kU5Vq2Hj4HfDISOU0DFFKticUMnCwLD5kn3nFGMKALppAr+wJAKB2y
ilnAJsWoBg9+xzQNn986KiKM/9hd14c6JmMZmazYorW71Ty2rEbskbkJWb5MYcPcts/2KEIIFM88
cmkXujnQNz2N3s1RTFfctVrOTPpgbeokqVwIomWUdYfZIm1q17xjSieM6Ep0bzDI/Dg4fjQORnTL
7EtJBS5o51O3+tZRpU52eMTgHEK+UFpfJGEv+V1JZr8Fyg5g7y3LbomL1pQVM7BTFUsC7creV0Xe
CXlwSl5keXcT4Vl4uJyUMrvpF6/1Iv1SfrCLrcJytYeKC27E4AeRM46JlLOE7foWe+VOFypKHNb7
yJKXUH7b4zVB/0WDm4bielfiyU/uLQn4DvmwJcYm00lbI4328D+WAA7LKuaumcpy5iejOcdMgwYR
4KACCjwTaiqliJQxCs0cugW/MSfnOiphEbX/L7lT5lVviJEZlQRnTQldHQIVU8T/ir5STy/4IwW1
deN8mCNwtms/5emiRvDVlZwj70fV2eUqKnuDUE0aZZgS7irYkVHmKApjXI9rsYyEaGhkx+VSNRzp
EjaRgV0wPnPFmMRnIZVFtok8jHQrGcZ8Mv8SapZDqZZwWG2K94HGlJvbEO0h+CDBzyLaDbhdDQDC
AsQp1nZ5W8NFmz/x9zkh9GlkZQdTAgeWliUGcA1LtBYrG2BRT1FbOatS5a0PgrXvuG4/LjsghuAO
DgfmCbrGqdS+bbmU8AFkZl/CzExuBgz6oBNuQIs7DFoOmNj/StoYmG9WxOFFSwTqZG+o85vVhZ1L
q1tidSY5SvmY9bHwxZSjCfuKXCzPHMmw5u6t7bhOFoLb5Zgo5Hl1VLBnirRKoF9qRHrQvggNxvEr
G8xprad7YpM1bGVwvD2tyvLJ7uU/0llsraXXSvQtcYIuDyZDspPrqmi+K5qrM7tukSn9pk3os8a7
385LMJAuP35xNouC8Ze8BBazsQFimCkLP37XzDZBrDyrSgngOKNQdrjljYJ0XpV2ot3kbNePBu3O
SBMw+zX//GOQoD5arwa0CvDU82E/ymMAijudOSQyslMe7aqRtst9IW4WjLmboMUqPLJuUxBqO9ya
hxyahuCfod6+joITPETFtzoxy5ldaTRHLh1B/CFUsitMqDFal2hRnrQ8HTcwi7anWAM8ixsl5zdv
I8trCddgJim7W4jT2s15wXzbAvk0UbL1doSDIBWP2XFmQnt4nvBOpNQX7TMzJL5CTsIuen+NwjIM
jJ1UU4liVlhaFH+NIveCtP4FvpG2euobitE1C2ctL0QbM+BLHHLJCJ+8Qzvyrc/vhwuxvZzlZaAU
g3mEu6IZnun7qCMAHUZMzYYlX4gBOzP/L2rJREanL8xiOdKiP9kpch3nDeeYoJDBmMJefL8DHqrO
0nVYuu1hUIKZot9n4ppWjCiCO8RjXsnLk+R5E+m6eW32hzDnk7A+yPaWoUdUNsf3It010WN4W7nl
EPwMETj+INsZ/vhsqvIZpczpTdHW0oj8jwrn9CLOSwWGdR8FeXlgZOW8vHTVbFUQSLlmJQLgPcKN
2tOv9eiWE7OymRoxOBNWbp1mqviJbok7F7t+DxWdXqAyGA+KeFi3cBrljSpzako3Ezgv5LtMICbv
h2LTMAYwp6jSXFK9cIG+PO9hMx9QCfqtLipiqQMwbG2ZNpNWDSM9hUNiCNUav5r5Sk9ARDGOpE+W
fqfzlmU9wGesuJZfyuI+e92oytjj17FHVPglkvcNyNNgI34irgCEaQkqxospy14WFTWvkzK7+W+L
C63avksX/hTJrqZgErTmjatqrh027GsQmYxcBWZBXwurseG/TilxmrEB5ODNKXwbbcH5dEuDWV3P
F6jOHbtg6bqfHvUvoX5xZ+qbUeh5g6bo5VtB5iji5kEIPyskOHg8wYxjcO8EDYfysdS+UzeUiZIk
zTp0R18arap0YHCyo3ORfiDHNh5Ok0mxuSQOnzbaXSqCydwLqGty+4CQj0c0VxuZcMrn0IHLv5nr
37ZPmrKjPj1YDkELKPKBZLgH3ZvrIwIyaoqc0WY0wrkhsU5sK9UoRzAUSkIjmO6D6iUFLUI6lOXu
72R21BFhDd+uyzaW2OQKG3K1314g4SNmksfasmRF610tODxs3DBTG7J+Hrm3PFe9LOEBXQHJDf0x
lT9LAlM/34qguWrZ2ZYtkXtT5oIkxAl6zkQqUhOV/4sJyLpgLF77GunEiu4Pf1auP6iTpmbuyAQ5
VQn/r6B4RkdHcLhDl9Wf6Ms7w4dcgZMpItZjUuykRTujJqze5HoHFNXztCAo/GORmgNPSr4jtIDL
pDTs7422TRCH1erzM+Vmy9CqcPTRz6qxnwbNphj4eSuGLhHCxB/6hxicmVyUqEwh4tOgs493AQsb
c+i5d+g2IDu702QC84uL2k0NvyqHw1cKYhWC4mIwFqJ6AN5x1AofjIyuZaTQVkIENSr31Tl5XwYF
a8x6Ktp8eWoLETR8kz0tw411IQQ+lxUwsp5lrGd0DDf/cwIHRyJVZ6raO8lROl+sr1gQzX4bGS50
GQDmfAuY4zX//Mrpy4CMK6Yn3csx+b0aRBy6Er4opTGpcPkzxr6uX3i8q5I9SIm25VcScIQXt6h7
6IET2WXUo2hx6jB5hhfoVmpg4u0AneUqprvVTBaO9OhExbRfjSjb0PYoxgTEHWMQZ8YnbQBZRIcJ
GZhqsnl7s89XSP8ppMb3JHp4CJiQoPELYxM3PkbCQymjxPRX0toj5FNVMUemdIht81jymR2khcbo
GH4yFh1LiZ5t2dR4goU9WL8Kk02BnKbVe4zQZMQATpDmDAhTpCAjknSYJjWWnQFoTq+aCTYq/KoS
Qo9xlisr801djO4EnaO/o0epCCrH3hdRjR+aXdyViULW/CD7DKmidK9FdH5lVV/YuTR2fenDQCt8
fnkq9tskDlc1/JRy51MzqoXfnmR+aSS/3vMKdiRwvKpZoP/qxmWkpHhuPlz4db8fT03YPypBCaYK
9+/8DuZuAKvhotw8agAKlEfaMb2rQfEk20TbxbLvSz4o9ehjsOWpYBi05oLwuMlu+oLYexBlS/7O
QMcdzG72PrFKpgELUiPj0Ud9qzMeSziv7Gw/kk2n/coUPzDwyJBl5k7xx2TUNtejHe22DK654OHC
XuprKTums7qWS0SyJq9Z+4wfqbKqMyFwgU7gfOPu+8IsZP/O3sfUi16TH4hXTZQp4iQJTqUi1tiU
rJT4zn/qwOLYg1ScfmWW3/O+I3yCmiRlu9vzYJKkR3KGiP7ftV/j1sdaLST9y/7xyMzsPRp0fAQE
mHv8Ufgx13BERFsS1HW/9M0a5KxeJejXJt6Nr+hZyq1/ENyvMp4vQsZTDgT8OOZqQQ5qJVOUngMW
uk+5f9hCGiH3sgzrxHWspGaWa/TmdSsh68pAeMXKFmkKyCwePNruRmc2uCeVHMk2s5zafSyJ01KS
tUtF3falHgbhHZn1ZxqgHYrghik9yINk6RlY35KYXHADKOtILpqcd2b29ucr4h0GKNjW3HAoEerj
81/H4Dq7YnqVVf4jyv84HeLApjvg/6TNlTewaoLyslGo84cHlO6KOtut6B+kO4QuwEhPzUVQoDen
U7+IAxV14iSfkYIXR8VKxJDEiqj0IUIv6W6WEgfnxvToLSNWafr2k7BnhEeS40YxzncFBDS0dQvU
qTc495siETd0R1c7vR1J9sfyZKnUlvkbCEBDtu8A2r/GeGf+QC5mom/WaDaPMh0dDfQRWuuTFJHT
HAN3yW0KfUyo2XOO6zScruuoedEhHyJtMjmzUrNv633m82yO8vBO1I14zj2S/2Oqj5/f6uMgrsYa
GJ7ox2nDrjIfCUf0+0ZaEVT5z6MjrwPxbSjzqbkDSFvDoZBL9v8HsvcgvAfpUVtciIdzAZ7ndgmQ
dBNgShQM51pRh+MTdyodO0QzM3Nh6FnGRk4acWVHq0upVMWR8L+6HOAZcvvtT6RwnTlEEJ6+xggR
cD2QZCqFDHqUH75XtV3I1RyDIw/0uYhXzBK7NejeQTTHXQUwIBc2tjc7+UxaKlQCqLH1gpqqGQme
4KBduPf9CLXZR6akFkQuTi2GDs2yOJMRGsRtYMOViK0mBia80ZJRGI+0EjkoLZqLkLyzwQnYqEXE
hXrzgEqiR57F3rgLY+r/xPMWUQtzeu2kxvxBeG8DqOfgQ63JKzYR3/kZ0EM6529V7fghu6M58Jpt
DZfqbeaEJQZJInlkEmNoSogUmxNagtX8b3u8F5weTO0GEMgt4iKPe6av+nlRQjSo5JDwdq0KtyS2
dWHYJiHLDaHnWuwi1Ldb5CVY4wKkJDuwr3wDxH1Pm9B2q5EkmEqroeU0C1ZZXJBOqFfuMKBqB7DL
8TGRei/zjt4P5qawbwznrX9KeI4z1zWccY08WXlQDMyUXnvhlLEoY42WxpdI54yseoS45rIfVr03
ILxmbMJIef42nHjsO+cye2nu6s+e5t4Y1eDmbbkkSrbPYW1O0jR8UAC/4oj+whcJ3AmkAo1ux1JP
GR1BAqYjNjbnBBTrkL0nbu+iGRW/KsJupsSpaNLxwrjiSeVm1GLVxqQ3FQ6sLswQ7m0NgTMGGrlc
GP/rRjh6DmHL7U+8tCMksv2oPGfuTst9XKVDbM8Q8U85MtfbQc2tyH57zz9aLseKfkI830QufN4d
r6ctNtjOxSXrOg4m7CtwD6uisQu3+BMauCVJihSxrYdtLo7x7z3c4hf1ivXrzXCtYWHXSGyn0TZ9
Lj1+uMSg/bMWWDFjG/obQj2WOjIjOLdNJ/gO3Uduwsyn0uSFQQSZGNc3OI1/KX6hl/I6NX0/o7j3
sYtYgzRzI9cErbHKz2fnJ9Rt6TuIr9fP+FbLmLchW6vYpMRMfx/FeBQmTa10UvnGHPPwvBx6UmK8
/JQhnAgjnZkkpvkT8sM25FUJrQfoRE5/fIpvTeuDuoqnQIu/AgY2uk5rIP4YDZ5BtKEnsqotBEPu
mqeW01v9EIKcmWV3dBPWxbbGpL3aymL5m1dmtRUQ6z80xbpknX39bvYWnmKbWOYhw3f0I6SEs0W7
fTL2EhXM29uSDUpXzzUS3yKOMZYB7x1/r+uHHQnUkkHBlB9ZHFhFnfVjHmHCDJUehg0KPJM0ASBj
0e+QSpDCDNaRmcqEwOY1+y+wyMGG9UoqjqhWXel6tXFstiCASgD1L/KMbOBTAFNCiSXx+1VFOd/q
/sJRR9LWqHeG9tdjKV2r9PszjE6QvWh9A/DO5NSKyGMrqFCwDEXQbIP7BcEzZjiqd0AjXQLtn6IY
o1mHQVCMUWg+rYX4+SMHPwrrVuOWLO73U6FPCmuE9BCZXcxPiWmdt4st6qfltptSiFXkMeTU7TBg
86HrIbUpkZD7DoTLhz8bW7oFHRqQxNW3v9a/Nb1GYcZTFwYRyXk5+7hhycl0mzrh2Wc1cYK2du0C
x8dCT8OYsByFfaaHrhg0rbBCyFXKxAUPZS4cRZhR+NGG5OC3qb9znv3FrIVe2SieQgMZ2LNIDs4i
dqX8xaSf3BxvYgc5qLvBXxpHDpgtZOY+oxZ5vXLgiROVGZeSPkkp+bLrcVXjQBxqcZVVGtf8PEr3
ehcHtMbGQ2g3Td4k7FIAahTaJO9SSxffE0WnN7g4+pJLdsaven4VPZJE7IM0aHAr9vDYVWaCn4GX
Naawodl3U2/5I2AppF/VhHHvekZnDKylkf7teOgA3nuGmA/t6BupHWKq5iY7v1wmuBaxYLO83xpj
I48agDCPNu63Pr3vpG9mbHwZFDrA2ZuGhUzhwULt2cfKUp8fR0FODF2wuat2Nvx2HLBVBqez2bU/
gxv4omHuVQ/fQxkldwZLThjZsldvTrgX2BXQXeE2PrtVRT+Ke0jy6SSFghgRyUj64m6Su7FE+Hjj
Jn5LQ8G1FdaHLX1gNlM/cNOfjleAt0DX+ixa9t1tE0arPBCQbi4mTLeBVUCxozg7ZtWb5/OV6yQP
MQK39GJHkYjZirZ8SGixsJc3vpzX35VLuIQPhNfwnkSqB8chkkhKvrApl8RI/U/MJEZhEbJMnL7d
Z4lZm/loNi8WlBNKzZpF17a9f/Vq9phLyb2Ge4GYF5g6XNl2h/3z//GddR3AuFkgO5pcrWsY2rZ7
do0fStCRUJCFuzjKdzok6GnT3s3K7plSamDp/gDphCJgpeNtVAuYS42JI0ndK9X3H7+hzKrUYV+k
bBTa0rnI1mJHWpLGWwa/yKuSNr8kxKALETo2t+tGgZEvbp+k7sfpKfHrCw42DQanJd7IBUY5syV4
1NX9lK9zsDAgMo4hhMiL1TmKTP2Tn89BhypTnJB/IY0AzBMsZEI7OC/SpEI65tDssfoDf4zKU34m
X7nadqIHg2LJ2SO4s1XORXgFydp/HDBPxFPGc549MRufzxCh1fx3q73VA2hfZQiKaTehk7p8vUQv
cyLiFgswnqny2dcvoz6qb/QZNrZ3EVFzY25bov/MxaXiu0EewjBJOxckws9cO+5DuffEPf+HqfF2
9xMjkaQUYv7AYRkJu9F7HPIHsKSmZ0wCHPufCShBIXHIwIMy7LCROe2XXqXWPS1+w7MD98yt2+CJ
eHlLM9DW5BHJ6UGK7wEnxnI/CoWLS/bHdwUIFg4QT9GNvq3STiZs+P5ZSSQBNjirFnCbUTxrzXqK
0f4UEM01bXa6LDoGCoC27Q1H37sfBTfbgwe9HV21lT/4oZLEDC1D2VJgMeP70Iguul4WfvVgDZGV
oL/hA0uw+vvp7xiHaSUQ5MVYyqkZ4mxkPdVmjQppVhrKIiK1sZnaWv2VhNEUHmxSfsMa3WTDQJX0
qabVkCG3HldHA7YzSi/QeKdI7em67u3NMm61f2MyKKQOG0xKZoRVGZ2yzuCOLyypQXDKUMXw+Wsl
glKFvnNmvtBhlYhGFeGUvOnZy9YJrvNx8+jtp/wVDRdEaquSCJVQjL5OWhutVHgmuXcIGigZqjml
rfpICOcSkERst8FJ9ucV1CwV1TIYiwhY1v4HNaFoDqY2DfT8mgFWi/RCz1BccZvgj8G9NZsu0rXe
//dLmMJUEJp/jHvxWBIKzGKEsfmu+x25oZIH78jADmCakt0y4pkSViM+rmx/R8s9owXyTdV8P3XI
hXgcb9mctodRNXCt3jCBOD4ir6nGpKH/uUyXa9H4f9kiMKsN2C9Lxi4vWH4q5RwdS4hIq4T1YecJ
5lDOSimKLcNQWaNh2bJdAWssHd23ba7bqXw35qOHkxKJWljBvkNt01V0d2HbQWWsScY3c1/FsiTL
YWf8wozmb8RoV7m5OtOB3vx7EQzxIGLxAGI0iyWSfgNi+3OSCfe3gmSVaIQCArdkApe8r0zhpa9z
ESPoBiPjX/lyIuxibCFHqLqeKBGKmPauKmDm7uwhhI0QWP6TOiHbabi9qeaFQxRlUQZEKywZbFhD
JiZujPHkRr5a1Ms6ez1bQ2eCI3D94ei9KAMkbyi1nu7EiWShy0C4WRTj7916On6FXMf5NIQLoogd
K4uFr7XxX8gwbGNqI30XMRyhRoGX4pO2wgXphalBpINwoBAs2ERuKasrhVcOUcovqVaQrWTXG5Be
DmV0MhZrHpmMFoTOYh5o6oEUFyQqqe7XrMOlCfv1Bw0E406AvJ5wHgKy0ub8NLPuxncD9iMccTgN
wfYAfbLWKEyprhNtI14nINhMiYtPtcPj6UfFUiVVbhiEd59M3SPCMbfXvEeh76C0H+ByJ5oiMDPE
dfinDd6P5CA9uxxoQ5zt+b6rdyhGUvzNTYDRi+sF4OgjjJI24LuCukUbRy58G4kmvFd2S6EbzuxC
NUEsg/yNEM1mmmrRwk0wNJgdRwCnxyciz3jP4y51LSDdlxCbpXsw95ywyeLA3aO4J2pWImSIbTa9
C3AYyBlrAPFWOEYCVLBAFwuwSb9w4CeIrDkVfPRYnAFQpJ3P8CF9zjSdg12aqiF2T9ZCSFptK7aC
HN7iZo11tjQc6FrlPU+HoUNn6/f3l7LBwrWj2ZYoDiJr0f31HlkPWVx+3sjSPvnrX7oRdS29dJKV
PQRqrAdCFXEUiT/T5Bc+sJHiKK6eJKX9Q/5qgqTHLOkvtUYFL3yVyMyo5m/hKs08fugASi+F1Xlu
SITx/gmo4w6d21jw9quC7wm699Q3ClF6dFJ7CbufGNZGVMEHIS5zlskx8/CxYDff9jn/0D97AHvu
K2zeGmuQbTjpnVq5kQJm4NyCbCX8JoiEC51/0GioL6hrXCCi8guYBk2M3cNzow8JFIL7UATSnLqW
EPN+5OpB3ARdfwl3s8QYDnl6zFWGI77znEDJBqJc/NFHyMZG6602/aHRzZPPnnQArDAhP7CdtUr5
N9NunCu0XeiEMHS7fv2jFb/xoxLUY3lqmiAEvV7YVz3U9eCSzOtrDxlaVQP9e7hv8ZjK8uqMkZpu
hXT/c08rggTyXoHbFeMvQ3fmZhDTi/0DV7RqVDVLOGivXQv/0+7wSiw1KY3d0+ldVfqQqq1C3o2+
Yu3oFpCyUYr6yxhgwdfzOHEc79sZ3Y9mMPpezNF2OvygQJDzlWWa/wLvWhz0N8rPjxeGY3+UMB1R
ZBij6bfk+yxBaxIvpY/Qn227FnG9YI3XGUO2JKsCeheGZiuXmoEiHnkNyW14JEVsdLycnC4kJQYw
PHKxND8QDBOijc3ISNG3PGDjG+I1BHenAf39Dpg22ApFWwf+Y2C/FQIi+l2dxKCaAhevvZAgwtN/
JVS8ZH1sOp01SMBB074RcXNKE08zlizbaz7zDzPQPCV3zutPYrA6W6NS3qXs+kft5qAnx6Rrgkdy
48B2085ec8VqhUSTWmXB/mthzoDG7B/L/6FeULj6rnrSntQFtdqnodlfotO+VPHFgzUOKysM1cH7
sBAntcypkCdkB6KhR/WQVfYL8//zHHz8jjN1Ity80htNCCUyh9VtnvrKe+39NiHJvMt+A2uhTzyM
GswS9Rxw9UbChaHR7A0/FJ2NK0DTgiR7IdkC3b8Uw+5ELxIyPHKzHgKllgTog7Q6U0+Mb+Xr5U8n
oxNs7bMrlbeBmIe/SPogN0L8tDL0uVfTjjNDE1kTOqAL26jmcOOWAkr3F2tyhxc8NkHV/j6vHj8S
QP446SHsYGohBmdfAbJACkw2RxBs0MFb4+p/NiRZ9iuR00l0PL/NBFVpWScN51FGu4a+Iu6IAUoN
TeMmOnOEwTx5q1AUK4RT1+xE2f/GyzNyfs2b3gMgogGZPHeeRUVn7HPi0/BYafUB2bTjWGSpFGH3
CInei7BR11nVYmytkLrIJuJHO0Li3p3xOgPTYEPxjgx5pVHTui8DlMFVUYmOa3lVmdJuA61Vc2jA
vjnuC0v6au3Xvkj9CKAZIi1+2SO+wzLJo9SzTtkndbmsnhp4SCpMDn1v/ADYRvMtCfmgAvA01d1E
ng9/Gd+HIPRjNDir3ueVvdtafTEOt5qKHRbw4D5de2PoVaAvmYzE5/RiTBZXVVIu2QzLY0XBSK9e
Fhx85wtJoMOAJqI2kCf3dK6L6q7/oHj0XzCGYNcpiarnX66qcEgFpbLj/U/qFnQr3BCAh3/Hph2F
jArU5KzAI+PdUHQ1QQOYgAlXwzkf358xb2KWVzwqd8tqydIAhSYMo0xcjn4Ophgg7FwVAwXvtHVM
b9ABqCHAFAcAZhEYr8IFbLgiiD4RtB8z1YJ+AAk57mxVtDr8r3Ov/e+Nzbv9EZ3ch6hWjtsdmCIE
gFE7S/TFyn4VrfuYTegvhxl8xQOUnsOsKaL3bL9HrptfIEiZ9BPALfJtsdSlwX63qoOoRZV+43Wr
rdol3LAWoc4fdyt4xLf+cz54kKg2KBZu24P7PghM0hlLqqjzF2QbkJ10WyL9kj/DmIRNKPOYcKeE
40b7w2OXFhAyt+UCysBojKQxrY0fxpNDHNXTXiTMhFxBJErHk1SElWCTHuMzqN8cM6caPwC9baYG
9V4m/KPaafLHRDnt4irVZm48ZG8P8HRtTiUAdURBNgpwN5x3yqe99ryMlN45W1dCO2qMvbwuBuFX
j32WqcNE5pI7F+vqpl/Hq61pymFCuwOZkfHGHaIErd7pY3wgAL71kZzFOSlGdDWhJtyamBJ6+KSS
WGkHbdaYb4tkSmDdDLEvJDSaYcnmCu/XG7jDG6QdBJVGBarD6kdgvSrh95I7BXylBsZj29qknl6Z
ndH0PPpTrjizs4cBWHE5zoE99qMyuIi6bcNL+XQthoAHm2bfRaxv3vX2BOwBLvcG/vodN9+6glDM
LKmRLbqtSCLBsFgEO+s8xZSS7l9dihS4E7yZyqA4/v/VMk/DaXkkY0G9rqvOChD84E3RSv1vkzV7
upkGGfioJzhhLSU9xEOLHfE48yTUfR3zFhP9az7Nam8srcPJJdGd9SZr04NssDDe9SBCabvOjtYI
/WYrUoAeKp8hyKxA0i8/yPbPJIpTv1Q5UWJdDx0bFhW39bW9z658E1wq04brRlOqb5Z5kgV9RdGX
GVMxekWyIFUa9zgN/XHlTNb1CCkFfap606vF6wHShE5992duutplorwylJrs/g9q95bCCE5/dWjH
bildgE+KkH+cMBEplnUk1O0rc1FnJLmOH+IhGaOjonuBpOUOb91cIoV6HW56UpynSMpHA6Bo9IMX
HIkyN05ZKqfVTBZpeo2wSbu/O/ouoIYV4vptmGN446O4optLLesMMM14vjJR7eKEL9TMO4sbq9el
XqTyyhpvspOFFSAl3DGzlHSc/cdGsxWNbBpuSVGfePhIXQ19HyFFquA+HkkvkYIKRf1sBVt5GF4P
tSwk+nisFfeAnmJrKgEuSURcDg6SX5ZUFqJ3yNfguHb6po4Q/HT2Xjx6v8SfSGCkG0xc8GZqeBER
+LnsfssAmTFDW2NKbpxSTalacMtdxc1fzQAf2oNEQiwSbk2URNWJlAGThb3HHdDi9zjwVc+POwql
iYQassNoYQ9EjCDrUeYBaHvHgnAVmRQDcdLpMF2TBkZWxiFsip8znUpDWoBg5uh3fQWq7G2cj2En
k6myuCKffWx0A7ktVBKg3WZWOvIUwbYxoON+75hZ/Um9kZhdfHxyChtMwsZpCH9/czCrpwhS/VC5
pF9cVJ8w4kGvRMdtaklXaAp6PI762PDrSisVaPyiPYj4PfGAap7m/1d275Qr5aa25AwsWvWonZPv
yZ8Cx6fJ4MBve/0dvAxdDcUqnXfOGbL6VKz7FH+943kNWgcwCvFv2fyL/PtTnMsYH/gY9jKxNLAb
MfqO+3R0ST2K/q+q6lv5ExVhEVuBGVMXC4M+rSUAIw/UDciwqBuH+LgTp8SCWN3nImEYg5DuV8+g
auYHEeGGpw+DPeAA/1x2qM6C0bMHRFAqMH0DEGmkwxL8LI1/4dKwtnO+NXtC8h4TXJrmlJZ/KJMp
lJGwtfh2CnRAsjlADrN/eiQbsh4jEdaHMGBNdqnil82K6araHcqjLrZGqzyDSPuVZJWk2l8jc55E
5jHQBM1hz1jQjHcjP1bEGZJZPzMKh9eicedm1bDQevYd41vQXgy3figo/r2zOL1vP9fSNDDykbjK
W6tkmMeLwh0FShvbzISyFn1hQd5Ir3i9hduX+aoxrIHqIn9MZqrhTupoQwumLMZ012aRSTFRt/Jt
CMdgLz6af/7CkY90tt6MRVIl3LSoON73c6zJm2Nw+ghZ+5b1gACTL/pZBuzCuRqVbTDG7kFqVdIq
zFWqXHv8H7kE/QHkozvY03xKwIUilY4bPrOGl/SA2zWsJsB76qKpp8vyChaHdY/lwLl+zShMd6lY
OGgfnxH3YQewmJxvwsv14y0aG8yUAEYna4NXbNrH4ePQoj9p08RTDQT+0QkCiWTqTCYaOEHlBm1x
FJKCexJFfQSoBfRTAqVZnuZOenI3jdsnNny6JM0ZGIf1d6X/8nPHZUvlHyEGdBdGZ1bqBqdrvqWq
svjzKea0DgTyR5MlFKeuWAaljQi7jyBqaCGxZAj2k2ZDcDvnk2yHE4cafOCygyBJblAd2jU9rJOg
fejleDE3y1zaZA7zePqpNbfRQrmcqT0Vy/CMLSycm/0PkRdVhDZb9kEJYNIlbn79G0oJgAZqUf68
HzgE36Fsdtf6TKmfEkrzNabD06tVYGiqwC/b/9gC8Yjg1BfXha1XgHRoXlyve/UNv4AuPirsGOSz
A4KITwPWpQIfGLsHwM3ERMO58IpP3kIofTWYb+GY4KOjtGtSZHXj/7VJMhe4VMkiEL37wfx6jJYM
DIJjj2dY0WEDXDFObOC6n9HR3KXaTJ1A0JMsWogzqCKJ3BfW4yTiOoGgrxykXiTtq6Rv2zMom1Rx
bF1gyAt9IbxedSCAmwRFpFBKfOyTIuSNrjNiwcIXYtCA5+T3zYmjvFek0a7IW2FOdU4YOBb8LQUQ
2jUdiT9pdqnwaKbbhulda91397Exi4RcGi6VJtpO/78XAZkZa5Y4Efh6D/Qb4HFULIX0KbVaz8C2
vG/kXNL0K82GmsOkWIFP7ashEfnukBziXRaB8My4cAz/oWDlQEfUqUa4u80VRyeOFaXfMd7UtBuE
om2INkYKhrXzGEYE0cQ+9pKHbG9xpxUf+bU7w/cUu7BaaZlVf/nIKRKqdUCitJG7mN9NZt+pUcQt
SaUF6bwFEqcyiyGnj1QWc7Y0PpmSPlWHMCUnO96h6vn1qEGfCEleToQIy75OIJYwlPpIS+AOhAXD
T9fSv+is/0SLpE9Kj/kTx+v3by3RQuV0TtqypT46rPrfoC9SLPvkquj6NIWQ/VPg3V3KBJBsSN/p
An/C3UiXrOck8E4R4EoQBNTBIdQH2asMUZoNgHrRp5DcbrOvvSDtL3cTPMj5T0BOFSt41ndOksAt
VCAuViZjLw7c4i6OY8XrlNUyCZkBJXvdPadirY7NiVunLYNeRuHCzXm0ovUEFRqmnWpAZ+dXi/L0
zXtjjaDSYUlQpAq6+JLGgel+t+yyuYikwAo7to1JuDFPySE1OFXgMor1ClsiDR0oAnRzT1QAAg6V
KREsIG+M9EDaQh9gn2w4LedPTYYQkI2B7P8NUdBUyx4dvPjtwZLJCu24R6Djed7NYngXxMDPF043
casYQfwf2MhMUIYi/FshfM5bWBL42aGGf9WzBsNksWYa5kZWb6wuqwPgzOI+2QQBTaYC8bSECmIP
cPLZ0eqRMZxFgVrvRUJC6/x44sd8ikLcfwUU5edfTTTYb1gds053z1ZtfQUqi5MhUf8u3kDrD8Mc
0ePl/IUAWell2OHt+qN6jYF++/grlzuW6+iRR51PCWqBL8WFghc0u24qdOogf2GEfKdiB1Z8x7FA
MNrIWf8lhMLSOprQJtjlX0fxpt+7kQYgX9lV+0wiaY+8+VSOhcdVqwgBaLlTaZPZfNr0R4TS1B0t
jCNTYA2qG8a9LoTQ7lGF5TXXSxZKezYJ9TOwT/SK45thTBaicd4weT0ZW2f8f8Q7DMCLbN2z0/qJ
ubleksuC2kRrAeA46KA3lq6UpdnBT26bHEl/5iGF3Kcq5Ez4Veswn5giRtyDC+i6ppQchryywuUT
ClFxRnFiTM+XmXdr5ul61Dusg+dw1VLmmZ/Z4dVTDmGy3X8f9VcFbAdIlGEjc/+C1nS7WSnTkMQ0
NCYC/4zwwTNLmIto5/apFuCNS2eKlRP9W0iu9QEdsYzlzUr/suIj9NMOUvD6SlGghTsnPVIvdzQG
Icrq2DMgMvbc+PnfTOKmmGYcO/FQJuyNhkfDbtOWGfCAFQ1/fJ9mIUMRln6yoC8C81+SsXyIz+L3
w3qUb09p+4qIBCwEK9DTESsWJm/4iQbIUe/CV7rmy226xobFMaTuuMs7pEphYowHNSp5Bc4WPdGI
nc8pBU4klAWe8MeBVZutiAl1qTiFLM5y5/sxEpHe33EFnje4u9l+lfcPAMojlTfCDnApVWSJhE15
qzgXewdUQK6dVwLlUKRM+HPofYYcIEOuRMjJYLtIKZY+hFrFPzAT4IYt/+OsSi7WMsTQBCsMgI+r
zg6QupxF8lzCfWSjmq7T1q9jS8GSNYkbRopU3RpMLxu8xwlyrNuuFJCMKktB6QUZZpNZKqC1Lpl+
cWh0VFNj7lqgzYzjZEsQI1Gpsmoo56MnoDWjpNsl1Ql+gvMnbdyqw3SIeCQLJs8S/tTtiHCp8slK
g4VM+WkGxq8iP/vbv6wPGDv0F2ATio6EcHfhJeC6QX8m+OC2jGMZfgKZ+WBokLjPaEuVpNYE7Xaw
JnhRUbwv3mqW+3Rfg+bTPys5DVyWnkETcbooIPEEGisEMdL5M12YHdk73ooHwqpczlc1s3WgS03u
wRlqki/EIoI2OnbiEVDs0LP+pqzb4asqZ/L21M0XtjC/j4rS/C6nbmkRgv29s6cE+FMSz/GhVIfZ
uBJ3wBPIU7c/XnYmI2u4QmYtINmdD+Qx/aSe+ytDXR0OyhTLncbaFxu9+zUaq5Y5B5w0LTjfAFe6
L4bp7JcwidWjUDli4XyHCI2K7AgAhkWCYevMrT2ZrAtsvjpEdASZ34QEtdEGTLw27GLbteMd/cZO
FVMNuEOSErpMU2LW6I47fgM+8+3DoHvhScAZS3cfaXjfXggGg33azosTi4CXkkU3HoeYh3vhVuZw
OHt1wrCt8a39AtbI36uw7KVeXQUD0y557lmLTS8Ld8kjzRo75GEtb8A+9xaxaRvtTvG0/50NadTW
uoFs/6s3KMNYzwLgLE3R86TdhSS2GjSxOzWvfp+GDMi8FFqp7qiNirEHc4jZg5LL+nCrFM+tWk/3
7eJQG27+l29K7XvOH0JRbiI9DnYCBIR00i7XumCgLdtIoPxL9J63XiFPvOCeBq5ch1y143uKJ0BC
/MZe7hFffqrC1AjFiFhBKvg4leHuSzM5KkunvtwFRNCUnao4luY1mX3ugQOfNsybG8m4mWFIUBmu
nNIXAynznladyfmsOMHZTDncgvhzwz/sd06XQHu/CGY5qCpzDcRKA0A7xju32hjL4jC1Zajk5tj5
idz0W3UFaq1UwgVycEooM89iWftIUhn9t+uZmE40deL0gE7me9Y4XTGo+4x8G+DfZUYCFCqhzXod
cqrRAAMXlFAnYjmy2wuGdwJiL0usofR9hCbEgxYpNu4QUh7S9Axy2kWKuZBRoNiMWL8nb+e6oy93
wFwW5oqrCMHpq4EK5V1RUR17ji54exH5Wl/1tgmSyYpfC3TLDfupT8P4RP+gJjtv07UYgZFCefWl
VsTCLbCaWF3c7gPkWaTi6dFitV7BUcKE03Q/7FGsLXzswLduyY4Pe/P8RkerJp4ZEkykrsXFJ0rd
nXNaJ1lI7UgY5SVpKChsjk8ttB8mCW/GVrn29cS9YoZ4YsqRef90eMk5C0ZuzOzowMFlQMmjTPhN
Y64pz/Sxw3PMOp64DP9NuUdKEMw6nvKG8wqNZ+wFqvZlXTo0itiYy4FuJcrB65H0RwuiMmKnU9DT
Aeudq9SatcMuOO0sUQws02pAjrzqEITqt4ftS43mpVgtIAc01CPIZ4a1DorRCt8PaeREwuGvlB8L
d8w22f93yVJk+EwE+78A7Ntod3pADtl5KTrSLdrKDwmExxqAdJ0+POuUSBGV93j/061XIa37Q5Fg
icg6O+bvENuKsWXzrR+bYnze8chB6p/5ins40VZSQ4LFKXaa2S6I400qav+Ua11kYfq1KK2s9OKn
DbUFoiHAptBCZ4XjR+oCmzod65Sb9fR9WJu1esectSPs8TN9Tu/0O+STgYHrk1gfPEA9lvPK2RxU
Yc9OJjotj0f/dEJ7o1CmxWMhBdxsufziwSGbr2lj5aDXOCkN7vgce5gPekLWn1Kl+IPKUnAIIx1I
f3Iq7YehpAptu5SzIjpgldp4aCDMPw95ujNKbNRdwDsPVkLp7tJ/Sg3/ql4odCEK1OG3JWnnX2cr
Wv/7/B57/UWTFnF+LzK7WRyAnjIAk3ak0WvLNTiy+zuAkV/BNBm8z1v3fv3JAdcXhG4nfMSCZB98
9O/bIsghRrJYlYh6NNO4TT8hN8VFZvouLuAiIau9CuLbjW+5ma2LIkDmBUjV5UMu+d+biEO0EcBt
vOuPU9z+RIM3QKdktlgT3EvUEW92C9FKCfAzpOyFjgtHU201a+Gl9DZuRI43yT7h8RwH9DD+fn+A
aTo5VGK1zbcrVEVllTb9k15c+jIKFtWGFGqzgb5ryem782AvOdzbzDAGMcwvGBWyGlQD49W8WTd0
hiu8w05NPju9qH6X0Iglb7wdBN9jbk81ZMqiBoX/lfKm+0/qDvgcyZ+zeb8N1Olv1/QMt6nIp8M6
LV9Cj06TsjqotP4Ob4ZsGDOYJdMZfRevQX09IzVNWkq57zC1beGAdWC5MXAXss3BEQgiZtrJGDON
fJjF51f8QCoySiWvIjttE2dfvbjjS3KbjkQ2Gc1xUkMCelKLevVVIvEi0QX83+sGNd4HFNpOt7Uj
CAEV6cF+0oS7Olms4RnhjbNDSboHemdiVwJFJbQiVH5phnvB8EZHDg9V5bNS6ErJHhOL4oVGWmb6
gYTalCz4BXu6uiQ1yoF+MeH6arEvjXE3BpsEMgy/Za9CI+vyyk65RM45i77zvVQ+ACyw4XMSeKnG
m4FZrLqjdlyg6BUVlqEsp9w52k543Y59hQOJRV340g4iM2BfjeeXesUVgDizGNmQ74Sb8DZfkJra
9qpr7mEDvW/bicNxxsOUGNZnrdC9z+RUAqj5faQNjWmuYf6BbapIjFLoqIPslYjDTpNww5o2t33A
6QlhJLfSJHJ9Qkc/Jiqnp4Ym7AAU0ySrLO9S32kb9V69BiQvkfz+QscctWiowG3uqeIEvH2sQZPe
AjJzvOUv57Cjgg/Ku6JGbKgynyFPZ/ryOBhhk4IbGLZ5Du0RsfVHFXNh0awOYTGV85r95euHMkHm
cGoLvrom1F001GuOq6m0gYG/49c3pYJ5cl/jy1AORSRqS7/hiPbjEPgK/Ctsxh1e32+iKgBuydL3
8bV35lFSrUN6QKPkryOuOMYuliezR46TZf4cYlPcTw3Q+MjYkQ9uhKgRtvRMk9zw1OqlxjcuhhsW
RTlgZjU6R7UazkLsxH5CdMJNrVHzOSKxSYROoIXh9ox0CiFRNrY19idOtzFCtz/+EeZ+0mc4Epdr
08T8400DenEvkJIYZiOKZcvW1Vyow+1rpoJVDUcZHbyAfW16UcfP5ciUWWHbWdoxd3q6EE6nJqHF
XRwuEZfFhlxEGNV8qYJOGkfQC+DEjEbOSw7vwwu3JIKgXY+nxByRrO48WRL3U9c/ztBo66i0hsQk
eySGkzr7Vyu+rRKL/IDRBnsMYiZyF9pTt0Tla9Pr/SmcEse2vGlhHAkfSbTmdSS1M0xYJV0eSpcC
usFi2WZlPEyndOlvlEUQfh4SBr+dh/Itbuo5MURGak+nGokI0sDeJGhUDeV2TgophZZkC6qEzYyT
KO7NbmYDEGBPq4eosRKznqjir+Q6flQXAUwi+N6C5CbCdJ8qg7WUiavQyUW0TEh3vTJumXILvFNP
kZZ92LccxXLNRipYz7mLRmk95EyzH6oKPhX71Wq7s9gA7Qsk4Poga+vTuQQ3AtUMwhW/xPrhnObu
lhzuXMLguyQmX/gnxVX+n+w6FnS9zNBH6qg9XnRtOR3VE8z8I80Lv9dPplJHfzRfqFmexUWf082/
L+Is6pybfnUzlfNZR5K/3gA8HQRD4k3OVyl+g7+KxZPaSYq1Nk+6nX7U1E0+BKJoeTecJijJ9+ET
XcznnWIq06t7Zt/OnkxosYQAc2WwpWoAQ8fJm5rAwMck7ob5a5qwBvgOS9SI/j3tc5FMUPo3qegu
VPLddWJteDXeNHk592KhsF0LPV2EGHJS8A8qu4z/yg2IRTj8rwWQLg1zq+ORA6M3BQxQxw7TS92Q
f5jZjJpXenmWyt944quMQXT+eUsp2AWBk7jxpV5V9qMD3BD0eHwaXxQXwhrVUVUvXKLDakAMcxio
klTL0PoyaYEOptQj4f7iY8Sw1/pqqhTo1Hr8ugOs+L4/ZfXLuhgwMdsrZDgrO5vd70TxRk/lm//X
RSaUfsTTqwsV4R4PK9jFsDN54AHrwwStIr1sm5ecjSqgHI56pB4BQTQMP5djhPVFLaxR4VSoL2On
IQa8QkATWjKKT+m95wdPZW4e+fz48qfCBeQiPiK2YoLUzOFufqQFOJE1D43HYKbppvf5gLWf7OJM
OApCEmFrwUuCN0BDtwd3/wKbRgXC5/9eglpWzpAz+eJ45ahq4t5wl3EyrCvt5TWTzVd2TaRk1dqz
TqdIiFrxYs26Afs7rNK1mibJAp6DLWZF9ENItcAALVN9U9mLrDBCNgI7NH2GzV2t4RwtFQ4BCfDn
8/CucCdO6PYebLHmIxRX2v/1lMNe1qNWrAkidLHTH3MuhS04NJCbEX7oW/feNFWU4jueAesTLdxZ
Qy6Km9v1RNtBWpiHqAMOz0AtUgcEUV/+GiLqpW0NFFqiRC0KDPr2b7tXCtJEFubbTHKitVF2dnl7
LnGdXiWVgv+XPlaEp7FdUxWDvKnHkl6dtxMvy7WUTUjdTliU9iFbLB1CMmEOUakTmpBBI0MPYKHs
pHku3Bh4BClx+93MsoVHzzJEulHlZAKkfN0SuOmhX9S9ThXE3xZowhhDLHM/T7eNdy1l+zXUS2m7
rC7m6MwfrDqoDp2lAc1tv42s9tcdAQb8bsatQJ1Kk10DJ3A3DxdU6R58Juqsrbp0uoTecEfesulJ
m3OxIuxgalJDP5hvmuYjYeGf0gatfxy1Lhn/7NXLDmeuF/y6vx3N1ZMs0/uH6Yra99Ji02GVERI5
V0PyvyJFYOjRZ9JPLMjHan0+Ift9y3g8zPJ2CJDLCpwabAfwE6Fgrh+RZP/qiaOvg24QPVl9euEN
p5Ynzve+mMqPg503QLJXV2MmnqdGpI0kdZe9h3WJwAtu4RZaiJfwZl+1hKIQwp67q//XZMuC2WTc
qJcm0QEp94cfieGPa/wZNDCf3ddxo1UKyikyHANHnqtLN2s+xnDnZNdTEOSvJlpSrqtipZ6Tmh39
Qkf9tz+M/ioU3/okCHvtsREk6UVbvLIJTnAMVW0OuS7HIvk6+wrWPalGWVJwmP//ylzQ3kArxP+h
MAvOL70j+XoHZj6il6Q+rdR7l3M3xXMoHrFCx4EEqkJSk/xGgNjfLIgiKz5o+4G4EJR0v7QPBjWc
L/yB1ysTrqtc3Pmp9wrhtn4Z0mMPGOpVOaQ+sBJ94GZByzzHpLbMr++QIv0Hz9TDnTFQiQrk5Gll
JU5dwoWg7gBNCGxCK5p3gf+mIyIE5C+2C76iC4ea3yCxug6nNwwErwz+3Z8CRM2WbX3wOJ/quLCy
9i8dkDiQatubmzVsCUm0ItnDRCAcKid8T7SkMleLjMvpEp4v6GDtQLp1WOKdkSiLhBP8h7+B5fJd
USZzfOe6NJTBU/KdUOt8L/F5hwtAHPH6AdlWr+N4QG1q5cLyPi5c1G7fpyF3wZckIwkYn4s9XMIU
1D7yLSQw6ZTiN7Q9QQ84TdCvy6tVL773gCN5PLPy5uCvPAqJce0AWfAqu/bp8+qpK4bU6tDaqPPd
x8TGsYsX5HRGsAS6BZFp7XkH4D0wyaq+oepFYzjs6sNRkvggCh7UTgggVr4GXvQAWzS+XmTwKqK2
8KMxNjIZ/JHIGBG1i6MrFZLlWR7/EVHHfOIGWYy+bvUNpvswtRQVSM3SL3Ie60Tnhy3Sp5JR7iCV
mJR45vStIWxicDaeuKRYAoEOCzQkbK+kembuGEpt4RIhb32pYolGwA9pgrNGBwmqpyJ4mmQhqH9g
sISDAK8F6UNKSMaQbjnmr31VDFUV/zZ1s1vajFCwX8UAy/UBPumm1zRi11Mhy57q4FgDDQAoda46
FuVCmND2vq0ZdDuP4N4u6og+XJcB7/5NxZbxDDV0audIc+pDLimV0neEF5E8puh7CFjRUcu8GbJl
9B5pMhynrnK85KsNkFttelRnJrAxioz/CbGpO+xckVAIOdValFytEC/5gESyxqTlO0YMf1prfEx4
2YgUsIme0A6mMiCWhoRh5xbs3n2c1zfUKkcYWAt01oPA9sOgeIP2IoUbHqt9cKYXpLYF9Xp6CxNS
tXIsslz8AMkSmvUP0bTy8XZ1o5Im+rZ3kOPL4JsihIN7J3N9JgAdJlQuigLrsVwcQqELOuXgwfZ1
r3+nrqd96mla9FK1XrkDUgD7C17nZZQQc6uOW8IrnBogNkMlZDyP9WvSVZoN4SQv/I0jGDNhkk2C
vJ9rNme6lfkYb/10f+Jhz1m91LWNS7CSTlNTJMKdwX99iKrhfSid6iGWSEQS9TOqfKBtWdTD2Eg2
bvph7zOrjw+qBvo0LmltOKg28EdiMrFnTsW14M+CUOqL3wSxEMdz30J7ZAUxOYNFKxSHx4+jYcu4
XrDeby+vxoTTS9tfhDiqAKnxHcjjaKfBZ4/WCVkUJT2u4SPyOzvo8Orpvv2vNQoIQ50478tKgsu0
OUlgdlTjHwKH+M/eSBLd+sVcEzPXmoPAm/J/iv4V0DmCZ5WL3rGMNeKYkSMIhF4zUQRlIJtZNghf
x4NgI8bS9MWx7w/ryrlJg6fYAFy2IQ2iKHdbpJK74D0H4UEYOaPJRcvaQYRHfYUSbmALm1GUvYA3
w3eDupLWimNHgOEGccPd03GFFG2o4NXFszdVVYwuN4/MfcwRN0VF6X4HT8NuQhNwiPWmHKL2xXnY
mRP6cATPJa2mJ5zN+1zcye2fHmLj5darrsnukOrw5ayBQLrRDSNGYumI1HRR0Vca4FgGx0bp3Xpg
Nx0Rvob27DHJa51rFVTpHq8kGQNQeUAb0jRggQ4sZ7+BkpGT2ymbU+RbZomKygbv+Iynr6S8+zL+
F6BLd/CGw50Ff8M1Mh7buo+aftBL4p/5Yb6a7kRrGYoUuijwzRcXvMQ6xs7RYC0jRI7clhCEDXLf
xQkUOAQ5RfUXRzkrCrCQmdEMiB5NtA9ciZ+VXaEYG/tyOMK9uErq7RAC5MPkXxEo8rOwMrkAATG9
MoW5uIf5wiw+9QzqaHifjA175iZ+0MMeTtXN2KBEMFbw7tlMh/SfuCXhvFAEmt6SUdO7tFHVPx6q
ToCb3sM5F4qacRPjTpWpBXS33RYqmvW5oY0TMESCMDsYOKentcHfbeUKLPl/YqMO9lKeD7O6chSr
a9RdjjHWOTTb4idJd88WU5LdlYzOoBDbLtSoHmNWOISzrKNSS64LeKqgLfk5PfHxMWfjAptEil+N
/KpUPCQ+M1tqJT7tLSNb5F3xVsfMFRxnz7C/Y2yVoFx7fnTB5GLDfrFEkg6szEqQLQWam6jDnsv0
iGDSOp9RavaUCLdlOyHxfTnfiV4lEGe2yVSgIjpZNt/AhoR82p1HWJxZvNfQl9Kq0j3lLZsjSqJ0
d4gqm5fdljMVMko92lrxiq/9mOn3AtkirK8zmW3LTGPFrkiZtnEL2AdC2g2VD9iTNNVDhvDnlrFR
7QQ3Vt8fa6bQIXSbD+P6OgpxaiY6JTLEmzR6UD0ncUyPoqCBPrpekD5nLgN+AHQ7S4DpGDnC+TlH
gEerXixV6fMGFa45rrXq5lCh6o2+nylEBO3dLQtI8YUvIZod6snYNzseNSG/rsYHYWJOSH4EC6+K
E1GCjCUR63mHjI73jOvDl5PdqAfVaWkIIH89DJm2POK0O+LgyB5hMoMhPyiN8tCRy5puxq3OES62
8x1wKkb+7uWajEEc2hvtqPQmeM9ZCN1IzhvnX8InZrayQwzthwUYRiyrW7oAIUA7ZPkiKCb79JVm
3TxL+Sbd0hHeVvE+DmVPFhDHI5DFgqKY9cPZgtAKZva2ngMz0lAe9PebiinwXwXVlt4a0eaTHRux
qAGgGAl1JZCtHliQZob5TUenTH0xyhYpFB44xDVDBdh2PbCl9fwR/Q7zHfYQ5Fa69+6eg9Bhb1FE
nFwxko6b5jn6NTfUsF3u69Fm7lgcNS1mzRdhLFApQxIN77sm6O0DS2aSBbLAp7LlKLsc0ibuE8Z5
iOOhCB3ljsnpWKs0Kai3k7AdQMgcMlVuVH6lJaHWsHgqVgOPwye39SaT2jl5W4RJmdSinEb2cJ+d
81Lb9IRYeuJUGdDVr4o7IWYoNZc1UCIZ2hpG9fDnX/CrXab4ggSMK7xzXR5GUE4zXDQKZhrEsdzy
eRm2hUmMF6tw3u1JCPR0QddhKcMmb6b/lLUbtQqIPAJqVXlp2sgejQpC+UUhe1HoLblsVOxByeEB
YQK4iK7AvjL0rb+QTtXXCgctWrRcyYNdiyRQM0gTwqW14umv+oTHwMhuQz0ryyZ3rplmQOayfXQE
gEEbr8iXE+LzKd/IrO/pZt1m+WAeJijpska9TIVByjq9mSTIkbL4LCVKAou9KHogJVfFXeQzfbw/
1Z5Fg90VdySKqwPyAtZCZ0h9aqAVvMYQ/D6rQkgcGLPWjkv6GVzRXfUqgq/YUFNUvyZKVaeOeyTr
unkh5P9WydV3vFGSybPgm62yBiO14x6kseiDDqC4ypHtdx3/hzWmgKBlrQdhOWr1bdKKPLr9Dxdw
qEmk7cA6tCT72Fa5d0R2PXBOFKOzvsxqYAoAJ++7RyN9SdOeRFlwwj+/7Ge1nHqknOT4B+ZHO9aU
vobLVXfq+68H77SHzDavAS8r8UldwrPyjn9/8Lt7sISVQxQFH/R/k+45Rpbt/LUEA0jZxZ+V1Cek
l98hqB1Qspa0+d88aXOpz+nqwEUjD9TowGq2OnCoahYgmog1sK0ppyAsAfdGsMtN+3Vc7IReQn1B
chJl9of3GBtiTOJ6UzUKOTSuI0NNxxTvMkvW7olvaSqhCsgXJS4fHVmhHDqBPxEqg3pdDVAGc2GC
swoUlDsUlA/xWnWuEB5PB+dNwMiU+6meLgXE5MyAncyfxToC7AQXe8bVFAjYrobQdoFpU81Sn5Z9
5o9MOmCLq+n/KURUd9G2uIYgywHGxv7oNMpTgzvfRIa6IV2kF67kxFpX5MH+68uQMCtXsiIFzGX3
sPlArrf9jCl84SJ+B/0LY7zBw8wubzCVQeb+lqU2yQgVyTCBFhUzbGDT4tlwP2arl2RI/QqDgyvP
SyMOhggmXCncI8RJGGWBhq0fbChjsgz9pAln3OjJ9ByWUuBXZSkmcPy/p1qYae1NJwoEHzB2+ivc
qmE2OLu+uoejFAG1rCiQaLUEVdnqzhUJchawgl7JclM+J/0LzgXyOk3Z+XF90oC0MvEMVw8J8YGH
ybxsJZJGhIYCWhMeGVBQQ5QHM457MDkwkhcpuicy6xlbTGMdIRtRAanypKvDzxFfsOhhUksI/sjr
2P0SihccnlXTUreoEC+baU7NZjic/guOi3sGQvGeJsi3eCNrOtn0tlRfn9BGxzYKHc1HElkQSCrE
5HkE1dEhtHx1mVynUnyBHYjtqPN4L3+6jvA/3WfmWA4edbIRYP7LrV3WwLY7Mql6wHFNk3n7ILt4
m0RMsmpZ7vLl6jtEwgkhCqicRM1YKJm6CKkDaNNk7KEKRNgZeq0KOMvVUzkJ2tWpLu0v4Wq3uOdE
h107araPAgb5qHCOjChK8Mlo9/lzNJhFgnCl8la2EcuYqrC5JnmZHXX1KRUlB2Nx2dU/iIaHIhIw
nUbszTG9WnH/HdcC05AR5ntZu2fm67cGcYvlSFiGJKJ/YsgdnyVACxmVkA8BvopYPjz9jbMYQm4O
T1PiBFrX0mEK4wSoz9UlFzM4LMafzw0ry2MMsELCdFFTD0NsvCmTI3vYaqt8TNxUiB4894+w+lR/
qwe1VrOEeY97wkECnqQzDWnfwUJ2Fp0ZXy3EhapC41neIVha10xu/6JZKnbbwE6s2ex9geJvL0qg
iWKMgekOrZf1TaCiCtvkpqWgzomlD93h5rfx/XbMP7QHUY6VvUUyaj6q+I9xqokuscN3GmqFtEOi
cazfiZpZ7MU0PFchVR701qSAa5s0ujJvNmyeo2o7j6DKfNlYQAtxT7CjZD6ACeiJOrqHo3NdeP6R
dISLXSfqhClBPmEJY2ND0nYsxEx6inVDW49hgF7IZozA+QqAUHe6SinWomwZhXvrjjkbuqYHJtEQ
BNGUjM8YzxQ6syy2eg3PAFFpkJOpVdgUlIYF3gJGnacQ4Hsu0Vj5Ukm7wnsc18t91Te0MIx1rVwU
1HDmAjB2n0nK3ZBOezFp8UF9slQGM7+Zl8dCuqiFY6L6Hk+FohEYt29rNehjkfux8WwHBML1PyLs
zHT5LPGcGt4FLq00NuwyESKrNOS3dzoqGDjlVkutIKBsPH5L/MbrtlVpkovhpTrLmsePOMqYeS33
EtyXyl7bWLGFLFvPuZffDrCX1NsoGmXmH8ijzt77QAlu+ra81sygxfXbkC5OwEceSgWQY678hJhx
MMiKzuWb4DmYcUqwMD8lFu/36lgSb59Wm6WzhGKc2VZgfl7bNjiz1Hc1OILuvjI0PgLorqIdPGd7
d6IVBqq579CkOMiIf0Xq4msM5B8BkH+WhP63eMb4y85sRR8092rWcbUArUV0rPvFg5SNov0+iYyd
5e/0LFEHjcC7+ddnmMVVOpUJD/fgx+1eoOqFZ4nw3bDHl3WYSS0r0bStf8ejoZzL9oSe5CI/tCJg
zvBLWTioFlTTDBUWGR2qIAhbqgpockNH4kQkODvYIZrxhsvg6z/X5uNCZnhuNJPYZzfvELCLKiq0
y/G/YJ5OzhN0NCN3rrGUNBzhftzczl5d8Gh8wLPQKBQxJQX6nG0nk+BZ0DyIwyZ1Nf0up+bNZ0mL
vRBzbBCa6+1meZfS+e/M7UYDP2kXRbRpNCuUk9EYTHSQgFD4vFzjQ/8a7tcB3Cn93ZsCovG/mCjF
ivu3XrRYzwgNeimEJN9fEkVT8nDu9KnG//Ct8EUNVEmD6dwgz7i+QInKDij5FWC861S0G3rIg1ul
aVupn4MWRw49ADPH1nPHBMK5Qqvk3xuSZVWGnSCwi4Ovap6m0lnCI9n+76aLonNHR7cgGK1YNYD6
s8mCqJs2kuITUCJZrKj4wzC0+VeeEYxvzh3wLVAWiFLDMHhYMCAxhS0xiB8858livx/A9iYgY0+M
lN50vTVa912yXCLX7JPWwcPBBPmaKrKd9QuJUqAJV7p9od/C+gEHWfl9p6CnkBa+APXPYTTPeSYp
rnIiCJFQLP4R+Bt0Sr56AGNVmUSfPMGr+JnjO5ZVNyiA1U6CpDWmQR2SrVPs0qWmqupvXNHqeNVV
hbY7vs3wzaA1t8Rc36jMT9HgETQiwWTzpMDzv2GRu2hmbS3NNZ59Kou9S4mobaNMPlk45kaFcQcl
+nn15LMtfdUXzNikCZXJjQTwtD9GqGIAz+K2mYhlz6T/yDDhJVzYcTnwyMpEi1ktHRXFzyIQVqqv
M0F50vEXWv1++aRN/ddpKP1G+Xqhmxi9PDx7VG84Urw3EpiQgTYfXffv8KcDj+rbMDkMFK26ARfa
2egMiwWBtphsMjnNZ28YJBIFZ6aNqNyadrj1CSe3IclUjROSoV7eLnUg2cNLXyEwWT163Gx+E4bc
8EMjW/LazCtsbVLjDNe2lR+PMU9gjiMtw9AtXYX7RdRzPuyGxGG4ngbAPbRIVrx7QzqG2DXxKQWj
VlNf8Q5JxzZ8rndkMI9GsFyQaOCfKoVEVzSAp5Qn9C5mAg1uMmBNUgecevWRD912Cu4nTeKnM3Bm
B9MkhrTwI3tjnAZiOwyEkr/lcPkM2hsojmvrRBSSg7/iCW7bO6Pv5WbfLnhCaQ0MjbwvW71DPyLy
aJ27rE0Zr8KTNThuYc1yTcP/QxcAOHytawcPKS22Sv/02fZ6xviL6Vwrl40JXVxzCb5bOGSyl4Hh
zLujEkDtoPRQCCBoZnZsPkjv5nt/At5IVneniQJGPlMBH3GiamL7/goTUMj0MpHcYu/QJpu3VwWY
Bpl2rHaZAkDx0KLr/lAKMO9Lb56rjjp2zXwizOrqy5kx/XLU2peM2wH5ndzRnEiBfeJJzlIerBHT
x9m2vz1IxQHgS/CZlyPFMYpIiDndeii55SnqkM9L2Ciso+6twIVjVGyECI8BxxY9N8ONpedVwt6g
vtuGc1eGtXnEDiVOXiahnUyicssDj3tyOiMhA/Eq0hvrBgaw1KS6MCo9LjA6SgjPM0gv+zPK6GZ2
eL6Ic89rse8UfQnOigYMxeDNHDw78E8xOsf0phYNzh0Bsozsv15I2yDqPxRwbed9CxSFLwUujLmO
575CsScOTYwTsx2J454BBSz5/Gevz4b9fE6ZfQ2teKG3UfIAlKDECmcdYmy6LHlw0SlqwETsiubo
Pyif7sFhNYJVNLjS5mxnI4dm6Xt2iJ5VC3AriWSA050twhlLl6VPQFhZ67AIlDawBR5e53cBwWtW
EyX7wlHWr0aud8V4NBPmmVc1U9VgwP+4Q/wi7cPfQdnpRhSAti3WHvUSIrN92jCRP3R4mZPeJF1X
ie2xc/ZM36j7zrKhYx93gXjg+BMJwmJKMNl7qWwRDgM+agGGGVQKT775+sruBLRXk7wC1PcdGNkg
yYgzhpQYZz0MBZiTi7XdZNbKrV8DSb24q0RJWdeWos0Zp9qVHlAoaIqXM9kQI/D45M+K8d3XPanp
tt3gWwrVgqIfSX/abn4QpDcI1jfC5pFwXz+8T5Zc0s56262FGq0DH4sw1yjAVKj9q7vSiDsgWEmx
b2XtVseW8ZtZHp09SpVQ1TngB8LC/YV2S9BET6iz3lOK/rZSZwwLtXCkm2Vn9a3IL7qwbAmZr9fN
y5+vr5+RMJnzvnZWnu5zC5h6pudJZKz24QoYYIq4quAnKoDQBMqU4NKcpqavyYAIHxG/oFU5AS1X
Jc4qFoSb5TT+bCkuhsyHbprirJxbhgkkYcSCXZQXRCKbX38aYs3iZVbsN9WMukrvCt8HWRgxQbb4
28C7okkJKP1+yr3nag9rTbaIgZiK/jFvPP9ygndCRyrCU/szJTbEFfFBWxqywnHPkICNizxmFfXS
GJIcDpsMyGoGS8aokG0qCt3xklktLKJtLVyJn5eQhnIMbfo6XNr6hv7F8reHGAhcdM7yYcvU79qx
CeHTJBCaNYWM2IGMsYdm9xsK3C5CYFDChJF805C9aCGPd4vwqVH+xPzyN7Be8tAsL75wNQ7jXbR4
GTqjN+KA1F/ivi6W7d/mNmxpwPm5lYS7xDWv1PMz7vhJx0fH3yoCf0EXEJeV8arkYS/aulDYtTMM
oP1JcWyUhP7ezU7QlQL5xnUY8t67M9nM+wqpSkj7j+XkFaR2TAf06v3DHJ8O9GQzDHcWFNmO2urz
pR/cp/RlpQstyjz3qyh6O8vIYEvuUQv/UZhKqavolxPI73+9JhKjPxBBUTIBuUi60d5hNa34kECK
+5ebitbb5jFYO5GsTAO594e8fpuuDRf/Io9XPucPQP9fSt5eVsiR15qMXdUmJdE97O565vv2doGp
ZMpVpbxrpavB0K1bHv3+g7O/+H+6qpVtLvrLwOAEtM4kuzxEHrg4FP8SBDy0Z571JO0Ly7yPI40W
XezR4Fgt1x4v23SMz2XoAGb03FbvPBYeGZbtYyeTsVAm9BesQ2Om8zDGZo1e6HnbItI+ALIsvr8t
UUowg3zSK1FFDUKWLDIZXsiq2LRatGXJk6xFooXYH1M46ZZ13zljWBi19AADXA2cyXWQbaJN5KqN
7eYYdXnmgKC4RtqcGCKr6aRYn0OTuPtY18IA5pr3/eNwLrgsxWI8P8Ot5G4Fhw4bIw71fV0OPEOF
Smg1jjGQvTX1VpfrVGcP1uoIsCvCXWAC9jgjK5sphg8BGnpEV6b0ypSwV04TwpjLIoB4gHvbcDc3
LDWZWzM4cwyo8qJYeBOlUlpe2kMoYpJIgZD1F9Zhs5XKAA3+85WiUSkq5OhsNGNNi+avLBPvLngr
J2rM9oQXvX9FaiRtzYe8L5+5JETwZTZPEFDFQ+uaZbNlNB5Jpn2zQQ5Ez5omG+SeNvlwI/UFu/9/
0G9qUjdd0dVrlIwoiIGipt1GG/+D2blm/dHhPeA+VSr1qgAnM62iBNv5xPfTC4ynxL1pXkHUw1f5
TGyJdTa/v1hpm00bGL3yYC8zUAwxw79hKGuRQJmdeQjcR46Wd4XLcF25CZG5Kn9eAOhrpLyojpN/
h7EOJb2Aov/KWd0UAWsuvfqulhXppLTnej81f15ye2wJIDa5zxPOEuL0B+7DF2yHn6IjnT+b5Oae
nueC89DyHfiZjkNSVrGw7pXITQAZtRaQSiEXfKk0FlByHw1Kd7KnQMpvZsSKUgOBB6ehoXa3AtqN
qnIkVxQQJvdZPI5+MJe1HF2MxrKXE9hcL56GKxleyQsykwzNnUJTe3Wkncg0gGh0kvrKzBJ9e1DC
6wcskdjCtXmRI1CdLSL0VttPx2n07NJL8HQAVmOO4W8jI+1XnyCgvx/VQh8MKwx5u3tBqNhoMEnV
jmL9WLvjri5Mnzxaa6q+vOVP60OuSqAxrWDnBp7d05YpfQbGbKLpTUvmvQHi4UR9hIYjWVbV05ye
urxP8eXQ6LyW1smiE6AGyfFzgH3bOhfZcC5QBwI2l9yrX51Aszehn5//pla4ngxzFM4mURhIpaFY
y4LX+4NQzJCKVexaPPgxuHEMJ3XGH3Nv0zYN8LmK4UY3i3oatOeWBc3r/tGssRzx4g9MvA5bC13F
i9dKhCgWGylHH4ruzje9KmMcLEf+hs0A38/3W6IgM0u3za0k5hpL/pQYns3cIp5FI3a+Y403+K3W
1kIn8TqiDJ9Fpf5HhqSy/tXwAxueAuWbq+TECoLirGV8io7u/VYpgAasbA8MIy5WiLb49LXlbtn9
TTO0tfsvalwuPzk0Oeuc90nPqRSggENdgzT0Q3hIwNutyVm4O8oZfk21/clw39VZT+fnapr1WiA8
H1qtL+YzoXihkxNaHWp0s4s6UxSMFg8Vp+TjMN5mVqtHTJHb+sDF3kPIW4on4y3O2W2P8c+WGCIP
YM7c3tF7TGgKf8iBXwotxGqNd5qh3Nb4yF8RkyRWmHYH4oJ3grW6mt4sKbE9Es+kFSPTvhDWRFiy
e9LgPDOn1jd30eZUoLaZ1Yvv9WoP6KO0jCSk70Zg8K/XWBReCfBTKM2wivJWzE2ddvM5Eu6WUhNX
05/GkZJbt1C56PZwBpuGdB6e12Tks+6jgISW13QRm8rYzUoINVIscaIiPHDWtzBFGKCU02T/hRmT
LrrJtZRBMGuipPTSGz/5RMj7Aj0Rpt+xdR4ABcNjv4asIKeCKT+qwonHamq7Jl73CJ3rOMLMrWc0
E900l7R9D7FFVNXiiO20WucZlhXla6MpnISWcNSnEBDIMFIJ28ngqufKrQWASzHjQiWliKqnF7o5
p0V26D946aluuijzKj/TaLAzqCR4U648a8Ynl+IkUCWU64JTwLjiXq+hmhGrtQGylCFODi7kahVa
osp/Boa6hkP8yoiBnz4pHjz2jz+4MxzyxtZYe2u5TsjQ9WgM9ceJNWqhtMpcJn4bjw2uBFo9M8GD
McJpb9MrByJJJwCzxvdbfWUk9miQQlZJEjVV9yQqXptnaBMIQQMrGNIukcrY53N+8Ft4ZT/2yMoC
yyabWxb1jPUERfjeYHoGV/m99kkxp5ItORCem0ErI4VC8jfuJTpZKC0bm8WP1T8/Ornb0quGdZg/
xTa9STLO6HelQHil3twQ5J+T3fs75Lp4bMxK6PYTRP/3f2CoXukabwUUTjAFKbmXaJFxISQI3SjR
5LOzPRWLGIOdTB1xH4NQqgCghOBQIGVFOd5slPF/mYGeDMfDQdghAYONfkT3/NMlz4kT1WzL16QU
OuawAvp/8TAzzKGPB79P6p+rxPEjghJUiLRRf9Jq0hCinrA3R0XjHN9fZ8d9DvtkYosTw3buijS9
iw6eFepizaPXdPF+G4DIW5ymKHsdOfdstGA9vBCgrtYF2QEX0j/LUQkOOJpS71GUJ9lCX7BaS/9X
lKN65ItdS4gZF7ss2PIe0oqDnSKU6dUc98a7ndnrOxhpFXgywiCR9bSZH2Tno0IEeAAFFDHuEpKX
W3FgT645d+ASHHhX0zBiKlut5lYxsGAaVU09DaQSqjZ91HD0kOJrqvxVVypGX74Sf3IqRfeckPko
36fIcOnk1UVM/Bjeg6ZYGtj2xYweYVd1Rnarr6wUFuFAi1A6AtY2LV4f7ywFJuN66hhKv1usyadD
aWvXA8J/bUM9jb8aPPeJQ34X7xOisDLV2cc3SuWJknd/ckvXodJXO9/IRJSJWU2q/wWGZrvrwemh
//x7kYdO2+jz5w754lrJfBBuyeROaa7qhEemI+fntVYUo8l80M3cnCc21Xd6RWAOmKetcNnUXbgk
fQ4FFi700e0iRnpBbaeMX4C6QIOyJ7FBe0m0W9XNDfUyMnDJMMzBa2iPN7s9SOupfbKtALjpDJsu
zQV1BUDE7BOWgqoibF7uM30/LOgRRka5EVANdRL4OTawNA0FajJGglqiRV7Pd3DPHqxKIsnRwKY8
Con5eQmXrmB5XPVU+73OBaC0Mbey61jDs5e/WMMOONTemtP8q4qq9Wj/z5X50ERswEhwRRiH33Yx
uR2dkPUJMKfg5jIF+kkjjm5MSieMn658TBMsCMXD3NGZ/vpvjphD7honPOj9E7aAYt3+8jxD/LiX
RgvzlDKo2K4kV05UDFU+iyI+9OoJpNcVeq/oo7mMT0aZKFtJDPoSajb8KTUrSI0+zeQO49qOEQED
+aN+ZDFqE8Y87iyUnMY+RPHND28P8QaqHk7Tc9g0GyEh7HK0PPaAVkix0EugYFCBTB8MVYq70231
9YvQX+kKtQwXNPC0ICoNLGH3dKuC/oxuVsWuTSf8ayTPDeziEzvHsknpeSNgaF0w7C0VnQpOR1rR
5YwiH9p019ANipNkXqBg1S8G64kyU6TjFiZLjX8NegrCiG4RMeS4c1VoiZB0hKtW4MmsBvTaXqMz
xk4Vh+aNIofYGdZZPqO8exoQVJ5VbjF8DPZ1rKwFbPHZujMda8fmfQ94GCN7ch3HvHm/NLE4x4RO
84i+F5Ot0i5ML7UGa6pUnYnGMjl2IcAV/F82SRTUabKgc6qw+sQBhECyCxfr93yrOe0stfBLuO11
Kg8SvY4Cc8CQ3CSLW5JeZdlpv1cdhYQAAQflAtXXsS0qeoq2CjYzuW73rOW1eb93WwMgy59jR28R
WjemtZxhwD4blm89WPJSJF0LfFpUFjEjYa4xZD8Ge9L0dKLGULYrqrwHrYP8gYIA0/2HBdbz290A
f8F5qe5kg77+JGH/kXSRszuP6q5toVsCvPxaL3cAUG+iUaI2i9Q2HbXjuLwcsLBi9IeRuHPxi11y
YaKMtaNynGKJ2EheAN2x/m+Y5dZw1f1cjBM3CtPSMhQcWEZERZQ6GizWHPCWxeDA+GxFxeNe3fvD
3WFDwAUWHw/Z6uE0gCePBMWySKdkqtt6gSj6in4jAm2ur3X5caoh4fJ8FOi32KVjDMt/b2Ce4s+k
nkivtSdccu65FA8TfTWg3zp90oEEVuSFg+9fi+ZMOX57h1NA047NlCmtoG3xH5GWmPJ59Qo8iZ7H
IMUDkY2EEXZ+zj2TNy9e5BCjGba6HxrEvVmsDKR3zMRO/OIXgNJ1MdydHIw1ucRKN7axlLgaMznJ
sP4aoJAwrMijV/nxEvouZQFYo9pBdA8Sk36LP3sBV6TiVfK9i33e9EEDC/f/cuoZUhEhsBB15jI8
erxNmiDgD2EmTUwRKsRtjdRbhkv1GUQx7RBFqChfZRR0uuC+d4daleOpodA9KqanYcuvqSxSo/dC
//EMlS+WoGIBiKCpFBlku06C1fCP8+CepwgzI9jhPMfc/ukl5moHz3MWrNPvjupI1iCNyfyCDAco
L2z8LSG7zhwvOl45StkOoyJ31tp+oYqUrZpemJ1tLNylVMCu0xX/BqUz0PDTs1wufKB4dulcg3ym
L155pX+JbHfKfj4PhUPBAuzKYBChCfUVG3LSAU3FMHTznpqcFlCfYtV8e5Fc5tyZdUM5v++ZXDmS
6Ywj4c/yv3AJiNr9PLt7uYFf9B/Sw70mLxAPXrjwEdKK1c5QJxS/zgp1EdI6Idu8X52A25LMKmbG
32agfFrJsCWG7Vp8QO4Q36kJ21++DcYKBpU2lWOPgbPYbEVVM20yXw/CGvyvDQ5tIxMjYATvuucY
8uhCBCaKnVIcZ7VG/GV0c3YiY6oJ0ungkk6lkVecb1B3T3r+4xMu1hawGhLdYreWhyzmbVeVf8KQ
26T8S3PJPkzFqfJ+HiccZ4h9LvneJ3NF/PJAuOC8pjery1WUfFt6JeStaGJll53oGdpmOBMQtCc6
0hZKnGQCmldOfkmbwcmJmFh6ZIMcT9wr6VTNWuk7oUTrp3kCKPL2+5OGURoJjnwtqJdlVHEkVZ3X
wH/zJUVg1976UX/Xf5WrMmZ9jzbSCpLpMagb0dF8C9mqKCZFTipFQYk9lX1y1C9k0FXZu/f0tvjH
weyydMOcPxaAq4ZFpdeCPAPelrbbEStGWXmKkDrmnQuBkUwC9etbArNr6V2woN30q/9K4IlL8Eio
oEBA7Vf4wgi1oETh3jkYYAeBhZk/mL59ejqbQsp67iuCXJ8M/1sQIIZFZfmpiGAFEzG+Vpw+CVrU
MS/vqyGbiQIJzkRAK1PBVML1hSD+3AbcI8Gb4pZNe5aUsPPG9ZIFqjZbwg5lYhBgqSbmBrORIHGF
miT9NRBHsVG0RWLl9hCEd2epAG8GkAPMgSyhCala3MVrv4q/MsoPaDfYHjRqkriu28zQv6daPLE9
KzqZ+kKbbrR0fJNCr6tPsDdPsbfQe8EYYpJOVG0S8e08wP4KZsXJOKac4j7O+sscIbLnrhRES7m1
EXYVK0MVoK8D53sYHacyYa7T86eE3ds8luQ3pY8vtaKf59QBODAQZYIO2P8ZpHMU2hsRvDLSz1Vu
3M7EuUWrxfKbJS+OFz+sLnHSNg4u0HZLJ6pfPNnRZ4NVxuxXXw3W8diuUIdsLRtAW9LS4It/t5rk
q7StgA8Z6KwbeLKFT7UI+riMiZ0wGczC3tkGOVWOtT6vhun7GMnxzi7+TbUqXuFn8J77YlU73qru
1JYqIyXhJ962s6PiI6liBKzDKa+Cy4WkQUe3c3+wltpvjvVMvlIGI1i4D+5MRnr/aYiFy65Hraeh
xkPtWIWy+Rq+V4HONtHQWrkwdtpQpPy75Rb9is63JnkGRiiJPpaeuRtxrFP5Ey1SRDOhxctUTjge
F5Vuykh11WrpYAoV+PBIEjC4f6IziUjDBDpkyJ1kj6nHR0QoVML3xL2EZMttW0gUFo0IHoTkhrnC
YhXmpoEZjxganAtByBhDriaIq/bpAWbgAKmaL74AO+hs28QsQX+F9/B6ZlfwisnNIroeX+ewjtVx
5M59uMv9A1e6lgGQYkwWrDPracwBs+9X19JwTvOtuh4Z8jW99Bz6C7Hdegz+J0zMeLuiM4Kt6XR9
rykSECmiNTEct9jLr8Ib5CwTNutRjET9dTS8J576jxNstf22KPodrF+vwVKH58s7Yx/ZR3zbQv9c
u5IPR/+iYjeQJDdbwoFyr2FDOxc/jQoL+0G9v4AWJloKqt6LpJyrm9jTxF39gv/HPHfNPzd1/TOr
h9ZJ45RB4rlMlKP8Wg4Ce8uy9LBN50jDIm6k2UxmCPlUG58ebJ9kRJOi9+uXGWe2URJ4UgMba8NA
2XFdITOch949Xc+Ay9cLPjvTSZUkugYNDlGnqFFK/fI4QQ4mRz7uaOawpTb7E1PfP/l61m2l3vix
WNAfpcWTzhr/kyOv2881I07hpbMxbpJaqASjaWa+2aQMYv/i68+n3vA7gOI444rsaYSrdEn3MmZG
0ruskUbdCToI/4IP9BMYYDs+0DqvXiqkbvZXpnqM2ER/aRGIydlZhcs4rBBIlba8vQF3uSeNlnXH
OQy8C/gvcTTo4i3nwFKcyfBGOtpJlPMVSvId1ApHSiQHjWITU+eQzU4L96DKXgSdt3nY/tdQpXcN
dvwyZtbtYmhC/l90WMa91CqmG0YVxZdYHnLFqOwuDHJ9dsg76b0oa3fltt4DaO90cgzKJvCqZyJe
OqyIaLK79f/0Wnd49d5T4PGMb0MX6h5HcnPVml0dVeWN1OOCvGF5Uu9lA62yf/ced0+oKidfaGCg
nBFg2cWvHvN1xOIWOgz1GSvx/EF+/1TTGiOjvpP3q6E5ErfQ852oFjW0iwdp7wrpYhACLcEzoav1
rRWl8jw/KKOov6MnY846qBvNYR0XW3VkAKVd+OtVjKX+dgEQn3ZGpa/nbQWmcYBvYMFXQ5ier2l/
3UzJ5Ksm2df+DMrCKv64XQVHVQzaqk/ysKcR57NljA32U99Z4JGURXAi9f5jvjjK6eJYFxcvIQ1G
B/v2oTNFKtkeq5T8zKPGMrHVnUrA+Y6ZZiGb/jelXXV19U+Am8H+3jthggEZI4Ab8DOSzoDLJGCL
1MyIzmD/ZEZD9nyFhpfNIX/Le1QnJ7mpqj+lXgx7or4DZPzDtsexQOYKO6P9qCYwWZ5IQF8knt7B
LdzZ/fVmE5kUWojYdfs9miOVgTWYNYnaR+wMExqjK2XDldnrke6N9voV8NnscWRzPNL6VnbqFFsf
ManyLxkEJzanDnnABgjjnxPRQn4bPeSJh0+TjB/NNUhxz00/prx01lVb/jC53Y3qNt8Num+eVPDW
ThzL+sESNVztggOQHhhD2I5E7P+BqxWD7C881Hae/PFVKy+dqYHMeq1eY6BCsXoeNb3dqDWZ9VXr
9nq7ovQHoFw6dbCdnES4iRo/Yzq7orYsQTnG2bo+qKOaPYg7GFpBOpcb3OoQxBnOgUigOP+vZAwt
q2gRO9CliCwQWjSaxdkdRxmEDIH+07oRWWCN5BJ6E/mxKQykPG4PnaYns93zZeKCXZ8fTeucf6dP
5etg1VhYExFUMnRaqn5wvthEbVrVMrAZNcrZKHVfVH8dcixZdG/L5jq/uvYh1G8NMaRHO2q3ziqP
NCbLJ3c7p1jFkffeKZd2rmlNXfmT4AuFkHb4eoMGRc2GYciGwPzBcLf/oRAKCU8+qoq/G8oBgOjN
1loRsG64xBkof6IVwAQDYfjA1D3Ao6OOIfCww3751VtOZPXGGyeeYKfBEt4i/pbVdBrC8fvwPyZU
S1WpficY2+609id2JWCH5Ri0qi+p7ZKykquOvuhFT40zfSNgSjJ+FjNG4lqQGoF97MG3GyoiAx/3
snrrE49UFbzrGL9kGfVsTfZoo6YUFgow/0PlTbOTlPOOUxv/1OoOVbrXhDZWeap9r4kBN5bu0sJf
zMHxSpEcuylVMYsTnld+VCf6KeHIT1fw1b+MDX2TbvB58YrCo1FKbBPI7vgnooRXg8kRLVXhKoff
mow7OLBhDAunSFji83XXwb4hxtxC2jAaUgUs0f2F2hi0+t/orGBsfp9cw1+zejKSWP6idrw4Sbbg
ASJ8fZ2fpObvcSfPUsgWPjavrXkF/DbzMX8BQrj+heT3eQZ7XEtubBhSBgNGqtRlduj+cSyDGxzO
WgJmJD9A1NTb2s3oVZdBndYvukUVhARnxHZVGiUjW3g+OP4bbrG9GJnTncidFGS2Gp5e9hHZyStr
+8vKxzRA8D9wEtQ8KbjX5kVqf8ocsfaekOqMwiTgVTQv/8r3Z1LMpT8cGF0LokPKZAKxkNEc0GpN
lrQ89GD2WM8b9ieRQDB2DXcbEcJ3sfcJ8aSW6CKilHqWaPF4e3d2vFQ0T5bMzb36KUFgjD6zoJbr
afAXC76KnTu0hBlstDYtvcfutxwUUQBtR9+yn1eeLOK15fxVCU/WAbK1mpt1pIevK3kD9sr/xW5F
XA+C+II+u5GLVMOrdyozIZRFCXoNipcyXaKTgieb+BLrm3bnd01XQ2339buy/RQd3FR4F6qS1UMl
QdJx/J0MxKJ8DeKqdjsxdWNapGcPLzmiar3cHMf37yhsYOqIWMKf2GtbrOdLYjQXiSLEtBKqc5Lv
C3UYNBy6VycJai/eccjICbragiL8tGPkmh9xiOoDRiUmolRibWC0ge0FUsxRLfYx+G07wtbuCAky
bdipwqYySI7Fld8/Z4x/gECkG22TXKR5rsRvgOsliByT+iLcj0IlMRgB3DDSUcoLCu5N01f85mmF
9tEK7iahafPraSEeHo1PGhnWdUcdTa83Krm7s13lHMihBCL11qKqIaAjeMme1zFgPuXS6ygEdX2W
qd+UzUWux5S6aVaO4B7hhVbwkMRQ3w09cS4eQqsZPe8Rc8GeaOoi0MtYmzfNq7T/QRX7GxyG2gGh
aLI+zT6iQjJym6d122L9I3W5TS+I9M1Td+bIyi0nSVthxl23I250TVR0LPozFhOlc61TLILq8J40
nFCbd5daPWBhd6+rG1mKrZgkFIEAFVfidx2z2188+iVUo1u+OX+nKe9vrztFjynQW90sQ2dcBamO
PXdNETWBd+ea2zXcsoN8n+AFoG/FlUmID2rCN49rpkDg3cBFry7mc3+IUibijpp9IuZPjJd1c1AY
0M5+sO+Np7h0T5R8A41TqX3a5f6n8P338k+JurtraJLi6NYPwNiE1Hg/bdL3mKouVzMnAin+kQ7x
IW2ykfTSYAczsOkXqNXAXR7aCaInvbLx3b4P+8C2VK06TqXt+jDm9LPYQLvdqEjV/pcO7t5acWn/
Z8p6dg4xUCyMoCgKawfWW75qIn7Y6Sno219Q18fk79aEnFfLRtMPXO4eJw8CBQjxI1cW5e6ze08X
ebGle4ICkiMixI7+BRpyP5jfn3F8xA9sanXROLcMwny8DRCXa9oTSWPG9iWLVQh/jnkQHbR9Ps3r
vEh58uuPV+VzE63uJL4VwuJwOtwdzqO5ucK36NyQ6fFi9TMXYpKBHfXN1M8a2/LGQkfyOWAP5O7S
BPBdVlaFqX2RZZzy++E3M3Army2tiilDrasmFakV3DKtzKo0CL9ruAMSWoonCUHIc7NN8ACDx//0
KRZav4EoXbzpmP8ICpQmmnL0csFsCzsmXjYcynst56ImJpAouJ7FMHLFdSMn4rC9CB4lgIbHFRF+
zk5JEYGgegxBLRb8y3rxA6SI8l5pJf2XOpnjGo/raQR3jlMAogEYmvr+Nd3psOm3/D5Nnkxq9ZVI
MvEG8YoQcdRHclor7GzgeoenT1pf7Bv1b8c7fJifLxj7FqivJBny7VjqSwLy1OnHv5z0Q6x6v9Wx
lyCd9BKldF1xaSoxtuw83pAeezl4ZVjEgkO8TMFNUeFMy1u2euAtjDLVER2PT6o27+jgv27xKDVF
e9Qy/sGLEgd7byX3x1kQdtYXtBSPYpwUpoUyEnMwFGgCIsRKrw15yMtt5VJHToyGZnbJqQKfqIQa
qIXqoOKmucSrtQowYRqxzPbWMTsQNqdYq3H5XElGST9CNk1mbUZhJ51TQ0CBnakKVKoDRkk91CaX
kCwAHIrhXSRTc9FsAsAFKfsLN0JXmIpFe0WwvIcnT/siSWIIsRyEJKhM+SY7B9B6sx+8/Wdb1/tP
+I/4mnPi7sixZ4Nra1nFtbHLFosfp8FVVjcTxec50TVcpKOVwAV9PTk2U15G8pvHmJszzqVnn7QA
dNcFOWZimpQREDigoeVwTeTCXcQgwFjV9AMHxRpUVgR/hp46zSp1sL9aJQg4RgMKc265CYHkmhKz
M2FQo/ihIgSGcpV/7YK+NsZsLXCxgm6/OzDYtydZ/dUtlPKTdiTBZKDYwR2Y1kqeMrdF1CMxEh+R
ykt+KOhVSiwq6dQRd7Rsd/h9qXUMYg+o7dOc2PRVqH4iNLMXz204ksjkWJs4hhIA0TD9lYGxrEa+
7kPAMtEi3x70gHPupIDTZnGFAVCw4YNW0ZSGrjwmxJMrOjYCYOZ3dfJgsc2tu/Sm6xDJEjLDRwDw
7Fn5E4I4PWwmkXTqcqFucBl91hrPRQGi2uYdLdROJMUZhGn6YjF/dzsn9rDGW5kcS5ET5e5t7NmF
rbcGd/YNE8qreZjX9cYOLQlUwT+dXDCD8q6230KZTzXoxHPO4yBP4j7X3uvA4upYndWPWsoHhydA
J5LIXg+6SAX3p9ltMG5ouIXJH/cAulwUD+SwjmAmFCejUOb6V0F0ZwEyqLS+nDGjlezXmoKHA3k0
x/oXeC4RgudBf0d9m2UyvaLhHG3Jff8zYeHoGqsZmzBlpaezbB5XUMkfWu4LYJkgl/dZIWhd3X/H
4RD99g6S2pwhBqooGDnnZSL6OSq/llz+UToNrtxrjUF15be5JB5ZlBGPnI3R7kt7I3kIZU61JQeF
TicK8+r278xRUam4Xw/7jjXgia3KyC+SQ25EUuqVhZxerR8720T7NRgPONRqGVSORZHiI0baLAkF
y3RTZ80SrHcjxKuKBrrdG7THP612NIWMl9CIPVmFq0qQYyR1jfzRVlfh41xaaS5RodI3ytkzwdsO
/1nPmlypMiXsvFJSlMQ18qEz6dN88j6jvJxX3NtbholCsOcIfkCNF6vKktZr7TSqHySgonjeDd+r
Z33ItOAtuJBPvBvdYkEI0HyUc1OAvOBenBoqOXG6lxQ6aMjAfAKB4QT1wqiyn/DBTRDVA0xOeFTt
LrN6Q5slC7jE/HSEEMvlEYaVU31fAT4KeIXA4GhktzyBqivuCaR7aBInnU6uMw+GcJXW7mKyHCXS
/oPs+wEn1y6t4EkAXb44HN3RFiDCrllJyXV4zimRPM8QbeX4Sv8kq6lu1jOmGT8Zm+NWCiIWO/m6
Tk5EHR0aQNLTtBUCSu7xsW+9/e/prYyon8Dv5ii7bq540fiPa57zbIKnL95uYJHra9TL5jT1iGXn
RbRVhchHRHKqiC7KAifmxpRpqyq0aKrsZyFjWNjVtUjwYJgGzkDxyKFR99hKYGiiBMrk2Qgwgl5Z
bTwBafJdZW4Rj/Sb60KvkdN0uKe7eY0LHEgoh+Xjyr6fvW/iwt/IQ5PF8m4Gp9X5XqSd0UbayRH2
5dAUkd+EPCm9NOKLYoj7IfZtXFOumdpScV3d7l0l5aT1+KzwGDIUJaEZlj3X6wicguP1ECHyZrFJ
vYXUMIkdoSBIPG5ccQm7TZi5RwuZOhQC3ydtvf/ruHeznZTxyueMz2vvp8/6SrYyNS6jyhZcVPTW
NNxDV7z1+cZnYMHlNxui49mgwY0bQDtCAwylVx0rCW5rfJH3KzYfcSOnppO1UBocRCVrTySCSGDf
oHGi5n9loQ00PYYpxiJpqx/8GrsdV8zrD+sQxbw6PR8jgVvNhF9i5VEWmbpg3B1/2vzA2Yx79Smx
YryDZpCwrbB6RlNyvpSnRpkCMjtmpHL4TL0qukAd/04TgQU/1wSPlK5eJE7DaS/tLnUjEPJVA+qs
8IlJ3/gU/hHxG9HmtBFpBlSs8hTTM1ZaEe0N8ozqqAXPF1+1SQQh+KSJp3DLDWoOtvEHcmsejMPI
5FzUCtx4IDKQP8dbqyR8kX7idw/ysWiDFrF/qz7LoBHK/GeSUzEIyu17a3i0FZA2iuACdGxz6XEa
Qer/CdANajA0BtchiFzHpPelXCHwnLdEY5QqmRGoNxL+EXNBZiVZt8Bk69PhXaOKkF6XD5Co3b2e
TNCekypaj1qrJ1KlnAupl61poGvrdllQ8PS63l0OMACdSkqdt+TrJUtC60p2GnJqKmgYSyYqoblO
yKRADlve5YBtMux9ij61gYKJ31FyjBBj56hrLCNxmStz9nVLQ+sboYhGkF/Q+ASzjwHF8cAhiS2B
fIvmzWtRqmhLixWgYBnzLY7m1R5JDQSbrn/1vvHbn7WDWLAMLeOpfx8wJ6yOMCkI17kv5IZbAQBS
Oz5h/2WdPhMzL/6EB+qBTiEAlXOE23HhzX7Cq/IyNT0X++EppSSqfuoWFl59MFWbUKpdj4ieO+AR
h7eHKerDh4cpVoMtjivxPel10TXAbZHPu+I8wEibmcnkJw+DAx0DkvyGTonYuR6Z68zESw6Odw0F
Me+d74OdL2mOolRTCUF6OafQfIJXRN6ABooU1t3veosAPd8fYv1QJtf9zMLHmiLNA5WxY2oBFfoJ
doGvfK9btpCQfCkhsZusNRcKxT1TTsXgulwvZKD/WBbLNWlKVsprnS0fBuwPBpoNDK6crvtaoxmS
NbaBqIgB/zNGB2+fJyrsuHBrnU6pOguDWyP/WYl5Gy9hykm8Rm7GDVSfkMTdp90RN0kzDi7EkfZU
iitexiTGA+pTlQIidDjAKLtGp3pgAeG1guEEev6+It3L8HOyEBdA8mtFUM58liYMI8/AVY/Yzi/a
3ZfE72A1bQ3A5fRJrHDX3r5Q8FoWImDiTpk56U1WepEwiSZvP4g9Yg3NPHDp44k/9T+KHwLIHpHe
Gb2S0J2zn9YcbxZl8fGThk7AdBHQ7uV2bnIb1WyjqlROm2OWVT4dtbxw2moVsflELWK1ZzWoZx2l
R3rKE4ivjjmiOSI9de8WqXE3wcRJTosiTox1lJMEXQ5rV+JwXYpch8liQShIJooNs0ijAvTQ2W6U
r+q3sqvRsTbHtEkNJIJ4ATVe4MCIM6T6JhjZnfWm5M0F6qnoyN+KKDzNVyYjRMEp5J3NpUhynplW
7rhXAE9OUJxRw/HHoVFVdMcUHowh5d1VUGL5AcselXjcG9L8vrQmM+DG3Ez8kpI0rElaTVXyDist
aNL2OZwNR3UEOpwbrELSkug152LNreQAnaRN0cAgjun3cOB4vYKUTjQgOW58u3TB/Gur9dGoluPN
SnWXK7NGvUiSN8pmrlgpqBthqhqb8ZWHf9cz+2A3RrdNRObqBWYcK9g7mr+FSIeMDOJteL0nFzlZ
IWj0ihoGSHln3IqYNvSlgrPc0Un3MjMYZOLdCWffzue5d3k/1XrUU1PUUAKcwMU56iEDuo7jwaMy
ohSuhhfiDytnMQEctzfPL9FTIq2FABlPlCwQe03QacLeyxrM6A6H9P7mo6boikAg7huM4gWli4YX
NcI35cLlgREB6FfbfKTtJOFovh88EuVvCck8dGJDYUtTM7kIgplXawM8FB9hylhKELE2MaLSvNez
O6wKvHDhib6Tfp/Br+Ci1nj71zHo3gekGc1cV0VthBEK2ga4OtdmrBHxdOYHLt7Mj/fs7BGzUbLc
yIILBoR+wGcDtmW5+Q7LsNkjqbIEBjb9KrVNnR9pj74u8F5uVBLsp9v3YY4stgn+WXPfzBXqtpKW
BKC9hS+PbqMtnvUu4644HKUE28+g2oZzQMtgNYU4WXuo3UvcpyxUrR6DOQKlPXmEQQ+o+9LQYaQO
yLNvI1MeT168Ton6BMAu95YAP0+fBO+Ika7r0kx8z/EPLWmJqhH358tuwSPKlrLQCtXQkGo00OS9
kUv4yjHMKfL/ZauhjqCC7dEHcyZrnaH6pjZwqDRU4MRVL/zCpiP43llfd1UYtrYDOfiQOKSJOT5e
VAje+4a/UJYxO73YvYzdSSfKOhAx5f3T3fFblTk6cNI81/OjlCa4opSZ7oL8JQMDnnr6Sr5jD1Lf
4T1Sj44//fhSqFZVOO+AUDnXsSHi7Scikr2SWo9cES030El+5oPukP+pdCs50d9UtvNA6uRmFhF0
QJGQcbRzQ2UaSAabXgkWN8Qv8o7DNA8OOsqQAcWbmh0j23UHOn7w9zXOYrN5eb/BGO7vyGYU3gaL
l6ZK2tGBKjh3ut8wdROheXeCNbPPeXutg+XtIfoOwWOt45uUmNEgftEsaOFFua/7qBdp67VEvcN5
jMZ2umw646uE2eP2t5EKsw5fGKLnSnsz9rWV4K3dLuXrl+C/6wo3FwEbkux7eZSv4ZioztD8YfJ2
d5QEBhVzdVxpU/V2ZeQhzDAfC8/KIaHFEicvqIfRlCNkV161AGfIqReKC8u/T5ttzcTDtWkXWeDo
n+g69mYLA7O079TTamgzt7m5tBDwqgjp7zQT//pxiF+OFeJ6ajh65UXVUlIfBc+JvnM3n9FshJ17
4ATwhqTxDO77eLADjO71Uw3I7l+hsPAYzWkctvawB18WszMihX6xTH/6ioOPDQR55/N+8llfc/4Z
RF3GS2x2fJzF2v4VDaOlPA+G+zz8zepMRQQxtwTpbq7VzLWS9Wl5nyRi/yYbOROb8qQY5QqCUee6
mszuvqehXFjOYc/yzenchpUmSA76hUNBI+yJuysrt969umc52aorDYj84cCunPZNpCqYhPkZwzhg
PIklH/P7QhZu7ybVtci/SGrtByvVHEhHN270obekeH/uE23Oc6Z5voK3GFmz0GjUFxO8SEiB6fio
c0iDufQwnLcHspWNjAM4vzLWL6sWgwbarVWAs9gwcvSZ9cZw86ARMMOMI7lrfIlefWsnSmSkVy8s
U6JounsfTGQxiYfeHy56CilNbRN94sa5fODmSKB2WCXH/1YJHtFuA12I7ERpYWc3nN9fx+KSA6mm
6W+1AGkdds+Is1QKh2N+V0VbgyP91zqBTVJlz5muCpjeLelK3fyGgSqNGhfgQMWbcpxgp04xXMiD
zfechpekitmLxoMSeEHwoXQJ1+SU5W3T4mXrrdqUQ+UNd9FBPkelBfeTA3/S1gRSUUSe/t10yHKN
XfAcE0xJNc+RJClnrE+A2cdTmGML5XLTyqozIwOTU1klldOUK4xNfDD006WvcKC12AF4+NoMkOdI
PCmxW+uvyVdyIEPc/mQRbrVsrC3xvU9RC+j0BCE7YckGnwZ73orRJ6QoCNsCFT2Ivng1zAgbKIfL
7UnuyYuJBV0Wt42sekT360i+ovHvBpo9RN1RsLtUa8lVpDZcToay06Z7e7vXp7jQut2j3TXOJt47
tm2qYcaLoYMfCMfyAT7X/B4FZ34fTUyeA7K0UYIQmoj1/bSDfqEm59I54w5sGGevApBNQeRhZ+UV
Malyknv6OkHOVhTGjM9baZ4FjtAmdY0mrMwTxWTXNjIptDxONA1/RJbF1OvRhLG3GC4q8oBgBxYs
5qFss1JvPe2a/QEWsvqnhWjZWag3z4mYs9LWHHnNT9C+cNIVfElLbzTNd96TlvGhfyxkPpC1P7/Y
xCjcJ9YZInoc8PwUgw++duRRZG9AeqnU83hMHMmtg1JwWHz+gjW9fAUMh6i+lPhLrnSuVs0C0HvR
6Aoc+QsMPoHLtAMZU/zAApUMNa1IH+h+wOWNYlEWC6+s7pfSJmFEkeelhOrD+skukfgkLuj0J9Qe
+hSJ+DM9Inw4nfeWIwD/4yeUacivtK5CQG9G1ibq3JeoPwvlHG0ix4zd49Xm9TnZn+qNKqhbegCR
p2TbDoDfbXrQI59SC37xYJQAvt/C76IlDJ9QzbVQcDwrJLx4hkZUqr1JLGhb15L3gN9WsfRYqv57
A2awpqk+GMI+N0B35MA31objZJEa2xRzHgIprAwgAvjDdrmJJf36/47+syBple7W+DLrCjsKHxn+
J2boWmwb5a9lsSI0VMPw8+M86adUdMb7Q2u9TXmU63B/HtMKkHCBabPUoejhXjUNrQHAcnyC2Efs
cRZdrvT6zYvgDslklXO8UF7BkdBRrQFpiB8qGMm7camt5+LvMDj9/7gNC7GAUrxHR0CkcuE35G5b
i4CwA8/RrMqn/1hr17XSyTUbrwoqHUi646YrvW+GxGRlzlch4TWpiCIOxxc8eYiHERSetBNLvdSY
+6O+Snib/pZXpfp+v1j8FrmPweUQZjlBawy1ZMt83LfBAQ3TIryuGartEyaBTXm42KaIb1M3pBTY
6NidTdlSLPsexlbytHPVXzC83NFaXZJNNOzA3e4uHyAvU/mGpEXremXFc1DRubX1wEIUzVzYGYWP
PJYgisQ0HizBRrbvhj9ZFMsDb4GkUELMasNm00trDZI2k5Ql3RQ4B8NnSbFFfevR5GGOn7yKwBtx
LiqBAhfCkw1oRHUmfZ2EG877bNovkqNSmJHxjzWpGIc5PFbUFz30dGT4ICxzeMAXlqUJeDNMvmpt
FCtkZ2bLoPnEhHfo8jM2i6UPTICbgK8qiW38Ujx7rb1mBDrxP2edj/8b6P1eD8Ch8sZn14lVCdlA
ys/djPG8wL45izdLYrPvcIaaq/6NVC9ohlZFOKnhoP6g4S1OBWYnj08LShDA9r11DZkVBG5igK6K
NrJCR4uZoG9kRmVHnkiLBDpl/63OrvaCvUrHJDYM1nKQ8kn/d4Ud5iD/N0aa2r79YBFNSfuS42Tu
t0mvMkowkPl1O+GnSyFr2MlmDpYl2SQ6+UoLOQTOnaQrv45z/+4PWBHQZD73BjhKTyRcwrZmPX8h
XrHVquwLIptydpsf9IHfyWZcQjiE84lufJrhNhqh3XJf2IIJZlZGGW1FH9+TAw8M0QERlwhZclQG
eYP79yd353IHBkDPOfeIciGprpjKSqCl53UfjkI1oAQcTCnH98L76zhVLWlnnP1r+8xv9ALeLyqM
h94Uv03oA0nQXhoSu4wJUNvWlpBys9La/wCxpTAkHtmE+UK+sCkOm9Eg7zrrwoQFpupOO682rt2I
89KLjaOonvsMbFAgcJKQaDzccUzjrjEBKR5RP0II8KwtBQlXNymbMLI5fBTgZ3VCR3BxbRskHjJn
M7AyN9NWZvOIggq5a0zaYdMsBDQmgcHyOEQLPH47lHWnD2yXMf6+bvLyyHp0HTR1d35KL4FAD1Dn
Ryk4l0E/aCf7KBn/dZqGqw5NM1sstqdooPxvgxiwFdVthALIn2d933Ifkaf2KlVrVXJXxGEUViUz
mvNxsxKc8XW6R+62qHpud16I+zqYTJCeBNV3qkLR+A/lcvY90GoeBR1KL0XM3zyDy29VhZTmPKrU
aRRySAwvhreSXkN0T2vpqz9c74AQUvWtao+ernlh6dBsWOGEyecBPAp0fmFO74Uf/GkEJqPRYj4r
KtfXBWQUqsFgxHiQk8wsofHhN8HjVJRFEfW9iCEMnHy463k9+6Dn0Q2sl2ZsCp3tI+O2knH4vLtk
CFsgaU0a4CDDn3bovgdr/YlfXwYxkltAUywWjwlVdaVfBXZemoie2dxgNfFnDHaLz5UJw8/uth4i
y/xC6JV/ycPp96VJ81u9nl0LGzGc6lzGE6v33/EIXOiUXUdxEpnjxRUXoP6PImvwGXNBhXlOwq9u
DrSvBmhCqxE7lu/0niF69F+aiPtY5x20lvMj7KTJyN2MDMXWMzQfnHAipjcU6Qc5RqNd13Z85tU3
T0s4wUNw9lTCLHBoFBuklL8Um+HwoUbV140BziwpId0zGrCawWV43e/bTZDaYc+vg26h7PF1i7eX
fqo+tDFDoGCxpBNgs4kSIEZupzIA6YOXO0z5tqZWgdA5Y2MzOCwcDz/AWga4RIvll80pxJAvu14Q
v/ptXdgIcOk+NL7V3GXdg8X0U9zz6hB9zUvgYuUFwNaXE1z6yQgIz2aYm8rcI+Im5sXbXYxfJIpM
Xjl76EUmWA5JoTQqXjod417QiTTbiDE8fyIMSowY607TTkz7n+32ucLigwuiATWN1N3R9BINXedE
YZQQjYFJ2YA9mmgu3b0w6TR8MmYObWIxFTRWpd7bDNPdjnHrFRH1ku+UMR24x2pt7fnRoFTjz1ac
WIuwHgonBrMy5SWWw8QQuP2KTF8VZ/R4ry0PjMt49GhWUambBhK1rfQnXTSUcprxOIkWlrvJmhzu
8597rG8JLS1Hch4Pvcv7d6Zc4ZF/4sBSEkmzCRUZ8RClMF8h3hXa2OEJqUwEL7rN4GWKWsIEw1LD
qPBb0kQnYsWHoAl0jAlgH13FyIAS6xohM/IWNCZdn/U+0yP9wkqvwRAg9AFZGsiaQULgzmV81Hj8
1pIj8zYgYU+ofmBG0JoKCOMs4d4qF4yIuQ9y5xH/eyN4jPV91LeUwtir4mSwjbrb+r1PTFZx3/FT
9jEHzNy0y//iQm61reHM2NSzvXpZrQsJcNcnwT07t+15A8bRTUG+LovB2lSkIUa1IkW4zHHJO38O
PS9zyvr4ebhRFBpEzBCZGZikZ86WedDtQaGDH3jgv1Ou9UX9E9aoBTeSubWO80pQug4M6yKO25AV
tSJYp+wcXVZB7LFvnYQ4Rf4kvA/I+Dst4n+F5bjsJPpnd92jiNspofovTyy+lGoZsPelRgzO80cw
gBtg6BSh+eOjahNY4rSzX4C51xJxqNZ8oYjK8WXrg+sSpchrjzb8WsQMMFmzec0ZNRp0lbOFuQtu
chYGawBIQfy+z7AZdPtfiaK0gaP1eZMUcmcbGZfI4Q7Hp5jZ6joX9IpMia7lhluTx4ueuysadOAq
ALJy17DxSst8Yb3Xpfxj9WEJY2hGKvb28hiPDdUAo3ICZqKC5z5JqSLjnH5/TMzeBjUIPPO0/DSw
OnhFLoKvqhjHVKU3Rli5goSqf28jQR9e8+gkNrTiDqToIU8x5r7/nYDhkq23teuXSpOwW1aiiwsi
8VvuD0AGZoCItRmZvHGP5C4lEG7axgOTq3M+PDAo3pMktQNDZY98kCF1O0K6kF27+aUpBaNA5DoA
LKf1a/toNd6TVTzw07f7eUbVjqhlwjroHz0PSS7nFcMpDUfhgINSmLFksPD7L2+jaXyrU/HHXl3T
ivlR0xXewdjQf9eR7ebrXRqcxQSy8VBHxlJwLg53crHHbZ9UPJ7LajwUqyTxVOBDZQJViJq6yG6/
ruQsfToiXnaeluwMO9pvREKvUcgUnnUJPn1FtXDF5Q9jno/Jox9cGrY5iQWYN+sc/Yf9d8RSqa9l
GKDuXIKgXFROUoZcUv7RGRwjvf0B0YByQKup+e+04erMRhXM7UUYSL813zSLaWjTgmtmMkHpLgjq
GoHZE5JykBOC8YKZkI3GFv90H3pqm9s6D9eZ4rrXnO6mRIEAUONcbpvH//+EgVKNHpfV8YLizHpD
IwZWaeQWsN6BnBO5YmZjk3hmkGs/pFmVVxWSXLeN/x0wCzmlgsKDTdpyznHVsCwxl8UzFcRAVDD8
+RszQqqTU192YYxzJwo6tqpZftICVTXZnJOaYmFRFHic1Q1PJggHSysMqIvVRtcGOZZWtvuk4DG+
qwgzdA8AjAJBxjQnA2HrLr9TH4y67b5vxpZEGxIULLU+JBsKq5FDArHaOrdcS09i9uac6S1R978R
bNnIS7z91Ef2rzUsv6ccxoNje+wOySbwsYcFYOGx2x5cPO7gsO7nPIUqtC1wK8UeOlkPwr5JDG60
anW1AudRAqmegzQjOscJSif1icH2qvoSb+THle19I5hHU0n02+Gkd/8ku+DdqiGkFI0Mo8FcrhZf
AbblCsdF3soLv/AOfBQQIBftlbcSwnHI7RIW7A4YQmtW7Dak9CaAeQgXN/ikDxjvlLKu2bCiTFJz
phnpVWpacGqNsvGsFqGV2u/kC5ycQJZYqE4nyzKXjdZNZa00d/gkv3W05dSJfaQITuytSlZS9Rto
A5yhpsrLsrPLajohtGXnpX48nxFC/y8o3SMztQurpdPiFFIHf3+j6BC3CGD1rg9c6gGaWj6eNtJi
xW19KifaHX4cIMgGO1zMDGZEpX/SuvI92zD6LKF0CIoz/Z6rl1tZ+CqPyybaicughBo7iRVtUa0I
CoUUopONErRw6gYaxkbYG1bJadWfaev8EcD2axhKaa2ofaEaXvzEE2i371+ON6TuFN8ddtClAwKf
CNwwIYzCuJ3wHmQV6n5MokyEx745OR8GMmjxXddQtWSU3SoWX/bMaNt6CIGDofSQeJUebPV0iUDL
Aj9JZmQDxImA8zZeAhDltFI1Swc4ZKq71KfoXvnalvVFNKiPh35epggiTi9HT+NrdD5FDFBuqyzF
WBL+JfEXS1Hz/GfWbpHvvmCjonwjufJcGPLnMwBTaSQQpGApj7WYMIzFIEBMxtkW9L46/N8UpgjP
oJhllpl2XRKdaTET891ZPgUJbaNjInJI5wgiIg1D/8ZjpXgGKeKrK5Boq5MooRxhF8Vmp03xm4fT
AkpDcUuDYUmEBfz6XkvM3FVDDgLcfrZuhMQrH5zp5a7Oo8F2Rc0ifTavXGjVNpHCEpG7FYFKobrT
PzHcA3mOCVFyV1J8gVZOzXgGFDiRYGCfH6t2tnN/g2Gd+vJcmt8Low3qnCNXrYkspSLgvQK0HxEj
vCYZeH28EnApNZC1viCMuPCYr8o21/r9HyX/pnXFFs7829WOQa7W9sIbXu1eqwiZFB1rAXdssUhx
jX753/JgmLFwbl3vCVpxd6FINRI2MZxOeLZ03wy4IiMR+r3i+WcK3WLOKy5BXKDwJndaVDi1KPd+
JIZ/5gLYFL8v4WSt63C2Vfg60ShJiT5IX7ZbHmXrSfy4XE9rfGDWXZjsrV3dh5UGOK7q9o5+0hHK
+S3M6RZCrcbJ5RKL3TB/5IIBtSKOcvY4m30aQu+4ldrM7MCqBFlSUNbF+kgMkqZj04h5nMzuvaRt
YOuKeYrbor7nTpi4JheTfb4Rsah/WSeYP1cU8Ym6XaO8Fwi7bPkE1hjmhyx8QLyOWgkRcdSaC/ad
CBH7KC17o0hjPKmSXgTpXLiIJELZsywnWp124p1AW7gZhSabbZT0QpcuZvmGtoqrJ5JyCMPmPdE/
xf0km+E+noYrDeKjdj3Rdc/JkX5P5QJx/XxE8M0SKMqp3wLHi3HcgM0MKcvXJHFV/K+eFRn4vTKQ
uu5RMqI/yMgoTi/AxerV6fONBA7b/a4nn/vE5RxhPJQrrY4qUPWRm7NxpQ390FXLj1DKzAzBjMjU
/oogRNQVdlbZQLdmjxvcaht4UbK/ZygSt4cIMjS9Qzhaveo1vep9wr7Y5On3Y6f2CBXHhRwop3fz
/Dj21lwAsLgAtKWQKwBQwI53QCOptUbzGFSlFXbRuwhsuB7K5USE+EFZcU2CmqOGBwTfbCdwVHhM
SpyJYSo/lfaFL2Aub74yTDPBum5LIF8tFgq3ZOmtFQd4lEfyvauu//27PChQlemvALkpN1+KBDO/
h6gPiBB4Nk0sZ4gtcFJqO0B0S3JSc9MUubNmmHQFC5HZO7V/b9/YCahFLi+ortWQxbvQSG5DFM8G
mZxUiOnqyTEL3n0tA5kfJwUT36lb9seDj2aj269ZLlsnLY3NcOmVwQQumTx2mRjUhZX2P5rmkcnt
V3hXcqhVyNrN8FdwjI4fMA9ifukipbLSMzb6s66UfwFchKxsgeXkc4dPLXBWEegcTu0VfDq+35iV
s+FPnyHrJ5Kzj0V9E+wKcjjgIExeVN44Qg+uTn48+SoGB3aGawmQ7/oJALPdZZSXcRGtgMWxgvD5
w9RrV1ihuH/W3Rj/MnRnYlaCHG9XVMAVJIKmNCAafwW+VJOFBXp4HJdDOlTp8BK5+5XW0iZh6Qlv
vn/gMqpGjdxO8tepUWN0PyeBLoWkZsjf5DnZ9CPxqYoXc72GAzxG59xWAu0CI0qqHauMFcwXWlbV
7+z0d4NICedJofH/3hsGCQK29Vd4+WBtGL1R9Pq4wmDNgSpq0VLxuJ8SfGLyYCtsSW3jaAinLwBa
ce9whINTq3krv69QKJCPCmORa+zldCaZGinObxV2Bwamam5F08lQX+BqGFKiVaig//HOco6zIHZS
MIzGgb6muT4p95/+eqdx9opHAs82P3X9jO/7n6ObOkcznnjHk+X11deQhMm7W2mlhOx4fixNl2ZC
Pu6TyBIkrJiXZq3EMavIieVNJUsIHtUepXY62e6U+ywqaXH0mPCFZtjRor5aHrIdAc8XETyONdpz
Z+4Lsr4iXstXFw1qv6pdSNbC+7b+YZWOL3YvRYDXaPDUOW4t1lnPDVaRBtf9gxQK4DClzSW304In
ll/zXwKSCGlfb/5qGWF2IMgXbqfTdW+oGtSPUtVtMfpn7yieBkVePQ2q2sRK01OHfX0kX6U2U9P7
ly7SdAalDUBYxGVb2Ba9Q5+drdJXoVFmW7DRhQbLsRI5bV65bxmFSTZz7qg+wmYpBPK+4IytK7Jh
GYplAZLWHu44vkpXcY04eA5oiGliGzMYMT+Ic0V/ZGb89+buAbu3NZ275LnYgA+6HbvMEAiFCQHc
dwZUQ7RAvjKHY5OCGRf2STY9XV4vIDuhn+CfdI1HMYGVyeXWXHJMvQ9i293lniPMuwUS20980RMS
IToEmB0EvMbB/clz1rWdYUmNweCMd/a0ML9DUfA3ElwJ7m+drQNCZkrFh3iFUCOX6ruCp+VuV9wQ
U4oqbsrbrMgSJ2WN6MngZD7OMsBDBiQ7pM+v44G5Wnum0vOONVJhOhkgrA4aCiPwsL9x8W0ZJwmn
51tBvZ50YYdf1S4pTCTKKDj6u0DFcPdRkGg7v+/2nIO5p9OEGwu/WvcYKH6w6GO+EegyeJz+/fY7
SNy/BoiKVMqvMAq1uWhB5BHa9DtkMYV64OSNJW+NizjwSERilpWaBrbx+4cXfDE9WN/uTdZxENBA
hLlTvrIMgJEEY2XkfyxsJd/kvjg5xm5LLcOQLhMVgZ3jJutAYlbsN7ZnioM22sMje/sVwI/wIQ+1
DJ0nnZpfZKSNz/4TZpm31eOUwN0/Q8LSSRCUacldwxTMLvDgIR4Vgb19zIqFpvwEqFwrBOhh1P0u
qtOBLKAcQdQZf6YElHpEZxPEmiqr5e/o+OWDuLIyy4crjNnMCNgzq/YVweIbxesdQgBRGIpiYEq0
8F98Id8zVQToQ88SLtF5v/w81PgHpM5+rXieIDktZCU+6GO3ZMMrB6iOsV33vm7AmewcyjaeAQZF
04zINWFdyLblJikfUcVsN/Qb7D2oA5oBsRP536F0Fjlz3JeTWhX0ulL9e9bxRMWpRA67HPZf/iCQ
VTDgaJQY4/wYmrkGo8QfyGCHRddUZsCZRlZdbMxLX/WtnAAk/MDCst1VB4Fnb6H6mCdC4U+IKGM4
UreuTK1yJxrDIlkPAZJ1coyw/0L864pfqoUX7ajtrv4g61gWAhfZiCFGguO0snkTB3vO8IR/bCGW
4oWj50Py/gVy4BvXxldbH3MG264OeOCSZOOtW3ej2fkT+2YZRBIm1pOVe1ceHH6BlyscIk0meKHV
oy2utOksgovvH/Ds3u+5lykqgKqfL1JKpi3E9cJy7uYHhg8CSA0KLBMfILtZ7L5USo7opFT1rB0q
F2ozYICVg2fVtf5aPhrIrT0+HAZUdi5ajF2nBDyCbM6mhnX3fVNPzzmU3laE9nPl70iBaDl7+DfT
vIn6RLZ2SU87lQ5bHHYHwRQETkByIr59zLmBqqgt4wO55B6roqz24VMfAzF/QcqxjHXFIGRrYzeK
nMwJnbvAeufS6EmHTP30IdixS5KoVAwWh7wc/VA3ILTVd6d6TJfBunfBjjIvF0e49TUz3RGPvv9a
8LG9Q3WlRwT7W5DVqz1dbRb4/1poblJJRevdvgLZyznILTnNLKrA4Z1swWvqG1tyB0CpHdRDgp5d
GaCDpnWRJM8O9BLS47TJg0TK82HwKv/UeMGTZQjY0Wkj//OUWevdm5oszMYqaAWLn9rtoe1cvAgA
IpVhv7iKnmeWgpUNkhsv6a3AkzIlChqXeHLPtbSJ+TiWoPp18h9fv/ylUW81bCKF6CKy4RakCAGq
iLOtp/y6iWMzT4sEKMio3H1wiOAITqXFGz2M4QKWtqZgP1XLjlxQUsRrYz2JJiBrFaClk8DkOIy4
hmfXyUF205HFRyiFV/9Ln1I7hw7nLR1CnCra8mKkcYOJHY9Tan5+Ekb4x+ak1ngLEJeLdON64+BG
TYoS9/Uv2sA4Hzk98w3Mmk8mT+pSAd5CYTRf1v89/mets9w+ud0qAyjk9SQana3L1MWRz/BtJWFU
N9Jtt6/XONpZT/AdRfTHuI8dOY2ddeiA9k0eRX2mfFzmGDCFhCsmfaXtrNRBn4gB34rP5doi3uit
2EGF5uTuPeQQ+lvR/CewpfoHBQbvDxMfiOMZTtAOAcu8Z+aZE+Nis9F1spwpvgxc+WWvcsih8Mvb
+uKfLwLIcv93n9CE9db64mA1FPPsFvplXFy2Unai8Js21/pdk8Hs+cLoAiUbjhpUQ8UEjPNcEIQS
6//Ogq5QtASB2FCY4gqQxkHvNocDWKJsRdvruqFi/RMl0YyYGXJ6ZHyWqcMSBbrZIB2pwB7N8E1+
MIfaAfvSpPNXdU3X27lnT2xSRZWK3XzLfzizsJlGe/ipb2y7Ni80cZ2lLvXukceLPpupMEKB5SVG
zKSiF2kPohM5ic8r4YnQeCRH1UhSB3Y5LrJAL84aSDCUOFfesu8lvte5O6WvnzVn3sDMzCK+yL66
DNVb21iYOzHzu0XaFAvAQ9A/bcnve7bI+xjXATEL8pkx6BbdPHgzUj/eGvVvPKZ1tvaVarVRCOYl
tYpIEl5PwKtYQrabRsm4q3r/MsHVncluvfiT+ug8w1f2Iii2eIfZ9Zx7gTYItk+r7BXfTXZs+DHd
2LsbRgJixYjYHrjOBdwzUZC2am/B+AuC0elXQK/kaNeKtFLBs8jwmLrPDFvalRX+hfe+TXfNwfCP
Y5ugPrNdNiOB9LsbdX1IYcD9b/7j3kTTochv9dA3ES6cqmrAvauS+lEc1zXgGycWNmfOeX24EyP8
r1XLiOrkvWjf0+fHDOXgRTiL+eHu1KYZdH7tppIY/SjE44LaSJOpFia0SE7hvwpUeivABEl5s15D
T33UlUIp2mjniNDqk07WkGep6mkk440wEKCpXhFG8DFPypnpyYhp4UBOSLbZksWVdflcGGoH9aEi
nZ/WhiGIaHpF3mZcGTxyI5tU6HI40dU+q97H3/C/gjidGlHDEV7Uow/ZxWGwxVww8UyPqpDhqXxT
Y51SMRnEvdqCS5CVXngC8/ZL8PCoxwA0N4L8SgzjuLEMiwmCF0ppBcmG4oEZzLwJhZyG9PgflgZL
B76QLKilf5UYcK1HEszaqInycGHWpX+Jv+xLjqWdtRnyeEaierSfhM7XLBldXQb5fFmTu/gW6zO4
SWIQJ9MbHNjHbOClQNPzTXhOtU2KY4ZzkR7zwYa8MSmaiFJuJ0tatwcEphlGrmyPGztaUJjmhtHF
8IvQEgXAKUujc8qAd7d1ynTsZwNbY0Kna10yjO9GHja+fvXuE081Xd/xt+zI3P0uWmrAJyhwAg64
1BR8NQIIZPw2K9/iVC/92VwjDESCqFO3MvfFaZ8zt27SJlBjRCS7nEKTn6e0dzrSM6lultrDbkAV
HiPE5tsQrB+NMyoAnXt86s4+oLBel6sXjtNewHmq0wFglF3o1c5sOU2tCUrNEeQxTHBFP/ma6HG0
RlQBpwB+fAc/o8+5sq88kvqAH1H1owlD6gDvNlyCc9jgAFAxPhylCKprgXY9Pv/E7wUVfRo3w/AF
RTJXxi/iy56qdm3H/D9cvmSt+oPTb8O7t/FLsBOjVKFfjL0ahPfXJz3Cb9ojw3Vg/GMvZIFWyr/t
Ug/oLysr8iy8TCGOkMNhyJjtO1RvbxURmhiT8agal7l8J36/VZHKq5dK2dPOXqwyUfjOWuDxRmIO
RKSKRG4pwNnIRLyZTPDpCYrSG8Rr2pjZ0wkZ0FSVJG7qjsKtphsBW65jrA5NSdbvvp6X3txgalQc
qZzC2P5XOu3p7Wq/X/AhqcaTdsP05KnsHkjNnpYbtqLvHt/Hoi1/lvOmdB9IjoVGh5aliv1NaGng
XcZNANNSxKNELobWsmX/HOYfiIds4++W46WS7RBheL7wbp122zRn5ljgZRNy4GC2nd8q0Uk1r4Ye
xXWMwppw76Am2WQNnbDEKllXkwi7EduMghEiAVk9s00fS65hrn1VchrOA1hGvcqNXRY0jf+bKY7q
a94PQp99IVscz9r5XROPPtCAk7oX2LOafyZ7xGjOmONqCE7XMpVDzEGdfLfEQOCKA3oGGKcO1nrS
WHLk1e0dj6oa5DcDmpYelLbPdiH2s7pBSWYXUZLL+ZFViGGD7LqYqS1sDhYm0VAQYRfGui8YqLoR
soOu+sQblowtqE392s7Fi6BtG+OUUYwsc+41EkrkFGRT8Bxo/jPhZSrnKIBYPXGOQpbpzeavgJpA
8ZzBj6yrUaudLqSkXdnyNiPRZNct7l51PRlw9Ov6zHoB99ayx7xKfHBwOyD0+7XDPz3arycIGPVw
Lmbm1i6ueNyWMr49knPibRarLOS0VMHh6cSnInfcrsrFQvxitERGhDK/h87CspPc9x7djWK0D/BI
SXRCkbV9KrjQ3iINA8m3nCbTjOalLm68t6S9CFFlj8eGTf4vk2qXyvCszI7KJrAme+ls/9tkNHAI
4ofyrUNY1ehylYDCfI56IiQ11epOLwIKqYoQyC27Ddq/TJZyWu/wxi7xdlDJCpOmL2NQPRsvq9M5
8vQlLfywyfP8xIPI1t6vg21dYv1WpzKVGb6I33yXVTozbefNqM608VXRds5xTVdFQcJ4QeK6T99s
MgFX8yUDF6IEzLs9aOpPDZl26G8qsfkzlMbwtCVLyjlXAVTp1NfvQvYEjptBJJW0L7fHw6LadV/V
AXyH1u+ClCGYFFmRAQhOkIx8VVL+f3K1Ns/FJZ6UxwLDYx3bQkDj2L7w14GwCN/Ydx2x6sskALeQ
waTdPtVRYJYkgOuVfE+4kSDNmQRfQbkxY8g5tKcb0Aw+Y2dhPy1qJYrv6tKCnq0jDeKNdkQvfUl1
begLB9Bw55fC+bwxhzi9VlXKj1Pa+1Mhijz/vDGAcGBDaQskWoiNWVdN39Q7vFc6yJpg7Nsg2A0T
XTHzWS5kA2dz08YZUhCuW9f3GrKaGAFx4yiiDiP9HyxFwXWHf7asGhWLwatjoXjv7rysY4TxHox7
Y4mxB4GSs618g8V6VFDsaF2YUG/zw2+XT+AgrJfTnwNPRlJr4jnqBlVffIqUKbQtR/tEZE82xRSQ
q4jIk5s6YZB/HmiSFhPdVNY6cobKc5N18L8YuzZoa2l1MHGZ6tufyg1HhOnxOgBn7agmCNf5JdwB
H/4c1dpHXnRB4OTI4AeecS/I4kKY+a5BSmdi38KSVwjtvQUOH3eo89ppkZbeDStvn/BUo1dS5qH5
iD/hn0LenRfB+LXm91TkAftOMahmJ3r4c+LIRdlC/gAlTXLi37Eq5JZFVemfqlEPphMRN3isWcqp
2SgsGkNAzd0sD5WO8/9NBPfSdoBvKmub5cDN8Vd3dlazeoCvlgq+LKKENfc4KFR5hA1ObvCPmAGX
8H4Zs0qYORtQ2aFqXz0hEzYdhHcLw1INv/Ru/5fIzWTT8VCKHcKeCsOyzfNYzkVldRTVXml5CtBp
wNbLVvtx0Opvy5T+DF0pAw2SgADklyNQiWTQXl0VCo/wR2Z4c/4RyrqHXNRbfFjIInVBYk2Rvfpt
CqGlVQGHVEPhD1mEtYNkaVCLm6wyDdzgT549tIHlYgEDs5J0fG3JMbUeEW+OK/ACgn4h4eyGYyTw
wh/BsyAv+LVb9SpUzOeHOkqngj+KJFXmMbhqmvnAzNA6YqjQy1/1SH0gvwBdzEWQ/P3XrFcK++8g
eBpRFja3zN3oBFGdIsUeum1gnB7WZhwXkf0t4/IKRYsHR6w9fbEOtlNupEIV0AtpcnkTCs6RybJZ
gO2Be2koetbtcklW4Kk92UBPLC+9qCN1dfmKcLq1RYkJUftWdlzK5YmWQew7lajIt3nbWbHi8Ae6
Jn473DlKXCmSB9Z9yQ8UveshzfnNy/Qcrhr3TohMFcnZdAemed1uJlsAjxGij06uPRFWqSOeQX0A
f07WiAc7hJdrIRDzyI53bhi/Zn+cxwgBAU+Bqbz1/mqNiILm0uaRF0fYkDgQg76iOfsHFC3ADst4
Me4HihUEXH/4N5Tm4+01f1u196yvHjH0M4/DxbPFEaS6EozOjp2hEwmXQu/OhW5hocgB9y6fBb22
5O4IQWXMT8P0hpTkry6rzgTum51x3PgyJjBlGz5xcYQ3u2OD3lBQY1OoGDdNd3xt0n0bvHc1c7+5
3ULc/i5lxPBak8EdeQ/Nl7gHyzouQrUqKiP0LDpqfdp1e/w+9V7X92ai3ADAjlWZr8KHMtOuMWkq
oF2El93GeULYe3YinZyZ7zK0G0rGjr/uf4yzo86+RcNS6b60D4ggE6xY2GoolCWG9N0HqgmUHWf/
wm4cU9vXErwjgAwuUUPdUd1QgSrvZ04kDB9150XQtsxSmgJkyQ7ZdvkutXSSi59DEF1EM0j/VMU/
sSYD2SfX/D8KhYWmH589dmkmMD+oNgQuUeRFVTlw/XMxe4Lfw/KF/Zp/73c3VSIwVUESAUV82P+r
OAEDx2NkL9PmJ383P/JxZ7icqZbjTCt/pqkETnaAS0XyN2pfXeOJ81Ryhc5dJjHd1uN6jka/vdIM
DewV0epPUr9oRFQXLtza5lPRz5y0LXc+puVGer2q2DxoQ/cl1dsWQ5lnLqtlDeXZchzJ55TQR8Nv
FZOGHH5RvpR1UJ/1MmHnsQn/Uel9VoErbBYMTQc6kgmKOktb/jJWG6gWnsWdE4b6eSNHdu43E43R
Xc4oW4qxry9oYGkeb7ljNyMqL419piPicmvu9WVASVHOoAodY8Yl3jXVTfnjRk2JU8F2nXrCThv/
zTY1RRASKCnd650BrhxT2LVQa8UmF6v4+BO1L0sqm9gOfgVGSXSpMnPueE/szZ8J/ZnUcbWjZHJo
Uhv8q7gvqUG5o4B/TPDuZW92RnMcXqz2bXrDASUpHQOmih0NyGIf6WvBBPNN6GQaTCj3lyaK8Ppi
3gPf9LfjiXIPAWVQmsfPWLFYGhLMOH+/JfFjxASUD/harpBtffA0gWYfK13j/Npg9usbUol0Aipn
VPe/14aHcOgpx01XeGuO81T8aqv95GENmOuGfAARrKIJFvM4Q8COxUnMO2T8OkKVP7jTB5wo1uID
PJwb6OY2jZtkN0Be7L6X3/3sKQQmoYYGQxhkF1MN/SbVfYeD9S7SLPkemYYIaLKaHZC2HQNYGbTi
4PdjFFbgvPv1m/yL5U81v0rDwjxv0hamdYTnf/qysfGLU+dfFX2s55+KjOyc2obm7d7Oy4FaeT55
hWPteWfEMcyY7hGqf0z5bti9bxT48FN0Ym8Iv6MEDX3Cxnv/zOPjdYBN+GFtEmVWQnRqtjdL2Bz6
y3eiRnerQEGjKZNcdEgflGzRSSzMDNAC2LQLVfzkBMjuRVwg2nhGaWOvIvgvmJ0WIvnh5J3eRWqb
XI2/AKvYOaC20m+tct6HTX/0NLg+4SKx1N8XYMt4yDtQekGclTrLV8pR3nRcmCivUq5GjD47t7cy
ZUtKjuzaIfeVthcueIbiQhkJwiroJsotzTieUXB4vdKIaJ79Yf9UAPAyMp2ZRCsjR+cZmIn068Bi
PfYKJCGviXUuvIsr5JN6F2OSwpxJZ2mWWMBVttSSWByVgwk/s12l8Eyj4yMColAtCbqkqVWSr9NK
5DkumpbnfVtWS/UXFSke2h/cRjLONzB+ZQkGbVy9m6n+KwCSB+BuZrj1sWU7OLYroKRdFTYsWOMD
IG865Do7X4tjIrLg9FyvdmdNVxpOIO9+EQcbotsmn11pHXJEunPkxnY/uw/jlaLF5ELgebuOhH5E
7ZfPyVwJeQtMaQIdFZi30/DVkEQXTW22Z7dRjyCZFub0xwfhxcKwwzuRzHRFUwoS1rvjeFmms+eO
WhVwgL5gipfEeL3bqv0urCyjJ8bE0JFq6+NspKV0iMM3TtVyPPteg1L6Mzheul5RxXHUw9Xrv8R7
A4oW2vufXIt21/pvlMV0H/qYiUrJDwOIWjDxfecjo4dhviWJ16RZBlBlUUS0mOrn9GDQE/kYXow2
Jg1ZF36nNQKREMg+gDULDI+eUe74NY6IgL0Hrhm+Ye3zFQGFhb0clyqqwzIQwJOmzQPPShx36POf
T1UeOz36LYF/M+3ZMYeoyBhx1h1VmZd8kbKhrjNbJAqjCFAND0n+DzMsTTlXiGejgpdyK6yniFqM
3EqAoKgLdywwVH21aqj/F1wcgB0pnZqB1j0G2MJlsCmqyp9HF4jKEdMfFCXYGyY9WQE89uXkrFk3
VKSZ2X6DdsHGDNvrDLQrSahdvqje1go5DlU0ymDJRSUAQ8hvj368C3OdnkMSGEiiOp1lWXEW5Zh1
ylLSOuczLKKChGRJFPTK1ApvcXC7jMVwN34Z30BFER9CEU3nW1MaxnQgtn3EsCA6Xuai+5svQ8xu
+CpTUY9WGmHow3dp6/Pm05RMwH4xNLCyHq9ByQQYJHjGryp0sSKoTZt4AIG7XrY3Uadb6vKWItnD
UcAwsfigEFgRJbaByHUu027bi9QhDBcr0Em+90RUaTzi3z7cnmRBl0cm6xUddyXgKyKEupD7grB+
24PKdu/dmM4Gp3zK7Chqyi3pQ/7tT5coWkku17JzHXVw3+dDUt5Ty8ToM/jFyP+CEzVap2jMYDLw
0RVzpnJjGwvFDIYE6nrIks2fZlaTBjU/+5nPP6z2uHZA0YnIWIkX6MZW/R+UN7ZyDWnuj4fPGG+M
nuC3N6lkAoALUWcyeCk+TjbbL4lACbjCUCGw2jTKhz+dsPg5JrjVR/ZuUhXdWgOusteihnuBtklA
fQg2WFvIpRKeDLPbq17KJ74nt8Lsi6pyo4GpYHcWExsDAstFuzJgMcM1W85ZU/b/Lla02cTUgnak
kekWBuxYMyiRqzdmXhZHgH/7i02+7dqlEFVvQI0xT28m2F5EX4rfo/RDKkubCftcMJ9g6YgavvxJ
J1pdh9dsAYUcGCgZMNeZsHAziA+usUTllY5h7JrVg6UshX63B9UnVfz/SRzeeXczoDtEqxQqb0Eg
6qiwUcAIs3whN+AsKAgb7QJPpcYoLbbUPSdbnsZ4Ckr+BuXUknKRv8lSCtQ4Ir4gwG1smuArmTS8
dAEulng3F4o68X6MB7gLPwN7EJZc1q6w+PaJdqDjHkkWe9eUUeS/JZ0VfL+JD/wixDIUDR2LUW7u
QstQ6BaXzCM0NMBOj8sH465DOUESWcg3MS7G9MIHFnRUKoGGuHPgyy/OxBzuGNispaWTs/CiEQ+j
FUUna48RsyaVvppXc3pEv3eHOlK1WJQJWF6j4Pc8g+qk1uYi6OWNqZtwSLj3F8e7o1g1RY+eAAog
DZOa5ZNL/44kQDGuR9X6pdyRBw7JgPspu9lGMq0WLgLen6ZoC2Wkqg+/6Tvezy7uD4Ho4wIgQm1f
IWvd9zFygM2NeUisoduNbcxnCu/KABZymtyaYH95b1TJoxs8iRAFSLhoOQMZx5WDdhd0OcB692ze
lnhSnR7XYBWB4G4XGr3nVjb0XPyBap5LzFcURd2aBhndm+kfHt0P7sO7GM2gvvLEEM5hQ/nwCReH
I7mTq16tyOREFvWJ+E0IpwfMOlHZVH6OrX73DSOgNMOKYhbZEB/k7qBXaOVVn/L9ED3hXEbTqQB3
xxRzDQqnfRMMGnXbwmDIfKJkzeEda9+ubp0Fm17v96RbEmCVHSqGgAWnEwOCzbFQCKg04/xLg9+K
wihB08c8XLq9EeMXqVueIoC7/JLa+v4klUzLThFimAw8tj2wZqv3B1lhMI99zQMbRTALlGChQr6B
7d7WozQtvIq/9HWKkJzZkQ9wAs6Bh5CygFLLvAeHdvugBsGTKUYGp/GYD8pXrW7h9TWgDcNxh7RA
tqcZBEsHH1JsAogAhBfWMKuBFaT12PKuF6kiG+Kd1rEXknqKemT8L0slxHP2JYh8xEc6CB3JY1Yb
Q2Ea/0Dqb7di8YkGh3f7uzbXxHL8UCVSSG+qWoLCxjcbO+idGGkBOI/W02cbsvqRNmZQGZAq0h62
ivUKsY00BvW0is8YS/ZW0krVMAf2yRuV2yDaJ9AdyuFUTtqlrCs4kCVdJwW6DWcbVHN8Dc4xsN1q
UUO6BH+ne3ZL7QyNdqltFui7d/WBhuOSepOR0pD7xyGtTup7iEr0++gPWrXGyjnP1zAWiQpYZOmO
HVjku9fOKKi2fitGhDJ0DEcZcj/CCQhuv0r1ImLMTDzBX31ccNTRWNUyKO2bWDEcV2uEv7EwmUsy
PepU50O9Cl4FUhYWwZvgHxJ89gPoGHTzFm9hseL9moBVk1Egke3J5ISDYVAHtarjyYICJ5EqLJJX
oAQQqKwo9WJiTOQx7SET3mu0ktqbRnbq5eFsxi1+igxClsGHwUFfWLoY0LpTNaMAbs8HyvXCsipv
z7rZo1aOWmDqaB2B4XTFDSguYB6prgKu5kMl3ulq5rbsjOmk1Vf7cL857lwYR7dwzDcXxxPXz8hQ
EiUa7XnkXVvB0k4iXyJsfvCBGKRN66lufIWhp9yU8kL66zl6rVjvvYL15LP9aCgbyFRH2XKEodt1
M80oAqzZ3iw+augS3qfT5ycWva0yo8X3/Xbp5QzlC9DpSjNDTudTeTYk5sDpObsahlgzv34mhugP
IBmO4qhevzf96ZNlJlAHINOaneX5ZzuZ6O8/ewqHmWOqG8cr74htUs+Lo/R0vm2oLwCc9TWhnZbj
eLXWCOs4MoeX36Lpe78neT35AKEO2wYKeTectpAdx2+5xaCSr26lm8ov1kkZxOcToMNK8hO6e+TM
oZXT4pnR4kaic9eQ3a2fEiZpIYHBRaTk3TRWh+ijfQHDXGEiqGqGXqaFPH1ULsjBrnemARueV0Ps
BS6VF4ijAkNmCAKdFwFZd/yUctaHFEgx60lWAQFzV6PYSHxBebKsG/HHzmgjSkWhQ3Oie5kGsQM9
41NCa/pDGZLbvJwkNFCRalEmAlT36atHfLKToBA5LotIRtrfkVVYvzUq5pBSDCZ9CTRGaAx5D4C3
9p9bOUTyXcgMHd9sJqla2/C0sSIYPzFMyn/t1uvH1aZyPaU804Prklj6AfKvoNdOCMMi3Q3LvLXU
8FImnIYkCDRGw2GaVdQS2eh5a7znHLQtCnEWfKfRZEdBkzOW6hCg7iIy8UR2LgMRDmUoB/9Y3Lzv
8yTu/mT8/RKwN6B+Ab5G/TxjtFUXn3He0X6QSjRpfCm+p2ccswPXlUptl3bGGUQ2yHNdJJrxvtls
DLxLGEcSu07SdL4+T43q60qTrHfTF9M1jqYbklYpYObui4DMHv1Di75h/jHRLHGR01tdoupQCoST
jdH1ekVyItLWspDdrErBtRe49z2M754YXJBq02Tatga49zTxLjOMT1kh4a+I3it11FMXxuEo5hM8
KpDAWOqR98MbF5nygK6Q7D6zmX5EJcAeLCgQicdP7r+r5AnDvwllXCjMkbY3ZeBgk7a3bemaPMjj
xEF9E2SU51L9gODOi5S2+BRMiBvCxhr16voUKnvL6oh3X1ANgEdhhwEF6nFsqmzTYFsGjncnSZIj
xQk/E9pZZGtjnkGaPWYkSEu0bGUI6AD2D+XVBm+5HuEiJO9mZrWW0f5KPx4eVJJ3aP3SvKP4zrEc
mzk0O5jGo5h4tUIDxlppsZtbChxlkTF8i4Joeb1vCTMNIudPDjxB+Y4qKSDaAVOCzy06omMlDWrz
I4XNK8vRehPKZbW4peCshUq+l9NEwFwGVj0BahXIb2kmUgv2J7anMnJoYIKzmNjbXUf03+3zgBmN
kCUozJtTone6dv9IoilMorNd0Qj9jN02CK7HEgNt5ivZPZPKxgKqA/8UpqqHBYdn+VC4EEc1oEH6
T8//2zJU0B9crpwqJy60/91BcgK958so48hD9QphpPhLFdH5wo9QqQWL7SpM/SpcnyA9SxCjk8yt
K2rrwdhy2/TARlNsFc5acQrTWN6UkB019WM4gh4lSxqfLGSATmShczpPto30R1dg/325hlCLg+Nk
ucOJQtW06dld47f+QrsloX2sjXpNJfoil9V9wwciI7s6vXwrO3VvWLB/PFRCZmEUJWanueh8SIw9
wQMU8+N2R18AIKTvC9QJV2/AycqcCgQAo+RKRrUEprGNI7hP6EHBk0OYSiMj/bEGIqHA0vhUxHiU
347IgHv6rj80XVQcP+6JJ47jjjIFfqR0S1d3ior5+D+mIS8v44wMBinjn3r6W6L1FdJnDqKhcdrI
awC1N16DwuziXAPub5Q54YmvvKWjLoYrgk8UQ2+S8OL+2wf4PHAlZN5rl/meKg/wXzcuzK6eNLiN
rrI8eK5L5T5dpC6cUqlVyda3+e8cBcCSd5h1gJLAdum07IxRdlGmnLEcrThES1LRblXelRmgEba8
2Qjyk7J9OvaOhrm/G6fqJnY9GfWW+93K6jcOkTcbJSQAU4NE9kQicjj14kQVfraJUTxNh6sn510d
jKOveiFHpL1wqHIZdyrdNKUnfUDHYrkVnpZQPwI/3gXhAK/6VCNTv/cgi2cq1xzdR6QK5KmDus9X
yfLBru7FCdHHKt3ZWnz0yjsuQFzOi0eVW7CghrdTXqChiO9pPyObpN1arApXHTImMfDtrSkulQjU
isXfMsj+ovEkeYdunGSk6ZG+LsNGHr6qfGoCa1JIMJ8fzUXCmc1uW+K37q+nj4eXT0SR9waHSBkV
m57SAkZ+8gsk8jeLuvDU7UHei6dWT5RamDwDNQhljKexMxZsoIEgiixzCF6RIzPKAPsbEg4pX3vt
ak3RcUKFGs+GL+QdRd9tddcyJjCfGUw9r6G+ZymMixbrlzFLr3TGsOTp80EtbyQ7mo2qhE4ec7O2
QYkJOznXWvXVrq+VMj0b4qi3ztCM6U1TloHaZKRmuu9g6d0nzmyu4KK7fEg7CYGgekokVg9P4Ss+
ed10rnjFF7fAj0dP5tqbfC5ArSQ4PPaUr+7dqnrzCM8PSLXqYeQaB96e6uTmsWz9seF4JqtFMCco
/Pg6pz6DsxqS7rNCyWJ3WKbo56fGVitrjKZ19SdFtVTPHRlQlid+bR1+dOU5QUfgfS4bSfpCbPsX
xrvnLwty18NTEc22lEuGbubmkC9Y1zHPaeNfVxFLRzfNyhznRMlVhTmnN0FtQaBlKvhbOwqSge4Y
thHPgHVVykn3K2YFjwmcutFCmrmSQDIbOfdLp22iRLYWTfSzWakVwQ/Sstqrj+3BlUIC9diqF4O0
UR/hNLaoDTq0E6n+jtjqkNV+0n6g39RcZhdhmxRok2yzXk4xvl2jCY0I5Z7VS9FnpHgkBdu0WnM/
5kOWbCevRZGMEwALCNoQzYUkXJWHnLRTPmeAmLArL7w0Hzs+KJXBeDC2RTomZCBVH+Bs4XHClWwU
DP2cVna8G5CAZD4hsfHIWVdmhWPsorYSz5MbBRIikwCCdUYh2B7f/UOlJpMCS9He/8UYx1QxjqRr
Qp1b5q3ScW8vAybolqkjOxI+lpm6Wn33EO0xltbSvy3OkL2X0smAr/C4HjCNrcODG5oD8Lv4gjFE
OSFxKHDEtq3M7Lz3fYDWLqOuGoMkZDB1V5X4Or0Iz/q0jMqGVfC0WHejWaG4ALjOnIC9wqVRim1x
ROgA0ahkfAybB8De4T82IsdwyniCNPDL0nRJ3XiAq4mAdaFc3jrtHvosZDTyPNlX+Rf6djW1hV/u
HbPjpiBv1RESDWlvDWZpKzwCuwl8vn/CbbyTViiOjWKTqU3UlSqGGd4tTvVaKdGIyxzpMfjypgbw
aMwWgHYZ93niYEAYtzSL/ZGwDZhH7gQ9UaZdksStyFyZGGkpyWAUv1OFmB2t256UemoJHMBJ/wUI
Q6PaMuyUEdDcUyz6/5kNvGiwEzIDgF0N1VpqWvNrXaTis07nFUmsYTyzi/3chTOFIGvMxD94qs/8
+P1LRitt4BML6LKfxgSHROxLtG+0E83zwx5eEhR76fMHCVIZadkjakHSZ0LG+PhRAKGs88+dcX0x
yjVRZhT7qXyzmfqbd/9hodvdFcRBJEq/u5p0MBsTfUpytK615P2m7jKJXSdMpe/kFmgjpZFJHNfc
AxKmKwBShpa0Rw9t2DEFHR8Fc6YSc+nve6Yya9J2y6ptxezff3CkGSmlqEr2UvVZfPtxOA+avPcV
WzWItrcDwVCUPT6YohlfMuy0h0yUSuLFYPRwx44XEWxGv37fkBl+AevPH6cDH8gqJ+61IegSm+Ar
x9Hdphr5SYx1qkAGFYZPk4Upewr71oxjYMN6DJf2zMU7qqfvcixoqSjb3zXeFXS5BDi3ujlTOzbA
gttlMmJtemw0j9EYt3+StlUOSLPwEy6BELR54IiGeceNi/iAFXoC3jBBZxKWmmJiUyEytt5DsViX
QDQxCKgouFEWhCNPtRX4sIk7pkYHrnxQaYxGA43r1eUe3pk8pIItYSlWw6txTHUi7Ki7Y+ecdGpJ
tXj+10UztjXBNTv3Z9q2QBvr2WlpWZbBXW8JIJHfOzj3T8PtYoNaYI2qZaVmruTv5R4L6IqYh/jv
JWtXT//W9lVYStX0IBXRZxzt55VjmS2ogFyRmtSca8OS2S+nQNR4CNK23+XDofHN4J0eb3d3I8r8
2XLwajGcG6dWo9PYBBdJ0AM4OEwHdAM1qn124kdy9KgLXevdTwlPwiH4cfsd18sjwl0I0cBqssUo
c5N2bxW3xjdi28LqhbnWwD+LI78NwhCgX6md8lSjXn9xdj9zvdMgPniC7tfj5CEzaYHD5lU5AOgO
kYCk6pu8VwY4aF9bSVbe6Bensrww8k184i16Q5UtIpu55/k7LB3tnBC4Y5SIyPrUglkzO0PpFrHQ
24oAAUjOHydZWtVcTEjw+eRsXWHQ/TLs/h2mLahCl4oIeEDad4lrQwQC1iK90cXUZ+aBPxVs9Trq
R88VfeBis615T5y7vAvbJuXRVMStGpcqc4XEGqS2L92wc7yYIJw8BZ4vDM7OEU0aXqFqj86TeB34
PslZFPZ5doOR7lW0qBa5mUPtHMJfV9M5sKDgDoBPW9Qg8NVFoDEy827lmUCUq8cNV03xu7X511IU
pucwbXZUR1iws7yf4OKey7DZRJZ8ZMc2BTa0uSP4Yf0VvTGkCDsT7q7EW10zi3BhwPRwFo46BC8i
Itbxh+kj2xUkctqxSG/B49cGGY16j1FFbbz/2OTy2TWs+kFkSFCzA0p3n84CUcIleChvOFpH4Mu2
ykd1wHb0pvXXZAa0Tk+m9NDtxW+QbMA8trLvAxw/zzb+VitDD0p/eQqYmpdYUkMCph2+y04ooYgv
cx7SM87zhlv1fSiHnbuE1CjTq0/szVr3RylWztyZ08+LOqQeyEKbsH/EIivc9IZRVzT/BVJgB/Y6
zVlSFgmx1L2SZoBFO8cWnWRt+cMdfvhYRDQWLNBxg5XIHpBVaDitnlfKO48wSApAnUwm3mC+MQgQ
yqSOsFDK77Rd4knEeWkdj9lEtGRegXTB7ts6XXAif8ObrVCvjISwuLrVjySRVqi3MFOHcH0b1nYI
5HdJiN1Kyz343H/nZ9xDcE+9R9o+GoLMP9VT9UCot2/EVxKPJTXs+8WvQwlQ15pabXxaUEiVXWXD
cIKGeU/rahCtfvJSNC3zhc79toKz37K9Nf5CCagapygh90pq+vsAHWtafz3v56yGBzHCZQj/EIvs
tVLBk8rHjM0Jt7eFgXIOfeNRrYOGMAI5c3bStehg/esebmHesu68li6t+RPpPdNXEs4gk0e0iles
tvpJVx9w24G0b9Zrk6LsX81v2RVU3BmU/+j1khGlb7k8Ke2Os/VWdfpw1VuFYONIIabZ4ZwLHu43
+lbMkWe1e0UC2UQoo/VWPVn9mr25AzUG3J9eOxfrv10QuI1Zp3iHlFKfZNhK9OeReCxNj02UEAGS
IZHVGJau6NahULwBAjQOWif3xbX/dz9TF2E6HVpr4UrEOuo8JEdWDDQ55Uckm0t5nmC/Tsm2CXwz
8oULR7gAJIBPUgoqXHRhX3+FT+e9LAk7D/oOeFJe+bAnFV27cvmXHnx40qDozTtOrItVwD4ES6Mo
VZP+cTl/nTuWvJvbP/SBaC988w8Rxau46Jex8dETlF0JWtDEBhQ/UXQhHlo2Xi8SCSeC3cIV2pKt
tT5mtodjPjhzrhaimRMgoddB8a0MW89S/N/QGKg4jCb2pJZt8C1q3Z3CGjWZRX4MXjcw1yPo9Iur
jnVkGvojfMpboAwPQ1indZDoU/2Vpaqw0gQAGv68V5y28splunDzLcvSUaSt15cCylJumYoKv0Qw
AWeYwiTX8L9ZUhMMky+W8yaIH6M8QqjS+lllXfwdMr9siurFyBSAZBBvFzzsxigfian+YVoSDNw0
Qd+z1GyQ8Hj4jq+4b0QJL67ZXuEA7GoB08nfouqX9rn+c/GPdC1+AB8F3kVPfX2bX6pidG/J2VNc
GJuvyFXbLcK4FmufXHaIgKBbIXVUJ9J07GUFO7rdlpkJHeta/JxcswVVg68p7ZPBCgYIA1TF+Uaa
AfKlIXPrwNsltQIxcB/dBspgYLGuajg/vl9X+QRlkFkyIyTWQ/vn9+uSwlDrOO717boe1DcGeKkL
Ab0Dcg+l1LrSXVmoGH7GsSWpMF1ODfhALGu7mFVucd4P35KYxGc5cMgYhvoBT/cFUOWWmbGty+PI
qxvND6EbeJHoxmLs++rYVNlEFLz7+EQO9iWRj0woqB8TLz1CuWlc2sW/3S6bfJ+lJirjdmkAmRfG
6M6NFnmmBZnwm8bqo278+/UANUwuXKKAqc81pRrOAJAuNQ3lKMup3budWZ0hs50su5mixifVjQNu
gkez4N/81XXsxWbxZLUFfedyYEAOdezRQrcnled0EiKBS8GWTNNCqzzeT3Ohq5SCwTtLq0Vv31Dm
9G5aoTgwXwhzygiaSs8Sm6U7QV10eRVe+1AaBB3IDFrenKGOKQg1z32b0Rt2qHXMqw8JVa/2gMZr
Og5XbHwzx6/TevipkpE8MG+H5WHmCvX56xce/ivorGmGBzWjXUHDWeEDZ3gqa3PCR4KeWzYL7OOX
VdbnY8weSJQYSJkDetUKjnIF3fwaBUGw+TbLAstUpd5Dw2+0wqX+NsQ9VSqIppAd+6BNjA1a6uFt
KTf4bRKQj6eaQ/ek2Z1HJw4+Ead1W9+NqhYoyg9t9xXLo1MFyFatI6xXIUDb43MHwlzhY9nMJ3FP
p0gozBezQgEJzfLVaDgGyqL2jyJoXIGQ2g+wBwZfVZ4U6Q7TgDCi2XzpUCpfTWgp8TChSXJTFG4f
k0+fqsnvGm5MVqII+gXyWFL7gdpKzIdaOvLfqcJiwEZ56IMqHfm7FHJJI5gseXaZcZu8jBDAylQE
iMsdMO7wiUTJV6mLs4jmu3SxVsKO2wJkTqT2ug9skZ2JzCBM/zUOKhn3dZAPeLCJ8MiEdBNGGimU
/5HnBP+xmkXY4fREROxVGnz3GPh6GXWucp8H1JZb8qqpbLrGfJBCLRGwaP/zzKeo+Gh9KHsYx75X
/FXFoDOZ25zxqafAwXjoEnRTkr9G3QwqsVZuSU4KujAuTDTrRg5kbobn2oNQTu7iO2ArJTOHTrYc
2aBrsqh+FPH29gg6cz4mFbQF5m+938nit9iog+mKS+M4Sa/HNGAg+d8cvCctX/oNfp1DarDU4Uty
wMUFE3z3rkbHyConXY9UHiX3Cw4/wH90xAHNlIhlvoYyCLoa0HuZpA614E7HrBOVDrYV4ZMWKFxw
92YBatTjl9HZSjULy8GSeGP8MDqDwzMpMIkSgRCodgbrR+KYEGdiZ4NYXswm5t4ShV1+j8nfeU6I
CIeaIy97KNSh6NRTN9FBkykGM5iy4C+fwiTpDV5iOtjh1io4iITIhqtlFxBpgwpGNfc8QZT/LF+U
yTie2XCX8tUpKF2b/ksoo1eRQHG3VD9VKfoa++rs9VkE8r+JXaf0uxACpqrR4hhc93VGr3B15yYY
e37Jhn2KAb7vrGHWtqF2AnadK7HyjyrswO/Q3cO4WQja2Y20EET20oHu5cIUJkzZGQnU6e0v2+vE
USJsL7AtNBq6h4jawDVo6htGesDSG+H+Nrv2sInz0zLZM7lU4mqbL1kBKXoIqGOezuBFRx6S6Iy3
8JuKpgWNPksEVcJIAPJNOC6K3sUZDcbGkaNkXL1EaW2sEwYc24RPEmPs2kYUDypNkXrmnbl6NLjx
o6aQ5VCn961vHprncFTCna20MAAx8ddBWhkl6X3vTK7ZKZid4F1xrO/3fESsloMVFv1aQqj1Y0Dv
IhARyJpQfI9brcYS1QG5zgjJSvfboAWlVDrgGLYlBQ8qVBQOZrZlrReOhAFY8FqN8zj6ovGSvp+/
zdpe7PB/cWV0ejHKnTPH0UVRw24oYcHsyLAjgRC0Gn1iM8oxNDw8/WU+cKQuSPS0HRBMo9r/GgVC
GHACf9OaZuALW4whEWyh/ygJop6W2GsHV9fz4gW+K5cJY3mxmMtTTRPONhrRPRNj3ymtZpfs3fsl
125uawBbzmJFVMqdS6LpLA4hawIyeg+AvJHor1yXDCY9xhTdGZO7s1WqgmPFMkE2KZexa9scH4fu
KaCEasH8XHA1KNDZDBpxA0//5925RkpDzxHSOTIKOY8pHbc6QETc3Q9JZwbMOEgegC0CgQWqB2Jd
L7ocktHVmrOAPPGWOn6i7LpP7Uk62L9Ei/LnPUmoyTXX2o+tfvplZpOvYXd9++kBWzzkjcIx8ktb
NiaFPFo8KZ89BjNf938EGWRpiubOnB3IuVCsjpmikSZL3V2RzN+n4CtBLo2WnJ44O/jCYMcpIFX5
wBE2898yx3etYl2IqSBPQD1ANTFWAx6d04A7MSzo5JmlXVZl0g9rW6PXfR08UIsGOrrJouLGt5Yf
uL7FDw39PrMutgmpVCoa6zdenxMg5eYOTH61hEVZ0y7qE2f8X4ClRKZb61YexKirrId1YBHoUi5r
ejdvpronEwLPp4oCf2y/piX3ShJH3stz77fDJEUfJRcFYYeRZmen2SEdPVoBHRCRvcvjvayJUPXo
qyXZAVSNJXY34xQEvEGe2pvZcvOe2JDEmVSYSMZI5XHe+yj95gtO6Nfvktyj+QKxycOnsWAfy46I
IZzHttv4gGWTNFR6ko08MxVxOfF7iOpFgD5KR4DDajqnU9L5+fuljcgmlrRj3freimSVpaSNf8DS
bMplD0/yEqjLLMb2Y/zPN/wIur1kV03ux5PKes5i3nE/KnIisI7lCfyq89hz3uy+t+AERSjp29TR
6TmdU4T0ErLze2XTbIV5cYcfU/WR2S5TzeTVTPWmycztVOgCf/CwjhKW/6ngtHj5ecjEEuOrw0tE
herGeH2u63vi3L/Iw/5rBzk9aj4QgaDcKRUHavumErnm70qetSpgB088CNkM20uHIt84KQtoOxGl
0LGVWZVQlX23UXZE1Tya5WrPZsZ+aAgUXl5lxtQyhQk9te/lC9LJfyOFv/nhUACUWE5+A1fFurRe
uzLzwkQMgyJ6vyF0YHn1w/xe/6JDwg0uJLSH0t3nbRJEs47TD0FpPgwH8cimwr3ntlekoUPWKpiB
WdB34b+beIpxRpXWbMpd5RLYwXy5ykmrP2D/jCpy/v0jaPyviolqoJ6u84FE4wCEW44qmuathYaX
EhqJHTHPbptWYFwVzC8RxlOt9wECSpsI8N4KzjnqkRVH46C8FIIRdlpSz+wcGbL7M0zNuLDN8sbp
g48i9tEFoANh83uL7XNnBrVIsI4vN5udPYHmqXffRlIsu4biaU1vQTLtKlXSXGnUEZGoL3bACagD
t4r4fdwZzVm+3xrcDCwTNpLA8lDeG6y8NZh4jceWcpOt3UysHvLIMS4Rn5vu8fzE1YLpVOXfqoIa
3A5ArbpU37UrUz+RwqHLzWnEjG6LXvNClF7M++ctLsn3hyMCLVwoClX0aVH+wv10oskb2CyI9/P3
Lc9Pnkoebo4N1LDV7KolXGlmhNF9g65CAfkwh6GS1nl7VwUb5oot6A2wDFOc2G4cpDoJU8AR+p0c
9vTyi6BS0OxYvQB0O/vLfotp6vA45wdD/3QqpFalxJ8qvivcMtNT0eqwvXKqqje+2xBvGjTGTrm1
d5cFPi8YO9vyLRIpsxNQpcs473DzkbwjohjEIRirEhE1gnlK6/gjjPgWmMC8km6ZRPxWFNnpanGr
Usj2wEHHEJKv6p5HJdwMkiOgmHmeVDNjpbNjtX52dQ45NfzeX5TAdOIntKzGv0J9qSgXpV99u6rJ
uiLa4d5FVPAjxooA7B9+FRy1c/al++XyNieTid0w7+h3NdtE6bK26r+XfR5vX1UOiMSvz/6vnokb
pYPmbMSbzEF+gSEyYrOgt2yYLvGLhOuspfavVGlyH7BTI9xPla2tK1YzP561Btx3tbxMzXLx8xSk
hRDjtP5hmSO9aLJsIPhf324F4t8I8ONFkshZA92vRlnI/OksW8f2ryqvIh04+q3jXWg7z5FMRfRe
iTZp9UlAs8Mvi/G+2tukGnW+6/MzWRCoU01vrzZgrZ3vUTLstYLfhbboRj8wrtb/0OGewC+R19TM
sXYTH1ikR+ITc/achJAWE4LpAIWH9AykAoF7r8mIKRBQRc11AX4cPfR89WDfNieOoOPyFqt6XTrE
X454JmrYDyt3GvbOdhqL9s0Yv0Z5sxD1Asu+uk/QCKVJXAq0bscUvW2OQYcoi56XVcH00Ac7KBg3
9PHhili9YNk7XafX5AZeKkxpfSfClOw7mpPNqIObiHKZy3REVw/DNvzlw4nVUmcOc183oAy/aAdE
RgRp1a1btPweG/NQ9Y3rDDcfPA3ubfEtiYDuRYWNduTGBg8e/XMwTu9IETafP2pIH1wPantjgEUr
DWiKg0FW92N7Z/vSG/nELy2znnLH1oZEfcGNiuOruIAr+x8sI78oA6YqExK2hmeO+Wtx/PGxrXwP
ZNe3QYTunvKppM3vuPjJf7sbbD9gIEQphz+IGWZAyEJ9lmF7zJ7eONr4Zxm/oGrHfxY2lkR9c0P2
WgtZjCrEkX3w1HsR+HIuH8T54ds1UyA8Jzj378OVl7eARYPPJE8LxCNcB7KzE+Be+uJN5LWhpwDy
BzyuirJW2UCl880NOCCq5QHujyHH7OF6yJUw44Ud0OEF/ZzSrIYSl4IpPVcPbfP3uxSijH0bSa8E
tWWK+jBt8Fs3oeYMSqNPuDz7ULUjYxeH86WX8sO+Tk3wjUeScsUUUZ0gehz6PphvXdoiBVm2vEEN
OYe95yqNjyHHODxeYvsE55ZwGBgbuXtXpfcV6YPjPcNX1fWLwF7nzqmpXnmD0C6HXUdCffWSd0M9
BtbxipFz3VYiPRa4STuWWWCVd8GTIlRr9aXdVtr4+1MDoFXtt5npkCAVyn/NrSbgWcZELlYMSwmx
5qHZ2FmZQLB9PG9WSEtiw5VGDtMVMjeO7FMoj/rIgVh3P9GxcDsWRdhnt2TQH7j03GPhkeRdQwO5
iHUNJHRfdE51DYrRVbCdcRyWqkzjQuarg84/UPovD8fBJcBwibcatx8nsQQzfJjUBQJc3U8ijmjt
FW5cqLab0CtlmTUHpH3IAtFV7OQ+dNYPn22y3eAHCV/kpfks5bTq8wUnDPjsoPs0Wwp98zbvtRuy
GHnw7WSXQ0gFYNomiynr0znl3/ickjT9YvgYa41QXxkgaIFbjkbwlOuhLMrOBuWJ5gSfG758AShf
Q2uXbPiUL4ZQ/UnXmZorlFGOHTnhR4so58jSX1+Gzfk7kE72TWnGD/t563dBUiRB7w6OZll58LZO
CZ7Bx2E34OHYEJ0X3q6HkeBQly+Bx8vP/aM1QocY1SZpcL3ct9Odj+rZeD74K1Sb41sxpKhbH087
3CBnt4UEaemmIm2bV/x/uB87glASDga/k1DrcANxGcELrdDDMYjs+3sPKKWyEdynGZ6SvnFK96oa
2woFpvsSWKeiIF+a/RwXOl3Nk5/xrLpW6K493AlODg+FIM0BdoMEfOw3WRDYoYGm6qB7fc5I8r2t
vhOPsxPZNmG0Vaywucldu8hebTWN10m+w6T7DIjrkbXLS4aFhke9VznUoey984A4gf1iN0hO76hS
2+lG+A8/L2a2ReERhvC8A4YncacNzT6eT+p67xH7CxRgzL8xMPQTFdd1rnlY9m7Yp4Ilo0nHYx3b
Y1ZxdpVFc6bSIMVXomEFXAy99BZHNlLQOwdZQ0TrZ2YOBg3TcyvOSeU6u/1KJmGR/eLCcxOxjZ2E
HRFwcIsXzaCuJkOHDgsW2ziUEXFEofbaaUwv+eg9Fbzhjf8zpxvx3nEEfKZw9tkwnWxUiP5HmZVH
gMwycJ2BNoh60xtq5TwFVcCJpOQunTNTZUD684pa8scXLJknsiV7puEHFfJ1xtvOneArzp5tVjp4
9knsf5Bl7Y8lFrxMkJMdHfTR6+BtQIgOUVn6Pxip4idv91EZE41P0yJXFZbHMUtBOTbD/hCNpmZq
r4s7POqpaK6BXkigcGMgte7TTXk8eGvTAvPKLiPrpq6g9tU36uelo21bYvsiPMwiICmDT33az7VG
SgzXi+UiUznie4DfHi37AdeXtjdz1YrQCjo+VyqUnxqmFhH1b8DM0FOEDCPSUl52iD5jcYVsEUtu
4+m++Ja2yve1L+L3R/6cFVTmsXC6I2TOhputkHCd6++Dcswsl7B+9ynhxvOXc9a8JQ9VGQeghdDE
e7fOJbBX01qDjd+alN383gB2S5bBOUI+snYyLhV7bD4xd3k1mSrr+z2/dNYFpW6MCtek0w+shorm
lLa0CG9DjNAY6q6b8tqYmQZxDaWrjrznuyI/z8x4LybonZ4GVMSF2ygSan8/AGNDf+0o0boGNlLG
i4SugFRMlu+WEwLD4IF17oRcOxoVn1eiAJhn0oZm+yfNZRRTrUDS8ti1Q8dtS9UbygpdxgJHKU2A
FOf6xpadZcdx3uKuUaTjkj1WEBdvjCrBuT3p6CHlwXUXWhIOLqaEtye66AJ0+xrTXOb+iLcwKbmg
2pc8kKzz06EXlpVv2ZGZYgADMz+i888rPd0Dy5IPk08iu+fj2mfEuyqYnpMteU1HtlQmI4oYyIPa
2k8wjWUUiXw4JLPXAqAd6k2WLD1uVKj5B6FUU+ecv8c6psHv3LaY6gBVHDqvtHkbUydBIwIA4PuA
WV8VKhtFJAS+D+zEXg6F0NCNQGIu4LbJq+73H5b7wIhhEPfPeAxgMGbsLQgTcZvX/nTuq9GDZlvO
0Dm6zWoScNZRBtdmUmV7/KB4WmDwiTah1R4blTOicnqwO4grPt0KtJvsmhK3ez92KYh6qVlMckQ1
KPOrgIWvRyxhufjziDj8GU0+U/nRK1hr7H2CXBNfcquAjbgJ1/TKCd54hUMUk4yQ2X1c7+fbk0sH
c82G7KlwMEXTLH+uLVCOic3qOx+wBQtYoDirIQpQ6tfNP9wl4xysrWy4UFVEd2YxiZ2lJm0ihHLv
ISI1UarKR6iiTSVQYNS3gXOSdO5vsRHTOvFy6d/EgBYoLCnmBbvsLHBUWoZaczTIn2To3L1RmCg4
v0igXGlKucpEA2R97Xo5kC1xrGFpIYkg2gxPguLfZi0IzWv/pwzIK1Wfhcfge100T5U6NuxwVQ48
WNrEVXnrwuV7NH6j8/LLnpev07G7vuwOMcaXxRvRxRY9XeKpZCrxqDdQlr4k03MOl6CcXZwCNOfP
pDz0GyppwA5NIX3A3adCLHXXvpl6PUf+L1V64ZFCb+c/bnRrOymU8DE22B1a9+QS9b8sYsHj63EK
unwAsmZ8Wdxn7Xz67Dnw2Vk4+pb7b5O6Eer9fDOQssJ5ZXI9lQONVoa5t2ahKfTbvVjb4MBsswSZ
UFS56ssNnJGmg0C3uMheLx8oCujj/NO3K3sU7fxJCCr1DnjM08HbwMqyCJXGOK2o2i0JbOT75IuA
BHk4AUDO74CFUQuvXMjVKxakPwhcuNn+Uz0lQ/Nu8HdyFJOJ8vHGU57moTYmX1/3BZ0TygTU8OUc
6WM342gzEnio9b+/D5Rc5CFn4LotG7ArTNDKjO/4IhW0Tc63O7EALnXuIh81F9GER8/7T8akLMDq
pbo1A/CWXwc69mwjoC7O0xM68tdbStuxHucU+ARYRXU5/SSsxPg2o4INjfUayRPIHgCrH6vJo3qf
FkiDUheiq6nE4QGrbBbAV71hqBOVJwFGlDumgZUQZVXErgnAKgYYnaet9hdf76hP2oH+cIGJhQJ2
nPQ9DVH7bypOrDPHgsCzPUy5HJbjN/sJL3ehxhWzP/mWTpgQCcuA/RfR05n5SEMgcj+tp5HDvGNn
ig3MrFg5jgPbPYhQKwOR/bnJBfEHGeSVvtELvnotxeSB/nNp0hmTJQUcdFcBkduV+uhmE/ZpKwwS
LhzPXJmSefJ1SBLG+RB3ViMlSNxg0sk2sHe4tscf9rlNLwV/xmcBHEg9fHm+R8MuajAk/qKFCeSc
vcUmwBZ4diYqxQcrHhtXo3t9vXUaYYUAgNjJkhyXNB8zOMvbdbzav4G7CtusjgzrsKqV1igKkyBY
WivAzxLTuBBqSAHUvgiTKZx1Zjztpv3gPJTAG0t4n+fIv6R+fIxCq4aEG4JSGDNymdzCadS95gRt
H+IutEy6HH0d9JwFfoCfJg7of9kyzWzgEMilxfH4wgzyTwb69aHrxc6Ce7a17gBIVGMNWhfvF167
gMKHZqyHS/1jXnjAi25oNrVSkr9JqZ25hGIgLxj3hZst8kBXzIbafGAIDnwTgq1b5HJ+nwZQMCNA
XlG4791eHy3mtMrVty2XxEpgbgVYfwuMwDf8nkDAJRs/DWW3ZuASNgfWHVgImSEJ+t+dt+ix8y4D
czpfI96yxkJ3Fv8WtF9VgIR7T9DcINvqq9a78uUG0x9tsbXkS1wK2vonV4iYjTPsG94doHo4ujej
4cJ7+I+VwVBLEl9NWhL1llqxLZMme/mEr/idbabu23TrqzOB8v0nFJuW5YzjngxLCNJ4l8JKC9QD
GT9cJNrKK8waUN/6erkbkb0A4Aitpjndarx4f3Y0Vm7E9X2Xt6ro25mHcJARDB573+xadlsW68+q
lW32KvdgsGfcSmBVbH53y530EIF+8TX4LAZ4tOsvB8u2nxOnOPZEx9XoUMHVmeLKVw/Fz83d372n
aLivPepOYejPxRk7JowAJo7jhOCcLYY8gkNEhusb7mxycEWeV339Rbbpi3jakpk083pjpaklxsyK
lApMDAd+zxI48c7pCKI2TajmR6qyIPPNL33hAefrXb9gDXq1l+IzfdZj6tuXE5v0DjJRRAnRFIsZ
jgb+fbZz47Wbrx/siwBv24AQN/8LSZ5iZkTc+I9EJxymDJ0eE2DTv1CQszSw/MVEpxYvcHe8CDxW
Yz7F1fCvkNdcY1RcDegMUNcGS+KmEgOqzcFMP3VQNqSbccZAkqrUf48ir6uJNI9TByTOyaRr9d2h
50Lkb0pjPVErcmV9TdRY7yjlcpnu+ijbD4f2luwsqjAAg/gdQ4KSH4OTwWWasA+APdd/sZuhYjav
Sn71xV+B7SnKYkTyAtkfwfcgsTvvG7He5JgS2nsKuIMpE6x/w4YJ0ROMbD339tj5Uy648Mf8oWzY
0p/ftme6JfzVethDWP/0u+muwpRjBSxtsimZFe3HNK6UDfvUjRPdMkxF5IcW5Q4fqiQ5oH2xkIdR
Paa29KK/nhcGo1MrA2FFYDVDoIUjntAN5t4GaWzXS4J+r78slHo36edYE3vkceuD+uN92Q+CkGou
1KViECEixN2vKC92eHGL0GAuMhJ3ALt6D1rtXI9pmgfYnjPNp3DYKxHnPhxteDS2VeErrIeSYABv
1RWWuIetKPn1nC2+98NmHasuiGTltb0sCIv6QIsFqMyGN1aiD/dT+18Bq8QSbtEGwMSpp0d41l1K
EbFczTf0XHnb+x/S2oV4NKv1BdK+bsIY+Qdha3LZ/Wwj9/SJK/Xbupe72fibGmnnPrQUcjMPF/OL
aKwbiJekR+PxeOmxaquG3lAff+zVj4qsnO395Cg6dJy+E4NYeepQtYk2h3eup00j8Glofu4Jrb/x
L+atq/nARa2mdBdgWidlD/VDvxwgAqBfI6U8bKsd/IxwmQQsbS6RLaBWatt5w3qwdD0KWtBlaqW4
Xv3gYvh1pYXkP72gnJr7g2kVL9s5R/lBEWvKS+p4bbojMLTbOQo+NoypWKqAfsOoE+efx6egGNya
MLFHAEjTPH0m0n91HMudaKfeMd8LyDdvYX6jQxdf70aZumbjG+DRhvu0f1T9VWeMulH4Y5uAvFuF
k0cOUWQ1RTsauEk/7s8rrHtQcAXHAsjndgF0udrv5ob9i9Gv3L38PbH35LE4CBT8X/B7eTrTmHii
tkFwSWbPjU5bgytxdoDPG/r6ipn9P0VpF8Mmql12vscYtC9ARWkYCIQ/3dK9HDC1DGEcf4faL+nE
dQLmjKX+Wg7/kelsZOWmJtTS5EcW62MFMq3tFkena7SQZKlKxzzhNgWwyZGSCYIxIeOEyhVNbWAP
4lW7Slrn+/xNGJB2aWqVRrKV3kU2WzhhDX7Bk89aDhNDWN/gnM98GfQC40E1aXJV6CZgofQHzsA3
qTrvpaxYYy0tpoUxy9jx/miARV7341VQ20Ti8mTxJ2TkS3SSpU3ZO1Rv7zA007BqmI6HolxvF7Xl
zr87kL/iIwK8aPZNSp+EMMY0P8CGGGX8IPHqCR7bazmIy8GIQ7uBXVarXDVskmFq7uyJ/QlrGbBY
7i0odT+uCMdRfhgLczr9zNFuOQLYdJ1C5v/RNj/I3tUa5WFuRRERgyzTxBgjbLHCbTo5fq7kkAlY
D4kzKcFPJc8DF8V8gxP6ANEagcf8zakPCZN79rS+1OGTKkI5wB7rxGclMLO6qIBdFXU9Vhng+B6x
on9EJTgoQUoTqJYsVHE9FxH4qv73SP/Rw94CR677bYy6XdDcNojUk2QqWJzw+AQdjP7pYgTNXir6
6uw7QQufg2yv+1n9glrzYccA48bopCvCicoHgsLcaFFnlQFj7GDhdMyt9NEcbOnzgQyALtd7TUJM
YPbsn6T4c3RVfZ+YJU22HS2f16IDklrOEl8rMHQmQt34ZZFxP7gw51krqc4P1U9dTF1Uxap7wdql
0u2B5RVy4AeRW+qFu30a+iEHXklYTJBqnaK+eRIwFxVbQjGpXFZNEcXzEcFHdSvscLAHh04fs9eQ
EagV7WmZ8LnFlgfWPIsgaqYeWwmWQqKfRkUTsqIC+nxIcRFwebTNTEC6JqR3nNbxqF3v3vo7KZQo
N3lwhZa1tyd+ofmVdptJKPsD2n2zEgb5bk8RepGNRfOikjcpA/2bex7pwsa0U8Egg1e9r3sbKHxY
9Hjg0ktF6fGWpYp86AXMcF/RhkBYkQys0CuT248LjLlzapytqKmhatTbRONacKVuTJ08fPbsugZp
beiXbJ2rtTjdybZMT9faQPyPsWuYkiNrrx8eutA6DOuh5aoU2gNNDiWQd92t5YU0XwwjBstZZCwP
A9UhUJVYMGSVSARrXufNEHWX6eRUuwRrubKMpxiaphT6qwQZ7MWc6LywzAGIE+hfN//AOrutM6/1
PV/2nQ78PbQznoSoCtYANEBzDO87nudlQrp4qhiwk7PzKpc7By4GoAAn4LPwIXSSg+PeZMCmK3EH
mhO4EVaRjiSb0n4BTQPySeeud8eVOsfx/JGYPXwCKff95kFLc5+3hfaR7NL6mqy01HbTmcS8qefe
CNQHb2Su6i3XnKy3HtCwujHIcjugKETj9gEB8I/rDDKmCf2teyxu60UNLWZS9h3fy5u/ZTiFFvAh
R7ocN5smRrqy2bGg9ygXGPf57PSJU+pcPyZzM9Stubjw4bsesn2POwFbKaIVAMIls4ab7EEvHPku
RJ039BreG5dsS8lJ08Z6L76K2ikvBdkTFXskmN5EFUaMmAPQWyYO80hFYu3ECDXoZ3QiRaJWlsxu
XhnGoK2EvZu0gZXz32tgRv3Nht0njzi4hHD51s2HeWDwyvSP1HTyCNPl9nOo5tJTscOgeNfIPm1R
YVH1Ii2+AOh1sUr9OUt2WS/sKJ+rjF3liXUQVusuGrgvjZy+yIAV3dLFOq67bTBF1DpHA1IsTRcJ
F5wRsSLZjqkPtBRZtDGwPe/NxsjO3HuWbnRqOJeMe/OwxJp3TDVKzNcO/CcBte5V6D2jmPbQ8MR5
TWmUuALUOklbTmOs7GKbRfgzDRSO6OlTpLUrliH+2h+qzfer33Z8vtrwNiXjrZeG5nAhPAYhToty
Lq18EkujoJf5yocpfqUlKwGglcCT7/pbwDkNzBn/0qXEETpPUiZIkCsAUvoDj8RBgtUR27V4aH9j
CAHtwevsyqmUrorLx2ymGl17jXk79L2XyGddrIO+cRiNFkNnmo7iZV+blq9dsRXHf/oE13CXkHKa
oyAKkU62wEcyGutxL4TODOrpvOrUnn5yFg2QJO66WRjDl1vX5kLJeixKWhHnPLahPyTQkNkHyhHt
gcj1YsDWVlTYUULi4MkKlzKY3d7TmZ+wJXu52C+D8f1Yf9W6mCAFZfGsII2yowCw90ysvZYIeknr
deHFDPzZDyOy6BO26nragP/XwY0QN41xbj1za7amLQ17PLcWcDQCYrRxnrzxbSyR5QipfVVEwqpU
YbW4uuCEjEfnh8BUcBr9ftwsVTmVDx4BMzzWU11zrk3Ik70HbOU2+NojbrIeXYT+YBhQqr+qUp+i
kxNT1jWc6tbHj3scl8cgT/6Fnk01Cmra29130g7XPfY5p+1fHnXjfvUoAZNB4wul1Uiyc9+9ru+n
Nx0URLeOvM6jHlKWSL9sVrhQg3mHgjBi+9ckykVVqaJLyB3ugKujC/KQtYIMRsbAh64+oW/NkVv5
07LbV7odFn8+jB0lc7JAx00mX7Z3Brkr8fg7sjrGB970jhpEMpJzIenzCLfWOpxHnZXdNDE17D8a
zZj8ok6O9Hg3++dd2MOX3+4vqpLnVfp+bjE/9M1S5WMNarevIhNP5LjZxtD3/FKuF9wrg22ywL3w
tjByGD6VfJhUwF7JYInOl2fN3F4drdXQT+TVZ+zS9zC5hVnWjW8qnqpHYDN0b6lP1KVpLgo45q49
rWKTjzXsAuDBtFe1EZj53KCM9bnT/IRJh8QQj509Bn66lNuaieRHVZil1JE7IKSFfTQ+ATX6mFEd
uzNisWhsfkh9k9dP4uQGoBTU53MLHR7UVzdRvC0tkSdG5sQAltGUNrlLRZdqx717SoJUHdjpzhUA
lN0qWKtRfsE5kvBWyNVeu/VfroxR8THAd1TjW9PXcnZ2z0cBmJMWJSfB+qbxpMb6fDxzWu3WBVJj
0dv3O+jjPoG6fWA/ilxdvS0CKOXLQsyIp0g8JwBX5vCGi1uy1pVby1bpIu9uJ6g+qNkAIoHCQ3wQ
/IgZQPnTgLOHOaJhRzKH/YthAj6kKKX/MLoyIwlzBHjWwn8k3i+/yejxgeFjYI6f8H6Bs2lIR8vN
j6yPFIXZvaARraNjkA5vsLHiPf5roVe+8pfZOXdQncd5DLoUIGqhoD8rMCfXShSro0FHPpAqwSIM
z1HP0Kc8TPj03tmDPp5h1uFcV63kTYoWB63npRFcuHZKWr5A8rCK4d4UZZKY5Ae4xprvHkdMxQKS
ne6nuxEEgmohnPtGZX/9WnLRQ4BB55t0kEZAKT2jsHXByWvzctAr6Nu8l4CR78szh2vLynVdJyBK
ieENs4TcZQlL1rqZTS2OF1hWyzGiYad8alIh35NlhvmbbRZOUfcknuq4S/JyuQR8+bqOqGnUPr/8
QTxZERYlijSuRNEPp8OkVZz9KhDSNVpXXxpYRGqqIRFOiUqjjH/wadK54t5aOGrMdArrWHsgoepQ
rMtzYjtLmWdF1P/s4P+HOpgwZR90rRYCpnEO9JN5IPoD6StCRAzDkweQs26Boz1ESkxCCsO9m9T3
mnh6fxoAAXSGfWyowolRSwjFv8VEx5NO+31HeLX87gYUEbuGmjMBQSu8IaL4u3Ws3rgozjQtGUgp
iiAqjeDt2UFsdBaobKaCPnrn5T3micimKZ0/gfBXYLzfMVNB2E6XaM0pgD1PLUTG6koYtkhaQHCX
xQFa3rX8iF0QsMSMxZ9EAUPzJ0LEvus8c23R8P8p+I7DTDQQhLFOSCSYjrt0EvPrSZkx4m0Cv4TC
xutftkWE2MNG96N4JUih6icaCmkeNG+gIlboGkt3uZXNYlWDGuXUWFC9Ee1hmxie37Us8Zm5io8t
iiysfdAZ8JXlxXk0bA7E5hLzFW9FBQlDrMXab6WSho4C+8CKvNXaGOiZczyZmUIuemRnNm1WEWRm
0aQ7FM5KTtzpmPQd/POslBpOtLfYfrwyQeszrfE2IBE2uggiobLoa2WOY9Pb/98SiS+MSB/a95se
UoB8egqu01rOrR+10wo3/YCWfVSX8fHhw/tLzrZUkX/6RSCv/1Cao5uPKB2cbloazSorC7/CJnXR
AUkBfUUaXYXQOXau8IFY0i2ZbfWIy0LcBrNG/+k9JvQzNAGr3/W1V7FT4r8aDvhU+hunPnfboqjq
/sYIE2jLgef5c1zZHpTKXavEsk/qu/WxY+/pzBzrkDEX0NNksgR3bphvZU7gaNWzx9w3JOhP0EZH
Cla5nNP9C3OwyHiCVb0PhUOnPHnl5yBXISb9qsxQ3q6ZCaiZ+9TSeiHlUH3Psk6eoeeuIgBC3D5v
Ei4ff0I6fun/52vElHdYbccwr7DiD2wJ3QhRezp61qckvzcvXBIh5XpA3ptFYlmlAQ6YYwPicAPh
nHoaMNRNad15/0ENe57IxuFEcwEBqqdY3btBN5FwmyU8Ro3Gm+Co2K6KgNZuYxUhe3qdrmREPaPE
DxKuY3uqhBfZosb4VxTnXYY+JJcm73s6v9wxQm5gyoCr+mhPBB+XBV6o7n0GOzFgFbcFMVBIcuZw
CRzRPlPM2R2y5Stgouv9ghaKMr7HxteuNpytmRfUwfYZFOupDyrpwACzgAGt3BGkYWXS2Pm1UIcg
UjYpFsmzwMTjudAWANpPANPKW8xEJl/kTBbwq6ScTrSbC+7/ifbuaTy5InhqdK/kFkA51Izvlb1m
g8nRKJI4UUhl2DrcQpq5HixAnRQvR+YjPXROC3hNPtkfRljBXb9mdCnTLHgh05RlV7+CwWkx2Ehq
ZNOw9brF4EzbCwlpVns6mki9ZBFP2XnML+vJMCnuP5xgFXfk1FkLwnN8zmsCkHnuXyyu7x3d8DAJ
vjXoFItkegCRAjvouZVtAxB9DAuRNa6rees6jhLJs74N44Tcy37+t3f0jWxPj4Zyt7LshE/8YChw
GIFrV6HCtqOpQxvmTX1diPlwqmd9UTCy95RDYJMj6SjP32dLL/FMHXZpi3xalsMX5jkRVvbUgalE
kHdsIRc/vWuV1QCsrDPwYhLDJF5zVQG74n1mCY9XQz39CaASPv8uqUkPnDggP8CW8yjL8nSX4IL7
p8Ls7GB8bgGiQKJZk1FyDrrkEdJm8/oYBZqJoWmXI6N2cdWe5K4EGh27a7ySs8DHlepbVG15n9sD
6soEcLeH7bmbi4n9lrDSo5dFkvV0eosfR6lIrqI4pI+0ZXYphpNXd7ov+Os4xhzS/jTuPvM5Ueo9
sBoorQs/ftEZGNmRUOpAE6zocG3Vs6E/2dJR1j0ChKUA42DyAQgUFG+Z2/ZA5vo8xNXY9vnWYvVZ
wp8Iv39Ajf5Q5mu0mLCWmJtKQZojIKyuLaN4iDHJNHUTv7Do0Sluj7+mTZCcCwwo2mi9wu9XDH36
qgEB9IeLZcb0MWq5CzmRoY6rgrOfZBFvRJKqZ2H/o+t3/Pi1cq3kYBopuvo/czd5YrH5M3BLzI39
lSqLrkzSBmW46idJ49fBljt0Hyvvm/aWKDNP4vXljuPbZEKIPdrdWxBinPpfkyBYiArpsMs/R5aC
zWG0MrwSmFbdf1fhI8DOTcPQkzxcnrkgVQx9maBxrOCmjfDj+QZmXCTFZTxfeGOWbJO9+J1HzBUW
ISPYPPWEc56uLVNyLaemtwytq/kc+XDT2C/RG6Ops3Ze4RAknlVkjS5L+WAR7Khfz5dtJ5jwHaLw
qAw6VmcbsMw+vEm643T7WeG+qV0qpmrW9/v1ZZpL6K5hhZ3TEKSL9TBHjux1O4u96ietxCDuw/bB
mHopD1FAjDNPYAmelNWvFNJ/dfKJ655FoMl9u69CQSpHWrTWdBuRn5fFiW0iQYBPFxEZJaEctKcg
D24+bch8olps2pQneyRqgsHjTnUIrYZzUIhTMnp3d/BRIervEsBl6U+JrINkErIscK7THzAn4Jrm
jEez1GVrxZQTpLXU22Br/2RreAB+Mc4EsLglZy1ciOoOiX8Fsnr3fUj8cD6wgCaQq0yc0+MikW7v
UKQIkhi+Syt093vp7AsdG/YelUMxwQ5hdvZW25v83vYUaP/ZaSM8LidF8N8CpiVs3iIGcv6jU8zc
Q0lgoQ1IGSkkvBr1fXHRBiMODiQiFA59Pr3zpkZ6JM7IGtb3fCTK1QcRrhvFhrsgnnL5Jl/WLow0
zUEsf3YvgAxkSyyKT2T1jQgp2Gmh6YLXLXaeJCCaCe4Btecl2WFZoqTPrEgMu4/UP92l0W9bAHuT
SB+JTAk9c7UZboHldr5D4lprQCrS0mMzc20ygqgKF2O2TvssvOexphUXdIYyB6KzQ8xFp40I1r0+
brSaIPyGurvK8fcLCmvMwbGgrCntdULkyivn0E6Hkq5WmFEoDqkbo2/AEdw2f0s9FHh+rKRuA3C0
3OT7KiRVe8p2mGfZXUOdR1E0x2B7HjD/ypPDeb6JWc0jZLf3UCK/iTe+Rphi/frDWeHg89CMSuKM
OIYJb60y3isVUPsafMQcb0wdmQIuFeCd8uM5Tg+2Qhoru1d8vlz/VfAiYgLHcymKmxJRz6XeLPxx
3i3PI7l1m9yG4zTpf8Rgr5OcpQIVZEmOxs0fb4vEVZ5j7g5gGRuEDYPIMPT1xcrFd9YLCojMHw4s
3kp+9z1J0v1QM7gc6IKBQg4u9pkJYTYfOy2mhqyJpcXCDFgKWEChjexlxlPASePk9BJxgt2K1x4y
vTvOCFfjPbxEdLuP2KKpt4ww5cpxaf/2VD31+zHkqg8ijbqZLCutBJrek1GTngnt6qopuVFzMOlz
766QrLyDsLPzsfr1/myz10he9DyCycsg0g6WV7+lcVk4WdUGSmHNDrNT7Ec/eLFbABnVktVwKq2z
QQJIRB4ZiOaXavfWO28kpQli/WNlU+Mg1Dbul2XJ6iwTnQk8XmWym1LYxTqoK2GUPiwchx8knIs1
j6h9E18rwhq16S/vfjZ+E+0Q9YUbTI3UzRCHIY3R7ct5JTVfvTe56IZHYhy8GDpTG2YXndoVD+J5
rBOQuKyRXvkoNNb0socw9JzavbqybLJdMLiZnv2GJHmyDhWKV2vOjtDjKxopSby7rEpuQw0hUMXR
uXOjyI13BykcwTDl3HvAcObfncgUqPcZ74TEYgxqmgMv3NoiLKgfiB8o7Oh+x6KDGB8y59KgkLQ+
xsKBIqk6jPCot2EAV3E+tMd9Fkm6ENx7w34dSuPXClUzzSj2llCaI3L7UQzVfExmbVUF5+4rV7VM
ogMJIbFQiSAAchhvXLodIbgPw4GuapyFV1ObkM3iEK5gTVQ/BG2VVqjA7i2APeyFsSp6fTrnw6WD
uGeDU93cNplPtB7v4SidZ/TZUU+1u4OTmX/L+6Sdkdp80UtZUQd2aSyEA9p2NaK2V0pAB5AnwyJ/
NulMP3LdPWP1mir1VHxsUb1F1ZxTo3/dFARVV+ywNlZCA5EgVApaVZbkmqZMXthlIJNRFxLTTAwL
6JDZ9RkqZq5eszx+ZKKClCHe9+4cz86vAmEYk1EWAQst5mVEuwnYiOIHKDVk/NilCO5bRGVuUDdR
GKRQuQPC5r7W8zAJhdZabsPPSRVgihAg9fbMaFvcLoZFZlB/dkoTAEiXb+gJEFarGRJfGtN04QcT
0dBfsMM2PmySgLh9Q/Bij2EHbE3u5hLol3gQ/xe5AeQeRBAMHyVgHvjkg25t6KJYBGMhex/2WoM1
hOwO+sXWhmc0TBs+6gJaHBh3++pNlTTNWvjUHmwhDAaam/LbvF5oTvGiVXQSX5UZQ1LKE0k+MLUc
eyoGLnApZlXCKHrMQ1o+UglJekHHRsdp5gWyaEspe8k2jR4pNji8aIZxsraV8JfhHhBtcaRcs/uq
dCM0Q0O9R2JJXvo7CHxmruP3dEf8tGs3s2CkxQW4E2SBhZw/indhkzEYvZECnVqkUFGAMJ4Rs2W/
VcpuakpVy/kcpB7mw2fLgMDewcbKxG0IHORLw+GmhqTvXjdIva7kfQSFH6mkO0vmhigPhkDEGiZ+
wxP2cXJQrkuNZQQohDXFtFa++nbzuHcaTGCoTfJLpatqX2120vaDNXndFfJOuztxc+0aL8XiQ6Cg
7BTyXPG3fz7aOgHBhz5e5E3KNXzzDOl5LwjOmUkUSZzGsTzE8VR0sqGfs9rIjT/1AvEKz6+a9Sde
rXf6KU9t/QWw3Q85vXQF76ES2cTCfvIqPD1Ji5I/QTXP2UoMEde7VaYSh8Flmled3LPwd0qEbAzd
C+ZzNlPrgL/MQuJ7r/mZDTsoXYPWowCpY6U5zTHUjMh4Hpc6tYwTKOyeB1OZOoB1mMrr8zqIsBKD
nkZXxTwuKjLApKkRbf/k+194j1Lp+naUk3Oe4TktQZaawPKL/1b5YS0vSXNYL52qmj51w9cPHd14
0yeHCPhamAxasiXb9ws4uTdzjNZuUCAuntKB7e5b2H6SBZnBy4ismseHcUFw0wU2Et3tsRy8H26h
eNtOu18YhVBfIJhyuu9KFX9jlLn40fRkqbqXJIiWolUAv9fCK4i4Hj1K+yDBqc1pYMB8CkhJXPKR
RbCXUCCnKFgdx67K8yKGHLr/tzBX1Pq2uIPJ5EMirUazRcQ4zQUx7sFjHtfcBQ+Ec+vhb4ActwDN
1sGcbI8uj+ucJ3e4VUSbO+4+KOi8lTqNHXPLgkKxt68fH7YJFNi48Qe6eHVHfThek1CMNquaE6lB
peuiwD9jtTCe9nk5R5EMQ6iIn4OYQ/ayEBSZek/CYUeihNn98D5SVNIZkOKG/mMF6C8sUdyGNZoD
FhAX1xeXCr2MT6OxmczRKEr4WYy/TVMtj+0gZw9itEgv8Opfq2IrvK691EWYAB9wUrkBEv+5BMi/
uzIV+1TyU72dAQwGozCeDZ9o5fCukpfPYqyG7pag9A+ERwGVA5+nIAQN7xQPNUlYbWVyR1lXmFeq
W2ow7bioSaFE8qdYgkHRNX/txWojsYsiXSGj7Z50GFpNdYdBqua/9DyYSXGRi/AVGfuQXII68nrK
xubr35aSxHz0sXSvUQFDiyZPlNp/h/jeNDDu5B9mjLBw/mXhqNUGwtEc7o8HvPZgaAj+9/3/uoCc
TjesgS3FHatq3zMw0PXkY/5v6F9/RORPfi0wx0iDsjebclDXikhFSlPlx+AlrdZpD8WbcvZ/m8Gv
jRtKgj1x97Kl+p1u+dz7CnRj6LMjFANbb0MqmG7AX/NOP4Rx/5Z+iZzEhn/SAfBk18gahanw0adO
qgoReNS6TlX0vy4MbKTfAv+cGueE0GlRmNg06eSgUmpdkav23qF7p4zlmdcLI906hcuSchAr9vus
XKrvr2Ckj9QblZt+qk9Djp3b9Cd22brGboUub/MZOXtbx2ubugcvhTRP76o2YRfrukYCBEag2QSV
Q9OmmW081JAsmYn28Ul7uVajKLUDzKnCXaYTmvFYejDmtHHEluKikWxWjkEkmGJFzC35DTUwishY
jNI8X5ZzAlYiAUhOpDwRPqbzArNmhGsFmAhWNxgJAsBcSp4l86uB13T7FJxKTBOpU23RmDfAvJqN
xQk3t/C6MpfkHosnpfGl8d8/8F49lL25SnNkVq1Wci26LNGDmfXujs/nV48WP0ZM56yOrYy6zMIg
B7eQm/8eqVl1OAF8DE/iu45HeJa3+zLuMGX975E6PYHt8M29gHiE8j0yLKaPqoq5A+N0qyZkW2xv
20KDC9L09oxbSWeYZWDiTcUyT/eui1zNGAhXVHjMR6jnpP2+GhDfGiLi/bGvpL4V5G9234HQH5AY
XXvuTiZTcl77cwvuaNhR48dKk37D7M7FRcOoDidiVmRODt+Hwb4DuQ9xS2ljXTM92mC7Q5wAFX6Z
IJHKzitlcn0TmBn/bL9c3S12j/4NJAFD2PxMC9Ml6Hvufte/pnuu8GsSuYWUp/9WHWVLTwbYDx0n
iNyjsnm1+Vrfv8OP+rkLUaKcL8UBb1cI6K8FVjf7phHk3ClBxO7oNuHsue6E1h51ms6ZI9Zobq1C
rmd/iaV2L3v3kiEZzp1hZjZgrzEHmrZKbjAh39Kj868ofHdGiPAjogohSC1idWwEzNDD5rxppKVN
jibHCvy3OgRV1N/aR2gIK1dOcegxlU3JkH+S/GfE79wwstoD+g5usAdoJmd60wO4qphi6hN/0c3K
rNA8WUvb2jWRpcscK6rmKScRkldRIhEapO/3X//kPFQxLHh31UsZjcdv/XPIzTzvmvqqph5gUkPn
FzSvgSshRL00l2XPjr/kPrzzUAQmF7D73RbRF22I/aCXEYFk+qFtEl9CvldS/m0OD7gHi/rHbNiF
kKb3LVaJf7M3FKqIFTWjqUaWW0rClhTmqrBgIwNgOQRYFA5RzwWTGqB9LKOAyoFaEGae1+lGddP8
C/HyvnwWlzrPjjVKOczbBWmHaZRujDJ7BqQ8nth/fzYhYKWC2LXpMYAPuLuTNJHxx8WwIqsHEPND
NHJVPU5/62oQsTS7tKQt/n6u1+ZjcqSlR3wWm/LZtj2NoaXHrGsp7yF8+UuyUqembsQ/n1VEYQ/p
RZ/lW5REzkwqQaxl8JHdaspT54VMLJGIEzr8Igjcpx3iGsYrE9aDrhP7SyT+tFL0kTYsjG35KcKr
IU3i7lZ5qp1ko+dBDiuQqTIZg3pHl3O4Rcuzp+ESmXM75typncbDc0YD+q4IuvMjVht3nw4ATO9w
rGzuz4cRvr4/Ev8IF9bnG5q4bthXLoqGWLjXmJHYpCEP+acvCyUf+Byt1e8s4Btp8aeRKMFksudk
PQFHCqR6M7UdUo2p/Yc+q3O2pJQvmCC3cOgtYBQQaITxAg9HYwGQ8HX1Txp0tVl821XxC3djnHbo
i3gnN+1YqI3Mkccy6HTAL0xlcPNECqRi2V3xN5+78ejGbdDsEs7rRLmpiGZHLkcOOPt0uDBLGlH6
EXvcIkeig1kct0Z0NSb2Oyq2qIgK89LoquskQ6CjgzN7GgkMZNWIQzsx3rE9EYcb2/czYZysiTDd
A/U0v3PaYzjxMHwguGk05sQn6MM/DQ0501PTJB46Oh6QDwe/3wmZ2QGr7hmFn1QbMGCjvedB4VOE
6zpm4A62hsDJt+5IYKfrTKPr00ZUkbrgOKuIp2ixjYe7y0WVgWV7n+6DInqCdztwMHYOiljusvcH
L/kLArj+i2mfemYW3+1AlwYg5zfqneoE1UTsiE/QsPDNnsdFqX5WsbeYst1IP+aaT7A+iuES7LPx
6DKWbY/jVbp3WKxSQHDoH6PNb2EW9Fnlk8aCy679viKLipWa9QZd3SvzGswxakFvApkKvwWni0Og
plpgv2EDuhw24IwEK5W3dQMkr6gJDGUSpcduu3MW3t0SPAaeGzJZi/zrvysxAdr6+0oFtWHEeFLL
ahKuqYEnaEqGkssi/9Pn4+bilZ1F6QD4NFGeBHLHqYoxNb2990MsM41/v/9ly5DbHNS2LHe0is6+
FNRqsCm/xnHnOePQV7G6cdo5js9I7RZcBcin4zkY0biV2Kg8n/zFU3PORAeMetuujN1cCiaBDYJq
UWAiLxt+3r6E72KiFzXds0qje95FgLr3ZJeGPLLF6lmWP6XWCa1cBtYn0kXNoZ/Gc/oF+ticO0F7
07XDBDbEai5ZFoI7rzpq+VAGIOjgdQ+BENln9jEgrRUivYrFCgxWF1NnVcWLYFfnoW68fLWTIWky
CZoeQ7ncerH1LIVoZo3w0RqkIWldtseLqJpDKSaGfAZVqPjWau4+VsZn1nSkVRw1cj41GDo9rlfb
Shi+cAuRH0kgWPCtmIKgO1i8rvKbr5JyA9CoNQkAqKoAiPlnh5Nw0hei4hdWIIFtKCZnE2aqlPT+
WsW5Bf/7EdGQRt7KCYqg+s26ocvkLIXPiNMBrJR0TP2TLylFtXAyyEoUiMK2qshwrwC4GLqryu+c
aEg6KCbae8ctGWSDxAZmZPIWQP9kU2efkAKI+ryfGBG8htMoeQPUDQKUcmUIxht9JEnbqydkUija
Utw//JOg8GEfvzKT5lTbMkOUYNIOx2Qgcd42EjDJPyjqey0qE0QSbXocg4dIlvEqz1UTl4KeRbIP
rNWWZbwoiVfaI4CmJM5r4n24upHkrLdGuvXlOqM1fvu+aOtaa6sNONvARhOyZ/Wt3ePi9zVXcW83
DzprueWqLiO7eI0dhkQLOZLMWHiJz28ByTpn32G0/T6Ye5TyzqclO8AaM74nWxAeIhtDskCdID1i
gxahg+8yKXhbYkg0KeZyHINyLNtchC9OKiGAR41OnvwpPrKk0UAlQ4onZeESXiFnkH3bhzYCGysz
SVadoM26coOS+COfPA//o5Als94aXvtdYu1XMjIo3UYTPklEVv7BjTZ/ZaZXWz+BF4XKdMhvzvcJ
xCsFEjbTqLU8t82Rt00hTmNU+fJyFngm9iGzsYoUlCeGytefpwO2adeuhwSSMsdVSPQzzhZr//w7
MMCHQImDLMqC++EZJ/IsVgzz/8GJwdhvQ0GigavUkzzHrZYIj7GbwXaTOOUvJ3K6kHQGLnFvQ9AD
eTlI09cHFIedESHhtY3siZAXcB7+tDXth8FFI6xzFBlaQtkV/GvPHC0F/nogNb+aJ5IZHJ2zzOkV
uWsnKLMJu9j6w4u0lqpbbM2fbXEx/s7Jz+MJYupr3AjYyop1CXnrilPcr78MgOU2GqPkMN3nxIZ5
Uf8S8wao2KAMPdS9UIeRzr8/viV85wTREhf45yTp0PBdThf3ZkKYqu2svtFuTGIAn6sIh7gXFnEz
G+9jJa6EMfqbRvKITxfoz4o7+JdHZBq4D0QQsP4+HfLqPm8OpLT3jIMeoA1GOHrc8l8Oi9Maibah
UqpAgfBdrquETrsUdi8Nx+/f9fwfebHls1lDT28B2nAZNVkLP3LLwhCR4W+wgWOZ/yDWq2+NVgBC
dr1eZd3Co2d6i5PDjWqzdlEl2M7ID4JQinGBbTbc6pqs+J3VQ43WhK1CB/VcPvsJQGaR2xk/cEnn
6kMOWlSM7gNS4ahc75MN3Vx0KvfdYqKgB5llMW0KGeKOBDv9e4WvhIyJJSzKW9rdGg1TfFTHK9VG
tloURWy8Y4EMLkxbnq8U3nU5LSn70bYmGi2HZs4ezTXTvWBPABNU8FA8GB4hCrizpL1rYRaePAWe
mjCM4+gi/6G5XByoYqMsLIEzDnsY95Mc5sawUmcbusWJfX0xfdhAObKkGFTmpT+ISHUY8KAVc8iw
EQK/z7Ny9vSunwQr4U4mQhGm/I3rtFTdMjumzb9r47QMCn8IdHfhyAftgEeefgIzNDTDAW77crar
rmjRO3Nrk0m0/KEB6lUCRd+i0gpkDQ23Lb6TqFjozDi7dLtkwzinUli/wtghCAZjMXNlF0FXq0rN
tDRPHzuMBZdGJAP95FTBLhmCuQBLiw6ZIWSHcKLKM5TqCXYf60pHKN1mGRfZ42DszGaEpGbZjM0h
ozjBq7TpVOuTliLNaDs9Dq5+TrwXBULEtidKZyARQmceH//qKK0ZLbGyaGKvDzHwKFoNBsLtdEax
dSg+RwfwTwyw2qZEJ1vFk22+2VLutNGUam6P4V/xvc8Toz+YIkxdhg0OKpKDQ7Y5LNMUFwGF8ZBV
Pq9bUUvSbLT6aWIgPAQ9pKt7E9Z7p51zFBnkHHPtpfAEaSPvuMTk9mB50JqIDfNOed6LA9uyVuT0
dvHr+sp79WgZUq7Tz+ztxb70UFQQkB/btDsNLxUe4ctg3MkGU/RvkwNYsOk4AoZU41N5ZnhusORt
9G0oVXZvZ3won0GvA5kDWrJH0rxBLZLf4aMDv/kpb2QksaYXU5OPVo8HASAe6WVOQDXC4PnOVdLA
odSXxYu3MPfpeSS/j5y9aAEkC8Ag9bnBccIgMcmV4h9s6CNcJ9zDh+3NfjD/tyHydyAgI7+iYYb+
WR0cLH8GF6S574zatIBVuRg5EKbyOFvQwFBNm1yws8Amf1YCUyTcjxXTxHnWZ0Uv4ibeJ2SZxtb6
Foa2W1vm3GeIxQd6FZMkqY8ga+ePmhveNsm/4fFbev2eqdmbgA54hbm/pphIv6uxb0kjg+8QWBBQ
xllbz02HCPZSuFo7zqFeRRAi/Icj1Z20fXV63uMPBWlMupG4W3ydJE3CLuI3a2orW7rkpZSXAOGa
vKzBiBae1JOg1YUxC3Wwz3sOXsdlBUsgj0/Bj3gEiN/NwRdCXXq7fwBAtMVxcgb3GpkE8VLGWcq7
v262jFAv+DMHonupUuxWLoVG0BLEULAtDhWn0tZDqDMa1dzZmU63SzXsk8r5V5qOLxOFy1Y3ASeu
OKIqU8mk7tOz3dmyk0xBbJC4Xu6hUUmVJqH/ZDl9WbzkQFFJzKg9M4BhNJ8+0SP9YtUeLFV1nRwb
Ej4ttPt1TwLK2B1slfwvK4Qio+cDziMmHzmN8WmXuHL9h2eGlki5Rg4NLBrWgfiBx0Mb52gvae6f
8iPMDAkRswFfOTVAvmazP6ilfIQ5qE4pJadRkT0Jw94W2lAJ2jtsVIXAj6opZ7nYKWzuoPyokS5Q
PjO2+Hge4F9YqRzG2ouQWsFZrGxOXSem12LbwG/O1xv2TGuvmwr/HvXN28LkLp0xeQkPwDKwE2as
zBmUlTYgNcfW9yg/tquf6uytOneC/Zpy9dXygUnNOVUq60DXelXOiTeI36IvP+GovRGO3tmMz3sB
POGUoufbJr9hs54sRK2dMHSZqTTyseF6rGOXUU3VtAA8oHCPtHKj/mwZweoqGNVoSxXD3Cn5+9dy
N00TIK9qO9AACPDdrVsHvfhjxnQ575t+Z49SzAEGFBzgk+/WLjqCQrl2+HKnSJhUHkbkluyvjpB3
J8/yAXJyK7e9AWo37uIFshiS7GIRsDHNRnJjGrwPNmvFR5ZR11T4IHUdml1DIOJ+1W9ts4YKjGcg
j/ELZAN6ML2eigUprkH+6qJwbobClWUPDKcscGOLAbXFBgzo4ZudlpZPorAKZFcsj0yFTIq8iHp4
ykkM7C8q+1PPHH1mLrueAbO/H2w5XYRFKbyLgWgx2MuQxHy/iI+nVIfS16kxJa18295ExnU4Lj2H
WzaxIrz5fx+giQsw2GIpE9VABvrPT02d6EVddfl6ltm0KrIe6fTKKjX+reIYOXtdvDJ9L81KxcgR
Nry3Bn9CxnX6RkAFhu42Rq+BRm7c4Zi/7vIPlIJcZtZzDgbiBSDAvvcJUMdgSYayFjncDxxAu2j/
QjNs6cSysfD7ak2kLIFXQjUY2L2s6H8px+OBR6nV8JPU939SPP0VKwQPnn8vVT/hLgobwuAus6nu
7nUozVS6OxYlVfrzT+ecq2R2oIZ4pEokdTTa5ECydcEc7uxbcRteDMTregIRx8ziaonxezQ3CfTw
NCvvKR+bJhY/wPJsTYHFnEQi9K9bChEBlWvdWIqmB9BH6H+QuRUu77M+yL1xvS5pwjVBKb0aXZz0
TP5RtbYmn25+GdnOo2bPYEDqLQ+AewlYItX2eGVX9PRmbzOW2jimAxA6Db8R44H7JuoPpEK4sk9D
VO490eCotAeDvottDPOyjIWzqA+Yu74tjLjyqx43yT60GuVhVAbn/JrQ8QTSNZyEo+VUIU+d8ICt
4e3SzE9FccDMIeYDLJInDffpMVFLjaqmcAeCs00j3kMP1dyeFgHsihixVKlRFvLSdfi7xc8nr2dj
FSpFgadmHVux8LXjvStcDOHCKCbU0ZXejCNW+9B2azR9DVBB3dHmno4PYsyfxRFYE/NhgmU0plkJ
P+bwbswJH+URNtEqYQGQvr7wUjNOesJfFmbMHiSbgsOaXn34v+9fLKv1IKWIEc4rBA32I64EQH/V
nAh31iYcTDkHihVoP/8iIwGQIAivFoyOE94sHRdretkU8iGSTu9XFPeI7IkUxfjdtLHxqxpXwEbR
OqpgQDWaNmEgcJN4nJILVSGYw02jqo6eEj1r2QQvVxHaAGBwXlFhmnTBBDpERYtmG44VA9XpHryv
XRtSOgj9CIMJRsPKchU4fy6zaSss21HBc2uo6eKgG3GnPSxdbj76zYMfrCul2h/nzzDyjpx6KY8r
WylJbg8YUdHKYVdU8Zmw1A+M/Gn53FHwIUnowPnjsT0oVD/6GeEwGAovVeVdo5Mg6Mh/YHOWVZh7
89SAFEsFwxP1lAr7vqOC2j+YJ7yPC0HznO09HPLsStHchxgZfER0QEQ31on1grBljJh0K/yaYMab
j/+WbuSONFVOhy7o+d7rsiqiy2QhPONHewgmZFrvueRZcJoPNziWsgfClB33POdb697y3ZD6uSAp
39hR2KMs0bi4c3tYXMTRQ7Quf4IWyUQulSHaOddjm5TCGRVeGFkZFvIi2HKCu4QX4ziegUoFQnTB
bpkBNnYYcwvw5Fv/LPZx3A+e/hsCX8QLmKHC1l7k3bBPpuQrDiRo2hpByTzGnhl+4j0KCYhwbpGl
HBxs5Q9lYclMWuKweDKg5OIagUgSGw+sNbUFSLd3PRZ1H4+tI+Alk58oGaubSgmpXaJTV2cj+VPy
cexwy9GyG5INhrbIAH8u/IR4OnAL7d5anrx6HOcVdoULv/UWDWdTfxE4P7xtWF1bPueH5h8EORYw
jjNj1alE7tktWX1YMdqEB+Rr/kVQXX6bbxawQ5pBDd/3NDa3Dpx6+Y+nyi1Ll0wasnZYRFQAOK4n
5ZPKR48ygchR1hedx4iFnI+nUtygsyYfJxDs857aYRiD6TGiefmRS+axLucgcG+Mfg5Yiu5XRKOJ
yTTmUqQrmUq7z9751DSmLZjcHjKrwOVyg+Spb4kjZKddn6J/xE31QOwm8S5L1RPMj64v/AaTtNik
5PWZ6pQOcDGXabpQr1oYXzMn55+AV/wG++GpwfSof7UPxtWqJdaoJDDs04Ypbp3MUZNJiftfgmsR
8DUA+VWt9OJQaKt2CDFXj8R1g0cW4pwHXTQEZuTWIEVRRyoUpkyW8CwfjBAjVwcXm+ZWdT8Jx+ZU
b8MWiM6Dvj1Tf4gJUcAdRJ3iodhR6GG5MwLncQLFleiy8I6awke7PUmNCmPloC3Gyr10OHAJi2Dl
e3oUr4jnj3GEr+VNUB2n5+SCGSuelVe5L0XUX/npelmvt6pxJFPZu0PqZ1f9L7q4kBmLvWshOEsh
Tt6/s9PZU/0fTwd8/tAvjrerQKo1DRtMC2Job6Nb8PzEPa16sHlbSFCyRlGKdFtNKdJgNGCDmIhT
XbE5YC+Ug/RxmDAnhoAEhFfeZ0SJeuypwFXTn4QkWcxtnfOpAGUOo9FBTqH8EuxE+XTFT4jy7032
2PkElSdJUlmAYUy/5DHhXgjz8mHh8lm/ZyAl0f7Edk3urx3PbKIjhlLOoaZkXkuyI9JsSNe9Ee+p
bh21PCUGirTLcHFJyitHbJsl1HyRvcPJB4fwCObZ2q8qqSvzvgT0Zq2d4ey+0S44ijJsvutllpnJ
FzzsMw5jcR9UPdhgx+lp7Txc8EA9DlyXbiIZ8QqOpgB/mNVJ1lDW37WIiJjUiymMxJPCDwDC89xZ
JgKZX8ccJp+EnY1wRrALXC7RkRZ5E1eHvh8lbwDcI4pd/rQdmsamtFlAbxNoWxERn581ENmBUxRt
JCDTc7CoGBVchDHPNtTSIlRwBgDMU1yL5TgAbEZjrwlZOWQtljVDeOxStlGFcFlxfgrijgFxDk/r
H+xY/seF7PmdeaMmBQGkfETeyWcqLRVd+m/sN39GAg1GiTmAeUCg8vBj8bG/MNJzWxfgD39n/8fd
yiDKkuK456xfCgSbNiylVgCv1Zstx7JCjnp13P7RdVubghlUtId6qMPo5bIEpA1v4V0fUcdrelid
aA5hpWnIQofdNkoAcTqPQy/lt3sbBDm2nEhUTy82SU3nkagkUPT9/LE2pBvoG/WMC6ZPU5kKtV3v
RHXwqb3LKPODYymcHNM5LXgBqrUvRVq7QY9e6E9Azi2cz1iQmLs/CQEvFkHo4XhtROEhRvHKLYG0
Cou2eGGdbSrfLxRGDFmzzf1zPe++3lsaMi/05fPSdrBCo34VLc/wriRmBurtdM2xqQSW4HDe7GWc
b7Zxn3y4d87ObRaGcYZGrYwXiPQ4r9BKcKbConQQbakNCusmAUabDj/uaXfnSxM1g2xBz0X+V6wG
aaQIK5Vrb4t6U1s9UqAkrm4Vx1Q0/MIVG9QTZpAlIiaigbwH5KzO5KSwnxOpYWcxJzPtFZDy1oTP
yNGxb64elZzWnU2Wy12UXaRPLeApJVDoVBiQNRmpwsCBH8lJdtXkHr+qrrZ+ojlS/a7XRk5hXl1P
0ELwO9SGaOI7pvS1CYv59rCTxe04stsgdYFZQrbV7xG1TITDwoEbsiO5LWNldHUPzqQXoDYWoUZq
/oCA9l8zJpskC7tVrykPsnDpwYfgBc2DlAs/8SB5229oDRTsvAjhRV0kqp5IB0b70YL1a13OVemL
1JxUhqzLySF88ZAxUHvobMx+RLLPm8+uNo+AxBvvku8fYvdHViZltllETayD5IpkXxxx4QwQgyiF
L9fBgNbENZy88k/0I73lSdGfySHFnnXNCMpYpHpGYVkZTX64x3k0BZjzCMGaCrPsgCbKtNTc6PrY
x3flEQgVHYHDav5zECOiY8Rohz1JL/Q5J3UbiuuX7SvkgHQmLWkyL1oNgMk/PJW+cG7SfMUMaMAr
oXvWs7sgT/H9TP4K98czP4edCximlgFRbia7N3HIdTUKlCLpcRHHrp9aXCqEeh2Hl6q8lydsmLv6
vQhAIJtJd44PsR+IO/ioZ53YUm/v4D0ryPSXYKfmE5kVmnXo8I9Z/oLUFEWAo+mNSwYCD+U6pOml
L+Mc79D00BvwfTBlS+I3sPP6qxoH6WPl2jIHgqL2ZKN2txYTq3GK8UrcCuXaXdPA4UY40mWLZmsp
oftkaTfHxlhoCq+22mNYtDQK7wiEHstqVseMtrtAEfyhvsho3z6Pw/hbAEccqULVg+9CF4kaCRzD
OxHFvSHqKkpHGC+kK7hEWNkDyQJK69R+SgoilGgsky2hLhPtilW7NRy7grCR4MpatototyC97S3Y
7gmwLgKjUEPhgyP4uZq5ONnIdLhO9mOKFKJtPIZ/1UUSKQPAcxNxQ38kuiG+tO2FiYgRwrLDqVbG
UUku3/hruRaKZ4gv/5YifA9ym8sfgKO9vc3Ie8e4uUgg+Eyydrs6/66+w+NlKMLms5AusB9Geo01
Dok+81ox2Qk8BhL7rj8TXtgc9b6OmRUQ6aJM6hwLiygqXcNZq329imkOSHlCrh4fSjHhL8uItG6I
dVbfCVHO/OgO1/oeTE8SbsFVl70NwXE0q2FhgOlXUYktL4TMoT9YxlIs0OQ6NiALdIxHGxqsGDUU
D0hhPL3mAkGaXBBbhd3UpUINgsT0Zxmw0EzcdlddNTOuHq14pcyRDVI4e0zuCgrtC9LKc2aMbMEP
rmuLIW3i3jGKvWbJxGg7is/c1V2hyBtUaJQ//T3yiCtj04nrsUN0gjdHjVkVgYuvIremGYaJGBbY
Mz5lGzL3k77tP5jQaHDdYZPsdkybo8QKqrkFPppYDVxHk4vMPoigsPyLgidiQFP9VO7wYtN00HYr
qmF2Xvuu3TL0clvRAHmW6kO8m1slDxgVsxSzSsKPtY38aViDyl+o5Vjg86KlwP8AfQn832rzNo3u
g8/sCaDxBugogk30FwU5K/e6kfkX+mqcTxI2f8cNsVhVxicm95ZmZi0UQWUhJyTxlqQwzkW7ko0t
PSk/vZVuSFrMzuf3rddZQXmsYDqJTEC/Gv+DInrCJa2LoFIeS/SgDo8FeEwDI8YrbnAZFLd+7VQh
C0rDVmbNPTkkug1ozUPD35XKoCXypFBo2rwZYh5DBJVEupgpqulOprILk/99RpZdT8E8nkZNBMJo
8cs4e1w/ngWVS+e464jygedUGc6zm+jsNPyEcQGQEyPBi9TWkfM9s50gCJYtub+lL/5nFDUqq8rU
a4aJgffyPPNH+y927PK15wyQVFt22Sb9THznsgTkAdLWLXt/WjzWavX7I82a1kqqz4Ods+3LFK2l
azvZoOzkqcDXsF/C3I/C+zsBcPaIjOkDBCAhDA6uZrP3R/8nISKIPPgivRmW8spLHCjz3AnR5Vkc
il4aYbraznJCnnoIQtB6WgbS7izSX0bOhN/Gmu9Uu51LuQ6shCTfxkCGJAt/xuI8GSsV6PFbkth2
EbEHwuImZha6WOoGYd8l9XfcM93Ed29n6buxBH/2IYeykvczsryIOM4qZQDGNlyTGuKjhCUAFJSw
mZ4qThbkZGC8SLCj0yobKK5kI0zplvkO00I1P0EIXprOHk7UzbR3IgJL76N9T7V/rC6XW5ojEdhX
a7FFreg21khy/xiU6iBVnAzhCkMDEYeuOZlrXEBO+EYfQZe4siTdwEthYKLcWPCzoxY2nlatosZ4
m7Gn9Poju7yBFZpQ9J2sK1f4ug7R1iloNlTVWcqcgSVQ3d1PZaGo1JI+z+D6hfsJosfn/grPaWVG
Cweue1nnXbFzN1sCm4TZ3Sj7DJ1kby27MEwFTikmqYPqMd+mo6uaoldZLoVMcMtuMHYumRjL2ytb
P4i/2o4P5x2EkiUwDm/r28w+AG5lkoJCrzGFgo1G6qyTp25l+hbrYVUATwYZ/jzjKUHOPY4VjgEm
ZhmFc66yExy1FOewzKR7ZthWJbijuBfJQk0lxilPsiBWtDexW8zWNs0IS1PCZoDpDeNz9ikLL0lt
emk1Evjbb649m+U+zBHUJsQX0QUDbFSkrwA4TXc7nLPDEtNO+VwGuQbk8g1wmEvkFcRkJ7cqkZbJ
0VwZixOoyDELxF8E21Nyu44D5+liPitS6KDHk3XN7WjRh3ZbgiDch/7wLNdUz/DpXCvm7FjtsDoR
eDo2wH8IGfsBqlAsAGloNAYELykLqREGnhTBLqQsHtTtLdNJx3DHHMrjck+82nHkh7x/dAWDLDbc
WvG88fGoSNeDnAwYAuHVzXhQdaVztDsmOr5EI7sy7cnAPsUBK3FS+0+1n0Tha5bN9aHMBCRPtBEB
yJDK+ATnwPgco5S93etNAsUSokSWAFKRG5hnsmD62oV+E775MQQE0/o2YkFTyWlIOXCEnaPuCij3
CBJh0JDpGeD7g9wa5czy+oUzvHk480XKyvYjHZ+UH/88R3wraeRl1HZO/ONeaLi2IX5f/W8mH+7v
dpnpVm75VsqIXBlpE0seYogRacKy0hl0ML/O4WpioP5SXR22yY9ApQjAtNiXhFk8KcOze3+k6xR+
3RMILDEeQ4bT1JsnJcEJ0/r0PI0lYWgzTpBXai2j8YP1JJ7AIhAO1eu+3uEicUakzz7EYI/YXvBV
RQ+YIIR9SPE/IZ6w8v21htVJwySujVN2wVduSVs1aFseZvd7DiRk6ZuYEafIsbSYLN/3l/7R/OWA
60haAc8F+T0XXXTdUb6EEsI9Q3SA+Sp6Fmy4EJQ2MAw93OwARDDX0ua/0BDn2Otl2pa5X4xDO7TM
dTXUbZPUhXVqghVhGT3kFhDg0qvdEhIRNbDNz1kPxaHiA/RQfr7nVFh0hLrJ1B7ISEsMzKlX9PGO
1oLCfzULTTVVzMtXo0HS0hVLaC8rO1zgg2Q1obLWbelEwFTAx6eapfkuQtAbeboHsksvdyXKDVcr
VOFO2mNIbCe7rmygFZKamVz7RsmznnOh+xQK8h67qVltmvIOWsnRK2VJrXesE7r1iW4Zh47M1Fla
HML96BmjRjim/nV2BUihJbyoun+7VXWePPnqhMZevGmLPy+EVCA3MIg2mjtY5wvNjann9G5Bk/Y7
OKXN6hk84xYdCPF+9COgalqOxJaeAy1Nbue5mXoF1Owp4qHUzpBw9b/JrGvnLed34Ofk0GpT7AyX
u2vTcoazFRdv9Ug46i2HakVmz8EHAhW93s+SyNY6PXfApxz4gnTMXdwxk8VOv92+smh9ilCQnAyX
MU+8iWYVF5uat5TBAbex/HhO2XFqVR6fuRh/xCUSuWu2TaKKA0pgNbfu4DiysT5VVcTfxR6QJPw8
2BnRQ2Pn2i9A3ZR8hn1ji5834qzNKlWciMvg/EPZ8fEV6KsOvr8g7JgXIUnVlJAUxM2U6+0WS/64
xfk/WE1PhIKoRsVXzWGFgoSoOhrsGhKmxCzZjAljB9y5y4vLgEViY3LUG2d3DJ054uY9+fwkUuZB
fh7iXcd7kBGqmhnndmVFibEYS6tjdkCihj+rB3K1d27+TH3XRv+yZghQ+j+rnK9Rk+X/joIMvTU7
6eTWVbgOt/E/w2eDUUHkKYcszwXx5F9SpO3p65eizw97uuUlGr9PW8WUNlYNh4Dus7tchVSNwmB5
3l47plpjRw6h8Jj1wpPniIMRNwsRGOaSpZAR+FP00BluUgxi7OyBbNdB/zWgP9JX1d3MccYp9h9N
WNVDRP0O7A1sC4qoQYw4cfWgRyNnO7pguooaJbf2F74pZtgnHx3T3UFLFjpoh721psbR51fY97s2
oxv+tF0mHEzmO2A5nMCqpWRVD2qHkJ6Ugp9R0QYPGt8W23NZJBhXNmlTwiFWGWwfLqcchdc9Y9fh
ev4HkBDWjS+3HYedmQnuxNU26Hmj6RbtUr2o0CCdiOcVT16jjYlrLGK2rYAqqBR7dYqSzbHyNc9/
VfbdC2xsfnQlMEb/iXQTvJssO62iD8XNEzjAn6BC25vFHt3k4iegEZ5fkONpkdOkkhDVuFHj1vLY
WEUgEo2mSP1IJbdYzivsr8HWCn1CRgDg7gMSJmKR5EEAoYX7vKaYr4LmKQrDLCNwMSwO1G5DTbrl
cGBOzbbwdiMzng8d41TLS/Ky2cBc5PnMJckiEpYgX3INyUV1Mf0PI9z8xmgEyYnQictjZ19zukJ2
jXQ/CcAJaOal9M6WFSR/ARX6xq8JjjgH1eHXoMgdi9+JHYJ8jhIkq4VbyQl57SKd68XXbffzQUtx
+HeA4Cml8Cqh3wSIubx6qCoxTZUJGiKDI7o3S0F5gWNlk1ycOL+PjBTyu7kamR0sVYhpti+xLUun
DapdprQNz7QLmUmuSH1qjR6aEsBjSKo/14vcvgzROBoJ5WUdVHFGblyLp+O4I3H5EV2lqwHUSBHM
KPZ+xf5r4xBHgoizWVsqTfIRvkYB3uqF3xVUp75t+Hc2a8sZC/49JwU659dSs4Sv6qKA5heek3hy
sOs2JQeb2w5Rc6ZcdZHkZEyGNdRxJG+ByeMwVk5WVgaPIpTyiz+ORtzkLwgoNjk8Jl9sif+MciDZ
+3VA2H/Ug0cVUyBac+lp77fXcBg8Q/OwUyo5s5zD4OUQfxpz0ldCuVNr8P1wmHoU2c0afNQbS8Ec
0CaxcH7Jn9clIkRPKLyZTSiuLGSss8iCvPi0T8ZUwKC1I78SeUYxTOjmJoR0mSNqeZaMMFvGjXn2
eVlbEihW0Y7zCl98X3Hjv15pbXWhvgmDTRJ0HLa/wP2WQNq8Izk+YFHxQZVDNJwU7R5E7n/fPqqg
lXAQ/VvIbx7sHv5tTRbWwfB9yU2vYcRhthry5gF2ruME4nOyhrUb7wbM3UZAuE8h3rlL4vGBLp3/
Nel31pCLFPt24rn+JHxHyP6tNu9vo17Fl7Ut5isIbaXOeYZGG6TKmz+7YOIeYYECXbRnWlEfTZwj
REWmnC56Kmwy3ttx2oBdnuB4lkBp1WfNuScI7CVnjUdkmUA8QEkdZ4A43RTNuvl8O+vC6mKEsm7z
vyZLGfpurSOI2CBCDT3qQdwQFpQ1nwrIzoDo1R5TBpjKuoEc2WysGiuvYieakkKb/qy590Ma1apY
oDTSB3MjOfPeZW/7uuV07FJTlmx/7tHzaab/mh26xqMJHU3P4FpB59tydb7VhD/x8uZtOH/rSpPs
ZYPMWiWXSosYOlnv04GTuAicxjl66fn74cXSiyJfPn0EGBsJAau4fuGoYv7HVULM3PwPu1ASneFB
PmDyTyJscEPt9pRVDJjMJrpOhkXvZdf0w1zFNeKiPfYQkBwbtU1EHsz+sa2ayLyQT9vrjwAnl4pD
kTKpJlGhI6eoT951+wo0q4TNBxVvmoowGVQYHlJsURc6zflZt2xXoH4PKrSlBw4hbAtC8sRj7ah9
1KH6OcRFGXlE6q5Ai9/MS9wXRBJ2Wh30cCIDB1PhKEjQ8AYWpFkPtUIiYq3T1iApxU+LvzhrfMvN
BYf+LlWM477G8CcJgcZirIarzn4Wfcz9vay3A8ayEfmvDNGoT0BO6vWs4HV2eDaa31ccsnqvXjWq
5jNrrpqdjesfn+M1IxaQqwbPYHuAbsCb8qGyOIQSBvElTqb8RScsYnHr0hCGhMiFnm/QcdTZMrdr
30Of2C0sksl1SOvcOgt/ghG4D6Ec+kG7HidMQPQbhAEDBjMCKU5UN56/nJKMscnCj8BeYuwvNXnK
aYNMvoF8kcHCVJwE8sjTacmNVr05/BNdrnT8C2wgmj45XSCqljDzaW3+5bEthyqBxwNVQs64d6UQ
xKevwm2v3Xo/m6UkrK7TRSg3QvNa8Fcq+Pg9GAw82FKG/3q5u6wHu4f9fDQ2e9MRRydB5W8GEP3J
ySomcGxCYTtHfPLcQ0I5zdKIsOpxwm5NrcLb1Ch1VK06Devdx+AtiDrwh0FLhMBIKRMnZguneiwb
IN0IwRHCx6i6uwLNy2ranIpSKr/9TXEHKvSDVqgDszYsCQtoSeBIq182yuXtMDTo/pG4XA0XsSG7
Ya/w0U8buyOFhsaehgJVKJP0q7tpPusux/ZFkXCbJneds3tastZ2IcIo2lqBv3Nw5YtemGp8Zii4
FTJLH9s5YU0Sh7xE6OYRUqtcwSK5SQlUXU4BzY4JmGpnhMXM90VDNmALRrR2uXCzKgHPywer9dXi
Ex/v5G9r6ItIRhe6E48EGxWFivB2pjBpQXbLbh9XvHr2aRpOGZ+bTcIDbaoQ0ZUv6VdbsJ2JeZjP
ik+4fCzS/yST1y9OMK4ca+SgKMltpnYRwGgGr3d9HTHcLP+N9yK3+Kt/9dbees6TIDfL25kVPiQF
3w5htbI9N3zKlofxMoDvJcyiOjcYgtC8QxhBPoEWcPx/Io7eACLX/JfCSjr+Kom++HQMFEx70Tse
0sK49rJF5ID40ivUzyiF3TPopvn+/qHuYVXl0HyO032T4Dh5PuJsCU+econAnnjAXfUFoD92m9oB
ImEYg7AsjqY8FCSJ0IsY8qixY4ECr3MAX+WcLiDIL89aahyfhgqz05SO8gEZ+5nBgmTWYfs5Ksu1
kPck9gcbg6g/2b2biS0RuMp8L19hPK7OxVuQRl+u7gZ4s3YwgQqA8rdy0DM3gz3bRlycvORb1NT5
JuKKtWK/E9I2OyF41jM7Iuimn/69WfrivqVJiXRG0Zdq8tKk63WNoKoqY/AZc6lZ8VKr8MTc8Yct
6G5T28an0rqAXTBLdjGNQjWY6oUtptqnUIB1LZxgetp9uOLqX565ehZJOcb98hDFI8nPltJ5UML6
jxK18tIeQcYNqRAquD/6HurNVFUyYdV7nuIt/BlFaoV8zBp8ons91rqmg/8wPkvWbNxsEU4tonLA
3RpG4KKwi8THnJABHJPlAU/STzlgC0BJCOH17ctv5/GxHE7fFsYJaDjQ4c8Y7s4bN7F1pnfbnvun
AFgAfBmCoyI/badsiFob4pgTuIRyXev/fxyTRqSWj1simsegjzSleNOT09HXsUWK/SFK5/GzATfA
SJxDHIlEsu8NZIjmJgZTfIkpZbplVu6BAFlCQTbTknq25zHn9W665JQkPTKmIP68gLkJRy04wVZ/
NQf86chGFzj/vB/K6PkGuP3W1fbddlKzwbRpzvXxGQcEnWk7EGLdFaNnWqKMEJOn6LWnrFDj2MZc
/aRevwG4kzoy5ThvmJEHR6ivEbhrSVJOBkhJ97wtPMXBozP9pde07bQ3vKezOai4Hnf3BzbAHUcg
ux+Md3p4TBLfg0v7Y5JbUqtqvAw+1OzF3OFOb0dFB/CF+JqUYimroFaqaUqiTpnb3icgN/DXetuk
6OApW3CbObe9S1ugxVFQ5ANbV+d0EXb3n6lwiRKeYOuE1FBOB5EEqZb8RTrkcIksxI0xAicP9XqH
LlTIwAP7A81F/uIjXuDo/e2hLPzo3Rj/rXoMMfln0V9Z7qrjhHEnLR1K3SCTJyEFnACT9oItb2Lf
/PZ5/G/FFltS2TuL+UqHWDs3NITiybFDBO81pXT9MfR0tZBan74DasUTFI3ieB/gcTOSWMacd/QR
THzKWrpplY+rrAvJ3Mx4oVgmKhtqT2pnlwciEdBNr5o9Qk4VMzNuiJI1mvtLxVl27gxrfzE3okTU
Ex5TrNvUu5CWWn7WgaQ7Macoz24w/H0gzdSu1dgB6dolw6CTa4ZaTNPM2AcGyOCJj3j5Kk7HoS32
vK56F8UVJecr8XFU/O43nOg5hGR6XU/i/CJvI009jbexdje+8n3qbBVZApbcPDslilaQjc9zSgWl
ETPaINVqeEBqVGRAPH5iTCR/ls8+7iwgRuwRXYFvOjmDB8hlDoHn5pl3sMNrqgcKAt4SykayjDfX
UI7u6lXw0zcjlbhDoZnyw2kLyEtOQ/j0i1fayFkLoytglOi4Hrk78Z2VQhM3kzMt3q2Lz+iQ0Tl/
N3MKEZjvCJBpZBwB29I9Wllo97/X8/RlaBNb34XJxT3PDog7A/BJztPHJKEr5Cuf1yIc/UiuA3Kb
0rMl+spNHEib7MyWBLQUNGak2mCtUMTf+Eosf+LlEwoDWll4/5i0yBpl0GC7M1mzPLDBbRL0/PkX
u3hM8Fn3QVNj95pQ/30FL8bbVYf4fMegQPMUpQWzMrrberVxEty3N1+vmRkLwHiBBVqzDiPVfMFM
AChKsyx46zZP0Q+KFkVtwBwee0WetCGibIMeHYNtruiJgOFyLaksyYT7orPeqaP0y+YlnT16IukD
mypaP0A6APmH9lDKpTVlXFQkbYuSyqlYphb25p5/JjUeEErb/nOPcNqTm9pP8ZG6+qeo5p+vENQc
hX4a7IrF44uqcsWR/tfquzMgX0SHch8QkQ0l6idHcEZ411X8jdR84VNTadZ98J2MNU3sZqqd5tkk
ZVEcwh0vzzsZfz+dDCMxHqD1R9V44HJPOZok0O5ClxOcVKE+94mt/TW2SHqHmCFoIiY5T6L7jrUF
QCVyrHVbjaCc9aFKt4LVhjKpqKG6+lcsbS3mtIJ7beggdUl7Wo6liiswRBFHqme3OCIWhH0Vn8ZH
RU5mly9Pxs1H5WdKG4AY41me5gS7YjxRgYmItKA+FpzbEyOoZEJ53y2kClQG85XSrKbpYSgynFWj
rT41AWt/5NxgWxko7y2ZuNrYbCyCuI0QeAKed5woR8jMdeKsVkQxFdtuxg/UqYezc1HmvXeZZTBF
Yo/kpkzhWH5eVI8TMRIaMucd15l1zFx2c9SLTbGSK+4/kdU/qg/2mhjrPR5QfTkPwREYCftpeKIm
50cO1mqu3brWhBaUGccxOcGJFJIMkddhcYIijVEYqC/7TyT7LYuzoZ3YYd07nF+GgFgPfwVK+cX8
x+tCNlI8tQnNTeY4Shy+t69aNgvKoTCTK7F7MW2jOaBngfG95NGQJu7knoUsOYJnrQfCaJMLEUad
GHXhUdGfj6ESVuwJViciNPCUdT2+CJG3FLG4Cu/0F7B8xUy01b6S0WbpP96flm2pXG9cJ46oLavg
0KzIypRLZlsjq9HHvWhcITmZz8xyMXx/PSC4aoyP2ADwU8ymNQzDirRkLHTTD/qZRAX/IVCDXos6
IRZM2QraMoV8MLPhpx+0gf2xy+pyyfVpX80uOUUgLkdZI3kjtomh/HIVYylCJ3r1ygLa2MSwgDWE
YXyi1J80N9+j+tQzViX15sjFpbppwFHcaWG68MXOUFTx14xsE/tsZJA+wqfCvsSnogU/OpeeLKzY
6YV4uGLlhoymWYTc1m9/j2luo91v4kErmByKkgJNunW9DLkzsVIDjxxqbjD+sYnJwBWniH4KMP4n
mw4Y88Ikf0E3Mg27y/7P0XezR+kcfuZ7GCetmPR0p6eMha2WkFDxNmh3UveV69+9IrZcKpBUs2Bk
ksqxd0im9g0TC6rh6XZUSw73fsLBgn9O4PMmJCYlIlUK5EWoSFBhJnmWavY9HZdFUtgr8/AoSR5/
FPuBntxkWBS4ZmRjrSSocSA+ubUL9T7Pz1K9KA9LxbyTIdDjFtbX3Ag8oRw5i6IxbjEAxiKR9yzl
gHWBIGFUNCHFB+CnFJajca2Ctz2hOfj+7mOS/dDRDIM7CsfnsFj2Yz4XwqWQ4DYdq9SM6ySV4/sP
oVoSYCINCsaMMq3mlmFJyc3sZjko1tK+0Y07JwDXUuS5S8lbZLcY8QVZu/pSeLba5sUykMX83ofv
GaogVVcgOvR8CUk3/rcFb1sv6Ty1f+ZVun4wnz45x1RbvdreVg14/I4AHzqnHZ+tU03G8oe5WKov
CMJCC4wRcHJS83Mun/wMrQRIaNX2MYqTVrqysEsuMoVf28ynNpAo4LIemM1u5Tu+8nSTB/1S+4Qs
NRxRkskkYl0ou0ILjCPGGfY/gJ8k144BcAVqVZVdiLmb6YjatoitLJDG7JWtfiFRkWhJaohx4LHd
2yq3297ns2XxC1ePywjn1GQloUOHqDNqfPRyMJAZJEYXXnmVHkIAi3Ny6DfymZ+2ppD0igEqrfrT
52IRP9T+Y7AMEE3odN+DDNsihEDf5cYCf1NtWJpI80jxKTXKrh6IASjZyhQgODNfB+RJdtx8ZaWf
blSGNwGdu42JpZwGwhv7Aia7Q+MddLJ9yjHCtwoAjWZbpucKsjZLpiOs4bAKHYy0FC90Frf5Ss+s
EebEoKY2PYcArPMFoPX/S5yTjL89YY+z9YbYwloj9smvxuuepkrosbnDFbsF0DUn+f3PxNIAMMHO
w2K0XRuDbiARPnO8y4u5nO8OUpzjXams2HyeH++GwgOnAZFusTtJCaVUaKtwwsX+YG0XTaAgQkOl
Dikly/hAj/9aQEJn6JwVJ2qWlbYJTZDshdkguvYko8BZ2FREnoWow50lfS4SDi1uvf3Pdx+QdE9i
XbmdJ8Y1S6/gdl/rh1F2YTbp4Ynrs6CBMNoX/BFbM562mS4IAwgVSZ3RgW4HMlDWWtaQuhMC35RI
c7JN9iHnDSfle7xT0L8sbWMexQnRKUFmNfjGWe6Vdcph0SvAmv2Y/eLe3M4DlVrk4zS+WbIESwMg
ri2WYzeCmoS4NFy56594ypLPDW2IizenjKMXH+7aoR8dhKnGEgz4gbLxKJFpgwbSKx3QIJzYfnGq
TqLmLbSxmUHQdafX3mK+tugu5ALwgrSWhiDxsw7yIfoa1p6sEkEgRrRG1LfaO5pisv9CaOj5FmiO
vwQrRUo6C95ZcpxHaqgzzb2NZFAa9/5FtTTTzMPejilpWIU9T6+iBIkzpJT9pjWQb5+40flfC5It
H6t9z1/WfvUJsBvQWro7UBKUSQkzJHJ0NKPro2mWjfT7Zx0uKa2VMmoTuLinkhaUeAoPn0svrb/E
5yvfMgq45pB1/hrGapTLlVnWFhqDrAlcwJnjPHKlVsfk866ckrVLvw/nZZTWP2uCC7Z4o1r/evv0
uR+XtMEepI+iHNZ6q3ZBWzEk8x8Remowh+VWg72hgdZD2WyAoZ8UUrYYK9hB/gGWFJZ6t6RKkT/c
0kvDMFQmueZ/zQuwdm6KX7cHaeZgdw3NPWFKdcNV8+tQ2UIJ4q4f2HwT14Jr/1dzecdYFxDq5oNJ
1oGm47jupik63ectoA1W7zfvnw7heSQxhZbENERy+G3q/a6sgk5EmUbvRKSVZ5V0Ii7yj6vD0CWG
RTVdM01a+lTpgm+MTUI69rKpxlnO4dKA6P/pvbJ6KLr+2x582w99nwtR7ZgrJfjJw5rKD5K+gGLW
pFXXzCif4Jr7FnqkxcQutAmCVO6p/Nk+DbzyEeITpHPXKCbbsGv26KP2eAaYQ2M1/1zWQLBBXuqM
BiKDJVvvq5IZeX1Ln9DeEh1aZH0UCKiL7QFJHYK/7sdG1qTEH9bNCL3it6wjMe2vM+v+/pDX/dtB
2SAmQmUHPSLjFrd/afcEud4JxkE0XW8gVRGcOWkGkdr8zOafDSnW1GHpwxkTzw0kSxdujdgmcNsn
GfXIEAmxOznxBW6ev16wPhwntI4K1kQkBWivtrm5cB8nfdtBgLzNcyhcnqtnx9jGsIb57lItLtFN
iJUkxPY981ZHq5qDOR0HxLF7bD0glnz2K1lkvD+PapgRz5/4NZfZ+3xaQTsJiJzH526iaTKfd7O8
36s0+z4QfazHkyuZwJmhF22xL5TCjTuTizkdcuSizagwHWuBWvBSrjnBXz1Kjxof//ZzSj1aEFlu
2AOtMnblcB6uDIy4kZJq3TrwYH6ItWCCcTbAblylSTHF6E6PZGOZHZhKpsiBzHduHtaIFUHcJ4i0
abCRoYoq/MBeO9ckbZ0Q08i92D7GpZc7FlwUl3BlarHe6IlIBYmSuUePCgmzt/Y3AaNvMYMUMrld
UQRoklcJqmMt6wTjte+zEXILCQCrG0CrMpqV7VbwL7Dg+Cf8ASj5E1ngTT6BhctkBItP/W9gX1Ow
8k+HbbVIaBE5gXUODL2b+sHzYHQ8V4TZEB8CkFxYTxUfqHPX84boOK1XAx3kO3QBUObjw3b25EeR
Vl2p+F6Fn6bVZrqERTsRaXRxAS2XHNHkZs2Ai4OsFP77j5QrSWh2CixHa6akxx3Dy7V30HugtpJZ
W6xAlgG5Sd3mBtYUqcXlyLMDjgJ1KXAZ3CM3/q03i+Hrw2aDdi2lyDfKMwptQlrZTXPmJJr4zVhD
+jesg2zKQ6QE4fD5Ct2/6KJVNYf8DhBGF5Y2vTpKjqqelRB30XdDlHqDR8lqSD5GPt+KAWDQsCmZ
bqQoe3Re3/8ODUW40suJ/YSKAIaddVCoFvN5Ezf2Y24tJsg8hkdoLJEgm+zLM59GgazowPdsDeTM
EEOG8i3C9hNZ9/joorkxCQHFIVgHizu6u08cRWsAh5neL9vfxx/aLOeuDdK2sL0tcqdreRX7PBuv
YeO8zZSFppzaWbCL7IsirMn4CGMf65bmqEC1Kctoa8LjgBduqbajKUFENqYZe9FVhZXlLrBzXtUR
HIrglLbpGXPs6SwHaPaz2fXGDCZ3hYPPSBGgVfu7x1P1DMy8+S5Gl6xkgoxc40728A9ydIyKvl/t
s32BDzkl5v+7ToyQHWA8npsi8gMKjBy6jBdsnKUk1q5jJEt0bH/a+2rKqDamT46L5uiQ8IuHlRlW
o1P0bOW8QxOdBX5zQChMIC4XMpdG/KjQVvGhGf5IdDq3NN56bHy7AEI/1YBS4kjt/qZpyMyWqQfZ
M59BJfdQaRrlKqp5qY0KiIvYtpq2VKgXbYA8DVI8UYSfJsWPbfhekZ/WnDgW/wiysFc4yw9X/qbg
R2p99W6rR4Zfcu4NpsnisM7FvZHofGSeD9PhH1uSNB0S+MtZGS5em3jktyz98feaBqZrgfisp2Kx
c0ESHDStOW7ZBvbAj/PtPx32HOWfnlzbDlX3YzZUwrtLUVvtCtNIfmjm9bnggDQ40N7giw5QlYZT
WQ//0mxV0OZptgpk1hUx4wnecskBRdxyI2beX+CsyIvFtN/V9Sd3HBiP5fXD9hn9kZiFR4GWXxZk
zmbCX6taaPVAHsgeSef9Jpfy7mJvkRSMwyujaiuO2eIqDY7NKSm03hjDZHqHk4hZPcJ563EXw3vg
18X5HwiYmlvFovrjmWhTF9uYzou//yds7EC0RRQJGzpyZkr61AEQ/b0AWvpXWXeN/RQh/FM3cqVA
STU/oj5KsHt6EnmYG/QP1tOYbGl/r6sLDpTucWU0S+fG3jily7Sqg5+JqHSqq2ixR2QWGLXsHXF1
J505+JWOEzPHwZjUklIECmdpDjjlo5xY1p2bxI7r59pzliZX5Ddj1nhZ7Bfy3+27KZgnVDVx1TNm
vj3aqT4BUALViBvC8QcUJU8ri/8MxLAx+3mxRBOAGQ0IGg6yWIaU4l76j/3yLi3gXTFz3e2K5ctO
hILOIPNJa/u9dt7tCLVFjT2FElcRDbmAfi14P5VdJMDjpP9xychP8ScbInQssmK5DTdvwYXnL9Or
NKA5LP5m4W2crkazNvGYAGFBC2z2Xl+IrdqhhexzJcCFTxchSBR+FNRkvguizenCbxxANcL4VU1v
Lwj1z9RUiA4BCwLe8x4vIdaTvWYnU5nUFhiZU+v5/AAlkF2Doldq3M5OkRMDYwv9JAeNV7M+pEDC
ZSu7PxZ8cBohnDmZFPXuRls6P9j6leNBOIiarfrNvOHFxqasVIFLMhaFvb6GjR9cAD1zFQaSfi7I
t9Ae1Sp9srXnK4ewfqC73KzF9k7NxhArNGLRyxGwi0LvUHzxxn+XM52Z4uWSbPYAJxD6G2e69k1w
arcKCs+TufHxVdCWXgTBNdp/6fnNzYtHAnDKa/uiaEvodEPfHdoFGwXCZ++FMqoEBTDyNuOjXZXB
NjJMrfM8WlTc+zHrKYhxuUcQt6ooSL8EiDjl0jLSWIVd1XlVCRd9EjjiQc/i/6OP9dtKVCHuZQOx
wCRC/PRMOmW3l7M2tM7QZPe9tYv1bA+KTnILMrQJWqGJd/mwohZbNHDAFUJ0Hnjekd0EeEYnvVez
/tEjloBmALaiWe6ZpbpSTHU3w3y3iDFO8uF2Ozcmvq0Rac5+4uck6wMN1WLuE/h04cEj1X6k2Q46
I+UVX31Jq61qQ/PNYG487TA1u4NSCdfgJD66SLghYYv6A3tVtB/sb8a/1tnzb85L/hLruweZ3OUc
zj1LkqBKRZ8GGc7xaJ4WEurjVI1Fm8QXKzx/2b2I9VmHDByWighrq1KeLCfrgRAkjuUaOiiXa5ZD
FcsjjusVVVml5zxv4Nm9DX9ZfSAd4Hvan0aKFz6rdMzN9cI5tmIsWGO9caX0Yuq3qmDys+A7l6mx
fBN9zS/taZLHvuAoZwviU0o4dJnofdAILa90rMwjlxrmAwko4l+GZzOOUJKbkTzIMR3tTE4UmHy6
M5n8FWPccGEVNl3tOk/A4p1oybub6WHepQqrtBBdcBPpYumcmM52oqJ5xs1pD0BBtmfV9xndf1Ba
pXAfnmwEJc0m8AOOa1jE1Ob4J412cPLmjzDTk5JQF0eLnk3x+QbajTmv+SXA8Z1vSBS+gtkngLWZ
BFvwL/8UCRmAXpfpASl+t83JYUf85JfV/ZDw+iFRxqX8qfMdqylqGlq1I4MBNGTDj0fLE00Xm1Ie
pMGOPfHPPwYtND0o3228iVUN2acnDq61Y/++FNBxGfuidlxwMCI0R78LknZtKytjhbg6TMeEqxOw
EEHkqTtGTFByGWMru/KQcmcIif6/S18ZccEnO0o74oKKDsLObryLGy7szqeYmrjrvLurrytcXVdY
oBCuT2OpQg9xO0bBiikdlOsxi87EZ0oTfCPCanWIw5BxYzmoR+gCviWLHOMmunLsQCojYbW66DHy
ogSLF4H1MT4R1dqCViX4hPOuVtRQVwKs3lDCR3d+7RcY8hXRETFSfE9Di0DqMKUOGqj7dqWdiZ/f
hz29FkD6r3H5D5vX3esoaypossr84AXi91+LI4LEVrSxXtjTBwGyeXtE+BPL9aZNZM4JTObi0Osr
N/xzvJ0YWjSh+lq50yEmZwjv7r/LJhMrGz1kPiKTBQwMwZ/ipKCddq4mpGLo1ceqSIndfwouvrKq
M9SxvuCbysWBQLOt1RtJY2hLJdr71gnSJFEE8IxEMVjZp0RrLuCWRxVVN1835jo/cAzlu6a57tos
LQmKxisjaIQDwcigbH+HN0D1JUDDYsZgUzJo+qPjDJJnUuaFLTJB/W556QOEha3dhI2YRKxfu+vR
vkD8Z5WFP9PGmLyHrlkT9WkgNCKAB85p3U0uCoXlLRsAe8LI+Th+ZwMfzEzpoQxw2KZxklc+S8cR
hhkfLP4iehMTEv4ZEipbmIc+6IxwT4bisuSDPLD0SeEzkSQ2S84ltHLSH2w94HVDYglmiFdWSN7C
p3i9cM9KztP9SKkKy4HKwBV8G0qhZ2fHvDY9Dk0NJMwePe3rNcZtNziXqEcxlSwCHahtsJGY4RYq
2ryP3VF/tQwQ01pBLI3TnE6oeTzyNk/l+Y4c6yFQMLx0wiodnGmByFtvFdPFcMngSPIrpLP6dZ4e
gPizHGjdPY3d2nXAkaqywaQvHmNXeHPFmASRK5+iGdMXKjQEcV7+ybWy3ce/3uGvy8vMqTjWSah2
+NhSKnbEFJ7DgNz3RSSsTYtF1qnqoFGwlBd5oQD8AU88JXCQ7YfXvvZFzGKWeCGnxrEuzPzDI8Nn
ZzYlfZAbg28U194nVjiF2DbYaiI6xghLh/TcfQsKk3OTunZxitayBvkc6YbfRo/ToZr9VgorFffR
n6r+qSHspVvgOoNtiDwaUYNPQmAIuD01YMXOFDt4rujBH+BcUFeVBlatV0GyoClQm1zlIxMBBfXO
5SOrreuB1R9yQyTdAegdOLeY6T8rZhW4P7bGMfBdchKVRk9XMcngdxFPdUTKUk41DWYNMzJ+FCx4
iFLiFGW+wcslcH69hlM7hTOGGtE4LcwCqd+lAQ5B5oyRKpOuyHeJmBFnexIzJBFpb0Drlt2kAQ9w
fDJX3ET/8Hp8QHLgRkzzAgFoW1j+539NVHWTSR/Z3Y5BBB11n1Zajl9fl0i7vMcDRjha0kxJKhQl
jGoh7FUtjQ3bx5QNf5o9akEoJ8vtqi6hvkVfCZHz8EyfKbXf9xOvonupua1gYYtMN7QdYGzIqn8B
hKmad53lXZuIi9en8b9puQPkroz6rcgY3kftNRO8T7Mij9pC426bwAf8D7az3Wls0vdu02Is/NnV
u4KjULgLYUPuRzBPYAAmvXB8zEAU8YUqvAR7LusoOphvUf0B7cEb4pd/ugRSQ9WfYrKVsP9SHYP3
pmz8LieAXL+Bby4da3kFemIkMp6AdB5feLeMIadplGlEhL0VQmJukc4qW1ZWKG5A6yOElXX6G+98
VEKoPpPhrWZQEXuLrgR2/cLMBITSy+rniOjeuEFlWt2dAjpCPXNMRLSAqsHnpBQCiqWbtPytjvZI
QkYjpxCx2usItY7gYCeQaGHc4digF5mC7Ny1xdqF1AVF46S51+ysqdOuG5qNkNqztY8qQAa7NXwI
OMYyoG5ASc+V4+H4fFyJTh1y0lHeOefXiSAPDGxgJpo9AiVSR1u3XAqaHIXG/rrkZzfV3NpiAO8W
OR3FDBahHQ/qBEdeBaxcpnBxsFC6GaFCI6CLa/1ad0PDj0Mj+8RlFM/XfTMtL0b/1JyCZpdfo+M0
CwdHk65pTnfymgYLCUdyih64yGja2peWRxQLdw6ycTKIj+Dhlc9pqhhen5+RJJlZvW82fl2+faib
jmWyw6RKGn1sL5I0TbiAot71aIC8WFaiFkVuCnl+oAr727oYLmprsusF2GYPgKSmRAvAVnOp4lGj
UZ7ezZzIWfXknA1+iQnfsp5hyPt89MxPA3KkTXuIy6KV5lmFZELdfvJDiiOOewRCqalnAA1mAFjk
pAKXF7l406BWzhfAxnp7ZpTcjMmunbsRFslo9OX90IYEBCj0XnorL4Nkl9SHUcUr3ikkg8SOn6IE
U1uVgKS5kIPX3xQkvCr0ctFP5ZaoTNwzpQZTulDFdWVyjVdUQMCVGyW5CQkO5StJbrZFTYJYfQK4
yDuXvKe1uPEMH29Wb+xk6zeKAxjJjKwtnmAZjlA+7qpm4JTIESMaHFIhr2zDMTkTUPXN6ShYruZi
ZFPVxLIKb/e/ddhNzo2mg0SPb5eJKcJF86oe+T56nXOTcJgSCWhQ+3dhAIgg+pYnYYQISSAG6c7U
9rknnixwQy1+DsODjWGWoL6BY4iGNs0SRKTQ0fl93bp64gMWB4V6ZBYjGAOMnqmwL9yitTwWiMZe
huHdzXicJXcC/AmZWYPEeh6pWiZUNfczxmMsRTBEnfB3I4xM43gcNeWbKPZ0ArzZPfUbgvPc9mlb
SxyHgcNIK47Z8Ti+qAC+h0uOIwDSbb04hI6JlxsU475buEYXF6OyhWlHMEuW99Xr4KAKF0xD3u3c
n+ePeegRg0QAawBR90WHF7hcSbZ2om3bZWfCw8CLfzX2HkzCrT1jru2W8domjc8kXA45CVL7jK0i
4LrmD5IKS/b9dJJcCpc0QBkkF6Qa2u1nxQD6LeMdAV1p9jiAwBmvlj5hbsA4hBXVSxk5+BGPPdRi
hXov/+OmAyaJrrS/5ziWe7Uz0TEnQmiCBIJn1GFlezQEPW4BjokDf0Bgf01QFfbsYYSZvvm14WQ+
JRRTsNLZb4GAeF/uO1Caxn+6gApT8SK+rccZ3deRL5xoYt4C0/1s6SuR9Y6WugyGDWnbO0/xNdy4
8IUVJ6iKQp61JQhGsG2wFFLPngLSbguw9GQVma5KymM7YERxyPcTR2QnHd5i9UTk2nYzK1fd0tA6
hjf+4XJGM7dLaE9U+n5yEXttAZsLAPTHU4FZbN/X/SFX8AQDFIwsIy4+oV5XEObZVTTznTTD0uv1
0KZB6I+hfaTgyGQFIiynHEGeHY7XbYGgHxK4Gqtdz6VYtIGWt4/jGJ5Mphl2uZHQNCICv9S5cnpF
cbVIwmi1zZ91mF8BSJxXSqw7rtWStW97oZNHKirAtH5ZQLbmmzhectb4p/xFviGdilRsKYSsaP00
M5FLAAp+jfV5o8Ul5clY7J9vT9y64ypFY3slFbYUi7zPT90vBpppDEX7u3EoSP0bdOvuGh6V2hqz
Y79/jo3CriesPqY7eCQHFAlBdJ855tW1hretl4ujF74Qy/qIjul2Gqwzp+U6rghv7bhxRzRy+s6P
jFuaKiPFA5AqU/PvJux8OWanVZJ9QrgZ6rwgz13TIBnEykpsX6nRFH8aI2i30aSU2oecX8eZzxnM
F8LjfF0dF9FY4zQ8YiGfoHYrObZk219HnxNZKmDFgL2HoJKCsmZyfotsKUfGb9Mm/X+NXKPtiOIc
p6eYJggOGmYGpx1H1Taeif+eTEZUdpczLm6echoTCtLMtOcipYjOTyxiP0JOlO7NbR8B59CGAbo7
OeHOK8wsMeZCuPQXls3SQqcvAd4euXeElW7sgYsb9XlzIXmLTgI6HlyW+Z6ikK79R9Boo8on6lp3
AbtmeJ+waFZqQ2jrWUYaKbspTKNti9+EcvVF7GrRwq+rw5eeblUDImRKQAex4gI0sbuEYDABmCr3
ohAcUa2hO4sUavEMlV7p4v3oII3pB/0iX7KErqk1Oxr3GAAb2emB7WUnT8wG4eMrAl5KkTlXW6Jg
uckaYuJXiG6GKJ4ZxEfmpKgWsrICoc3bHbD5LPOjqF48cCRj+mcrDZSQHcJ61FAy1j4gdsv7qwgH
HozjQygSMhfeTF8vxD1vyGKkj7m/EpDS9zaqyczoHyD9sKNkIA8t74HngqSOZtsxVq5qoIoZ52W1
62HNWEGo/bWkhbsqRBSLDL4Wpc7Z9OTJXELw7Tfw6Z6MogwWtwzvErsHDqqPgQw27Q43/BAudDAY
ABvNQfpTZ0DRVQv2jqerkGZsA5PkWLzqDvawuUW8ToYgodk14KvFpCeB07I+z+3+p7u3yD5BweTa
SSMwBC4+kSpVCpVef9sEXqaiJAtIq36yLNBv7INrfKPVbn4rdy5D3Tr8ViUpODjPRCR36fhRbZwI
ZnUVWkORW2VJRcKDpNcIOX6DUJRYDNjurYbeP0SlJrtl+6cVXjHpVp92ZlJ1Hl63zJIIZtjGBMr/
Q1/KmhEL3HtRwn56sAI1L7DRWpTjAeFjhUABQccaXFCcsMAT6HAj3jMmP92ZAiuLxLVaMnWZVyWx
Zu37WmUR5mmRYnr+fcZu8LphWn6BPq4S10Hdr9DWlYCSc4gZcQhT3RvpsJfee0qhTYwvnKV2VEiK
JueCd1PnNsj5n0nRAFXc+0sbD0KxxA4MyGR/Lc/TDH7bBzLQqDK3gvr6FJnkdcxoQbcLYWLBq1WZ
J0kxklohLE9Er1xWsBjLN5qkrYc5r3AwhxrQclt9A2YiWiFV77njmu+b95MXE9KkjV8xh4/TVv/2
kacVd90L9EMj1YjHMnARq6Tk/EP9i7eenzQyBpNBeLQqM7NI2Wszg/a+0mRNimRrdCu2ZvsJ6GQv
QqAuk8CiF9QYysAeyub/xPAc7XfjaOd7yrb7wdw+5amYtBIdx/k+V11aEiN61LMVOtjAC7W6OVGU
w9iP9+q1LxRJGIhpQ6XtIWRXL15bruLUd1LMiXVkcdeQdyVi9dP1QpW1JP1V80a40q5IG6UvklNI
/7Pcd90ytJbiAy3I/lW2B/Rb4gZasKtZH9N8M7frL3Pf53S/9bKCVT6OV9qDykOcsP1ROeqSP1Bu
s9QZcm9t3fSvQPHQRpDWCRLtIlledqp+j7smmCdVHlhkxVvilgFDWAHz810Yx25hAWdo6oBfTckU
6RA95pQ74FEWhP2a/SYGLfLxirZTWmhG7JnrLzmBRxP1y/uV62NRId5xOph043QIEFnPZ9REnnFo
rwTGKTGdGVoQF107PZsYOC1SrNA68LcR+7DaSJiCKCRb93Hn2F5s1rwpadagu7G9fL3Xutl15u/j
AsZvtvt01ac809mHtbw6mh0a2SUPTBrc6Y61RblDEYd0ZTiFoBxA/OVKx8JR/Ft04nH2mWrLEMgC
BTimF99cvGPU0P/vN/MIxrykl3GFtmX1fombZrtU+fZ0v2xrziw+Mu8Q6Cg0xplDlqRHFntoafKh
szRpfdKyQYco6AV1oN7+wJKhBv8ltK2NQA1cfYhvBNJplw3xffVHMM/3GKyd6Lul/OExdzpN4987
P54OUA4n8Cdu61HAdzirRWbP9B1wTLd/mE4vtqRPlSQgfm3IDmOEByC6krqh7ZyLrodPzC7uPNH7
sUfkgbM2hCVeMWNOC0WKesu//ut73YEbZJT3QX66uMbDTPqFXt8fOJAmCvNg8TveyrKBPblBXkfO
xz4XDWZ3GSdqakmL7pagwv8y8ddYIn9neWqT2Wgb6BeoWIfu+uu6FFd5lgmvhHzehOsNjiTii0Te
k0BBvxloxWNSCWB+drBDVndiIWOweR6JrWlE80nqcNZnKuGuczpzNyiF7Q7gxfnnfWnTUCgI2vkE
MBW7Tk1HGZ3ba2R6mCYB6Ns7hmlDNXZsyY+MZZx/SwqXivsMyj7+QSHlnTP7ptugEOUHwLN4ykiD
fqtqEGC+qn8dtjjuLmA10Fi+WpXIgcxbnwKx0jXMxdIF1HywQ0WtV7GtG0Q4yznVUILYAmcoRohn
6nTYpdVnH+qBsoCnyBt385Wv9i06a4hYW2/0/3+Y9hsUybd59a+ND6dUVKrFS3chNIhoxVENCNv0
Oj1YZOwgmZR6EmcmEPZcJB/Qgij5KPsUBttiTe5w7wbHPEitYt4sSN0CIxtFsvhHnaqTQQCMnSDM
yQ6/Evao23zdKDRNj5uLwBJmBASaQk/EGd15a+3NmygCGJUwdNWu7LDgpt2UYI5jHH3XEcHTC68m
kQzmuRocsN7i5RPl3uP74dZFFnj1D91N379XvFFw0MURQhSd3NmQkN2x0mBJ1nHnrh7zGl2YqMD/
MGIpLW29pEQMTNtsBz6Pa1q+AdPfQsWJZ2UANyfjhM2S+NHkL8Qy59fnh4tzbcvA6YKMMSAf0y28
fjK3GFxfmhR1ayHol0q9qG0kUVttnoMGdFdpcKLN+GIEkUtz0ZkQ/dzgR3zrHswv2vR/v2Pvg2Op
KdtGrFcMmL898hhKtSljyn54qY/rLPjc1uSBTtidyMi9kbAY0ZfTp6HmSNLalhxUsHeK0SPwIbCW
5RaLJjhE1kALZ69LU279AM2sHJ1k1yndaNVC1w8YB95kBh3/S3g76xwf18QMe4vXqAN7UajT+OCw
ZioC7WrXcFfHKSlmSYXV0db6vUN7D7qu9Qew3VmdCDLCg7dy1BU+N/kjd5qVvvcDol/By7Fo2LYM
SAsPNOk9Wtg+FwxEFfPky5eeiDzZFmI0oxZkKiXtVrzAaUbyxYINnLecpYn7isRNuy2Kn/aDEv82
BfrbaxmdZMUr8d+iIcjSyzkh/CSfGX+lr7+FdZo35UreMp/mxy1skA257FBmeQAY76ALA1NWfL4c
pNUMQfU3FeTyQF+YweVr4sN/fS11C6QYrrFpada8BlDhEtkBr6S63yLblYZliiV1i0YX+br28kJy
+Vgz02+joioGFrAFOti5pTulW7H1NSTWTsCIdCljhz9s/AUFuwAudKtQ1WyleQuec7GZuoQA1Hng
NTrggs0QC568YO2PdOOtUSG4GTq30DEpC9lkO4QjpHqXvuQIGg9agmpW7HIG8JPu8Exds3dqmODP
yHmSkAqR4J5aV5YSE28FOhspec/UPsy1aUNjVHMIkeIv4e4gmTBnHon4mtIpIh57c2jmTptMKE4C
mHHXb4whzFNLw2288wSzq00h1Jk/KqsBrywcqRmfSxaGFk/rhvwT/pPp+A0uDuWhc98tE3gVVMmd
Ct0nzBJgVmOzhvZVy+C1ZyBBRz1ARcZnqAvFRK+r+pAS5SSXTYmA6ffTubJ/feiSSAGCapYFSNDX
tXxTeHMSpZsuHlY7zQFeBU7tT4RJYYZAQCl/UJRswS9XVggwhwQMeGUYdj6QnSB0oFqOnHdLYQ9p
XyYpPumuxVFv0toaJKSAr0cYkvmvDcfOWpB4JusJ7MXhLgaQaGNRggkNoKIqtw/JZrANoWcLWtUh
6EQaOLCxK5LN4lNv22mMQ9T5jV/nnEOjgekyAzllyij4dcNZtHSdDVMFGyiZZPcOvNpeyGPeNh/d
xGLlUxaLU6yVGxmjMXa03poANRbPU2C9H2ktT7uutMMjTtJZ1j0XnbxeDOx/yBh8lq7aRioZo2bs
XWpqC4AQhwKi6s+/iZlwJdDzBN1fsTq229x0WzDFgktLt3zhOegNL2n2jquPst1h3bSmnUmOGrnc
mVwwO24c9lRP7aNiQi7C15uOrjcCY7JRCEJYJ3lKKAtrCV/M0Vt7rC3DL87EBmMInHMnWeeG3+26
jde+pPq8w5zCvh/H1G7MdpOeD6LPp+Mlea+ampsYxpMyv5PIrpBgYWtvnxmkjESfSQSEJ/LTqe8g
adaWdnfSQDCN5iRlZ13qTmau+sxXBY3ZbR7mYPae4pvKGMqfVDomjA4I8ISjvygpMLY4AN+RZprD
h3qoYAlJ0bcyIKZaD9v/4QOPv4Xk0SmDFnBYJwRqTdDIazEl69adSoLk7aoor471Cax5oMIFvC0z
I58g9x/AAYGJufFHWdzpRoDHEDxZH3VJPPil39wYKFYvLqDvjXMXJkqW7rt7SoJRa7/KwXv3q4tU
+1vzrij0TYUIy2V30BTC53eopHeJj4zMDOYoauPbQk6i/pk61DXEH0pfk9L7UhhWvpVnznUDiI1Z
jQcUwWGf1ERc9cd6S0Cr/qDzUyWtu12XrYKYuwR3a8Jqq243cumTeMlQep/iorkOrUoxj0Cad8zi
iOwRZ2hzv3hpdie0WoZ1F+r+xEP6Clw2myHMGYttojOcwnIlt+VJdv9ASPHvWSrWQiDHn8DEA+xX
W0OkK9rRQY+r6jwGZs8t8EswxqE6T38rqgufgTnKYycLtcUxtortMmOXQ4p3ZM1z2vd5zbTaZTPu
TuoNWlI5au9ctj7gQnvQsgkTCCSEM5PlBW+eekVwsFvwnI9OKpiQPEKWvhQnguhuLrepT/3trwGm
M4odqi9TQU5f3BB7v08RPSw8FOn6sOrlj4pM7nwqygJit0Y2wcOPl20z3NpBdZ55HTMpCiftyjZR
PyvXZIXy8koTWwGomIAQGUeMjnurahkalqPEdHp4wYX8mVcIANMav87P5kWFNyEtZM/GMWD8tKXe
5ju0C69Zy2KEyG4wW02WXNsbEUP0Ce3EOrNRqX9UzCtF6+H+ulypS4BTYxceNBNy5nROcxLC8ANR
uPSiuuNLZQlz5642Ct3WAY9jUv55z24AdKhKmHEewkh3XdN3DhLryY/ELTPmwEENJvxDTFAYPY1B
QUNrabl0rx9BUaddP1/+OajxS5FCwDIFF03TF+FdH3caVhfAEGRgUKqrtB/h72knMn3yqUAgRtMB
Ql4Cyrp7Xk8z+SJt+O79d1waHC9jK5keubJ/ZtauFefaZcEnjZx6SQcSykY0Mx7/ybrMTPgazjsV
ksY7m5puWfSvKkdgV5kxqsRU2JLQM6x/uxWl/SGJJlSWmu3K0ALPaVPyMjkqgjxRjcjr+RgAQdl7
+gRRgrs/SjHjzk7veKULbk1JeJII/SLc/G0SBG4FzKbCXYrCp/TR4+W0ZsNpJ7lDFkLpb8f5+MTz
scJtiGal2vEyo4Ux8EArwbYdg7pHCtjcjzXBV8UiZ/dn6eCqYBpHwLb602RwKmO7Ps/XUvQ3GGvC
kYTPXZiQMDd+BIJTRdBvXwRdMAQZ4C3hWSPM2NBMG0LS7wDNsy1mhcsrOiBn5qPAieJIbN+9vSOJ
Ge2CG86417KsoFDbwfPrIbB5IT5m62Zrxp+haVlCGQKF5zP2+3Wy+TWQwXTYiuh0i/Xg0BPN5iu6
9K+q9zNRISpfiQEyRKljqFnhQ00E1yNJDYMSWPvaiqQGLHQx6s17zGhRIVbTtnM1yIrrQuyPLJXe
/uBgJqhfuR+jLYvwEkWfpxRnYUcoZCEfdz6mbL7ae7UAuPap7jZ7F4LLlY7g6I+95tk6bDtPJwRb
XTUB8lvUb06SvzZLF1Qf54G8fFUHiSBKf6DAv0Xw/u/qnJzXaV7scKDJLmiKU7IVOEoEXNHoKZry
QsqHbqsQ6wXRso5nD0bBt+CBc4P6sn9X22yK+wcVrq5q9KbmcXlk/EfRr0tG3DsScNr4guaQLC7j
/BdUmGW9U3hT72YE6YvM0Ri9JpXM/B/ATsrufcewNCeU+Uiaal2zbjuSECZpHvb31TA32zef3Ci3
gfNDB8wWAwe0hwO2TRKi9cOh0kqFaeX3ZlCA2rR+fF8gGXWhEIxYTl8/i9SWZpESpQnfXUygFMnJ
Ibs4H9OvV6uzigszY9R+E5TaejMFmeX3qNbIdw8AfAJIYWplUL7g/NTbYgA1hZO06srXxFRrXTaO
qEggJ31Z1o/gMCbt41CLaFLXcWRz36nEgn/m1yn+Q7QPCJDn7+KfjTgw1/7LF+JCe/oTiRJVK1eP
cwCVIwyqMHrGISUwF4/8vZFeINdv2q+c9p0fqvAR3uJCIALRRx90j7H1ocotFotssWWQFFT0rTsj
6MQgdyLNHDBCA12khRva+QsHIPG+eIGPumZ0o5Ylgo3+R6qUVj2RA75l4WUb91G07x2zzGQe9QuU
Ozj2tPYWzYarMqtxXCoZCiHKOv8haNVcgTXcrXvF71pcbeWeQxwS9MD+Txe+pm19Vp/XkUHtfjnc
xEI0BSnJekiQEGmJnkDV/DQH1FKoa2RHt13WzvCQk2sej2mh/S/H8d6w3mWzElsuGECxsjGtZ05H
rcdp+jYNAaNJ50yMtu+TLbBwXeHmkLYS6OCZBgjGzNpMsdezA4rV4MTKprMx0QlCPSdOs+nlH0OJ
RZVUzZV3P6YYpMj7gsiUXq92WLbet22D5x6mI6OiL0o1jcoIydTK4v0jAd4cSIZQ3S6LNi9TbuRj
ZmIKDsbI28xGIWS7j3MfX1IVyrwpYcmzmx/QbSENcwMiwQSIa+ZTafpl+z4MJkxLXMammAHQbGc6
g46HCpJhDbE49AqLBLeIiAFYQPeiHtc1QaZp20FeQn1iioEQ0hQxNqPeBBpoK906ta93EIOON9pi
NDBnOJ4WVpbdSLnyRDbeTxG2+i8Tw9DYFF/XeYA8moUwz2QO8RkudZtkAQZtlIQE3twJhDZ/LGvy
PU4kOstZxSUKL9e4Sn1CNs41NmlHMT96sXO9kHhJLS9RjFS5UTGbuwskRuI/0lvEoFeSgwmgbetS
M1QNECLqODytZeU+UaNlUQRQnI/jkHNzUjrqq4aqlH523XTfD9MS+xRfjgFhTBlrEz8l735fShKv
TkyJ2PHohpr4JqCCxH8U0itExG+CtvReIooe9fD0OznroqU4TVZBUolvKFqDx7frIEA9RlJfcXin
nynRM3t9VRhcXGAJ0QIh9UHCoZmYSGxL/7KNWpo2KCirJWJ3ROrG4Gil3QuXYGBnCZdq2JnuvWMD
0ql9eKRs9R1QDDqQjtT1SiIBDT9bFjKFJaRrqVpcgDri7P6MKqpjzeZY+JSn4aSMvapAWIYUX9xI
x3hnH8egvgTjbfjmEgcI70bnL7djhp18q2Pj4kgFOVDYb7HZDnMda9LK9B6BMoxCWlelGKzOqII/
yeusjsvZ7WN34Qik7icxgbIvdwfUXeg6JmsYGzXB2wW2FFHJxAsLXxhCa0FDf1Jd0UMxT4def/ML
sF3v5jbTQdCe25QQlBJeVWlUVvVNA5+/mkX/im4uXpYNwV1NX5WJeR/kwqfbwGTEfVXJzdGSAoRO
qy1MWYK0FvCkf3IQWhTa4QEaG1/wWKvea7EDyjsyydLassCN9RxYhxYksM8wKnxp01wE4eG+CdYi
aeGPC7jvdFhkq+0BeN1vJEo/aNJjfDaoUWYvmLzjwNyHNdlnMy1bDAlYdK9+ZkzsiHAth6anpm37
qkQBQBCQx1oz/Ppkdbi+SfI+u/9nm3W7Mh3mWJSLFMJw+4mO3LpVh19YjJIos9+2mDNGj1sfRPm4
czLIEDm3t3VTrhhLEord0iMCUU/txE0yHjbXnkaD7kJJp/E7koVec9zKiytt0HGFBsLVHYdLitzS
TOs/qX7rOjT1hmviDlOLmb2ZrV2u9xPM8zVPR6uBhYAygV9ohhXw6HWAm5BANbKzgWL60uaEbUx9
LQ39g8gxOXPOaunxkFfDwtco5xqOeKartgwWM+qAnes95wtxn66iCFe1xbZ8gyRAtHJzfIeLgzUQ
MIoDe19X+9ydYfStdA2D0NYZs7ShlgHfYYsq2jnx0Za79XHDtvbQkQVvY+4n3sRSivz1l/1fkCGH
OKg7GvqeawI+nMaaa7gk2hNh4eOVBSVVFOQhlIx0Aret4ehx+k+jau14gkO4MMZFlrfSxExNMNTw
DFZ2VAZdfID4gLmaq1aqFxo1QAPxuFtIN/jjR/ZNCwAt+0Y5p7d1U669YzKUbBY4wJwtuHGxKYC0
0EnCFdFFYGEtp1a0cuBmeSxk7eOSY/xC6vnFwiFRXo5ffk2Zmki79NMB5tcWUsMLxTWJxSrJvokF
xt3DNYLVZOzz0tnHz3yBo2mtuQYGGAC12gnC9l/sIWm2KSByZfsr4AIXKcWAk3G3CqGULTUhhRL6
mfdvqtfMn0ahE/AeRFnNT8jt+D19rJMIt8HrjpPJwKQVCbVjKTmDNxCX66lNbt6PxF6h7ythZEWa
rHFPiGGhe0V1IDNNKr7h0LOjtzQ93LCC2FQy+cFAneMpmBuZApx1eqM7VRq5CwQgnzAtvOF76207
FQlmS05UQ2XoWBW1Ml3WJt7HUjnXFnd1g9/nQqs3BCe+wuO5WERtJEmrn0Ju5w5eaN9ptQZknhYu
TJpCNIOp+/gaaxIgnmF2ACYz0rVCK5O5kTugj8zpjlj6UyU9x9eirgUkTkmjFv31h0w9cliJoBoO
xT7GGjDTc4wV3WmgSNZfnTeTHo5gmJhR3pa0HEtNdFNrKSA/iFy4yLgTvrDwU7N4EgW3aEfQ2iC3
+2dWVc6MpFFUET/GsYEftmoWBfjUDHS9DJ3ymVH4zGfRWiH6GMglxBGZs5Ico8yuVZHZwkdxHziC
8JsGFqdATto1ko845zKnVzthLPnaHNr9jYF4geukzZ+n7evfEZXnQTYdsG/qcn3dq0Qq3XjTxVql
rCXQ53NJw2jn8tMY+L87ff6v4/jJ8QmDfOI+kT1QIUF055llzPAZwC0w8cMedQldoRcuMY54qiVk
/EWaN5rM5ydNtbyodmPquh3btGpHBtdpO+8egNMrqzKuY153x0q1UtIUe8f5nrc7jTOgt+8lfv2L
LOJtukFHW54o2sxRS5YbHZg66RwpO3EJanUZFH6L5OBQ6IhM8mUG3Z1sw3s1oiXTB6KRxQ7Ccb16
qrtrjYs/YF/PSvCtWsUmTqW6NjMevDqP9E15sxXBQUcAu/df2WYky3App+d7NXc8weVxjIzyYiUL
gD1R0iBiWvWrjHczTZy+OyEZDEO7h5LXHsR5sKs0JSofkcppPSuilicpwkzuXS7rgFlbd9+gTmq1
hsnZ6urd5E5xu8qPsaRdl5li85hjLrXsqGx1PaSBvwIUnXunI1pv76gr6TzfXn5NsF7w6pegexTt
J78JwHeNhA8OafrykhvY1iXAKQZr8GbKy8eGhDZtE79P6yIDmg/JnaTkT8lLh2c9S4Nik3MdnhHA
zbWRK4TTFcrRAXH9kUY7x55CICNxnhyANffkSrNXXRlg7lMo6BkU60SaKPwUElRR7V21798Yn1JH
p4XB21LslRaRqWVwThXXZQZUqP4FdDmYoeFhCt/7Vt7Tsb+0nUUfN8FCrDudJcB3KtaGcaj89zg0
N8xanSihe07G0WmUiaaqPCMkSCCHerRlgnD18AhJVuMepnl9w8jlODyOLINi8Onh7HU+ErRtETBU
ShSpXQSh5iIwn7DhixrqoNBO3M9y4BBTUko1CIAgbHKl/tMQEuCG1TdZcSMbEZOnEer5JpG2qbzF
z03MXWJTjcNvqEqRZ5JOZHTuqskrfPJyBvIIgn/3F7/oH2XtlZtx0usSJgtPS7wTdlenNkiNpRj2
qJ33WqmHuI/3CbWDbINzA+h7foEXN1V1rvcjfTcAUhAMLS2Vg8Q1ffc7lpr9ktByePC49KSgR+TT
yOOb3uUtNCUzwT9PFD+lavTdE9SwfMcyGUTZxDT1mSCggG5Ch1Z9ePXZ0VQM82SRlmbNfgPdntIK
HgxQ6Q6ATnUo+u+IqbszBYh78Y1NaLs9ogmUX/+vFELWmvDJUIuF2xWMIAUCL9TgIdq51QxaHA5x
Cn+VqBaOOzGetnY1EUdZge80/h6hOHNaEVd6hi7gi1vGlDgElWh9DxVapIlpQ+RbE+ht1ic877uF
W1mbg/y6e1vS50GmsiwFnH9y3xaLJEQBy4C973lFNwVXmQ2XCti6AcVyMjsMsEcgyFX5scmP0uIK
5fykB9UPqw9L5LDdeEJb8sVnKs/RB4PeIpzplsx5onRKyqTe3PKbiV/vkyPXngIXCgE5Mkp67EDJ
2MzJO+AKAA9y7vSCa0Y16K08gZFSYgSnwxWgya5FmjxlOdXWoI+XL0zxFdnHZtp9XBV/m1whkNfz
brralirYgLNEp9qDYTJCQDSykCkz22REsbmmSKmlsVfqUfvK/xRI9cdW3NzP9NHWIAbFiddA7BpV
F7bVU4Tf6swVxH46f6b5fuz6r+6rvR4Tqj5V58MxVf49uFU6PtIO0Dxnd+mtzss38wewy/rCpuux
TEOv+QdG+SjuPfFUTqg4VIwFmBWpa8k5sWkuSkz680Oj/VKnb80oKdY71flzBzZ90zHm3n8gV3dU
BjUQE0MMXdeGqIh25hVNLMpk5/lllTU+cFqGw1BiMjTFR8px4dNumjY+8eYJyxgyUbN7I7+1ugGm
uIAMYWw5vbKMdZr1smqA8bRP/kBCKy0WdJ/K0FoLaNFlARWvFe/Fut/BAMXqRjLpC7JYN26Ff/iS
Fyqw5k9L6eLG4cj6a5Y10y1xJbLXqA456VDuV8W6iPjTJSkTQOrEuA0r7pUlXKn6OsYbrjuTzUuo
NX2q25Pkxx/pPAUlUTe1Ehx5qrbEmDS+Io6CuBoTARnzNi1I6vNZfhN+uYsAee4xwS6KpIsGvsYI
muhsK2O6hbKc1nMEc6BA4OxmcKfHC51cFJvzSEHojAeW51+rZ0L9Nd9LqhspF95+7KTkiHXNWetJ
Ln5vetRGsEG/U8agXUsMYJ3rWEqQPLoiF+DxC8VNFQsOzcYvT6rg/dlDkaq8gVpxJFzvPSpVstgp
54B2h+y8Ehex67Kqwx9INDzlXc71f/yhGGHGMqZg+Ob3ZtDIsZmsyjVWO/fsY4elYuzS9cahlK23
Pqb4qxYmAypwEh/3iQLNmLv1AoHeF0UImJOQNqn07uvDVyqDgphshyfHb7ZgcnMNfmGTpGf7OFvl
+HXGH+JI3GfDDVvyyQ/WygZx75SxmHL0zVq7tyl2hovynj5SlQq9GOy2JRaCkp9XPzI/gYv8k5gp
VkRWs9K4XzM81NgyFf1ylrWp8LVIiggsPsUdC/pEZ4V6vRxP0FV2FFF6F0OsdizSAJnE0hlJ9fRR
YvqgcJy7IrJI8wm/YxpHLAoebagIwl2LgPixjg5GsKLrbHFdTrlB7BrHTHR+NXwENQgBDDLtYdr1
x17m6M+cablfvvEA3gIw56QFJ1GeqI+g6gptpbPwC1PML8kIRy4tgzUk/WHf6cg8cpZp737UBk/O
dGB7iHWyaP8yoiQPkyklxuQK3O8HZoovxggRNd9qhK+AkJn8424VHOvXoifE4tF3zq/LLdT/9TdQ
sgL4xHMziNIN56KXnLZSsZszgykT92mESb/oN/SKBW1T5Bv2TxzPqBbCknQilfpVST8vfRzB5w0r
8N7hjVo5LJ4SeIFyEAoKrBt5KA15HNI8rF+qIBxvNzXZRgK4TxY9UT38Qz0Xn+baBHo1Ls9AmotM
/48ILA+yrxDEn8cQVWCwA1e7WeIMjACM540kA4VCcmBMq1xf4wtatO7JeTClksIyJnG/mdBZWqaQ
4xQU67K9Xb0VIWvnHd7cg+LTorPLAaAtBDo09/nv//FLR0MQ1HfXW2s1dOp/7EGUcVhD62NAqZXU
JXtUS5xy3UL1tBw7bAa3AZ9ed/LD6V5SZcWz7TNKqsAK4iA2izytZ/nNOxEwJSz1vG68h7uJsYUr
GH68jJ4dJLTyuj/utjSM4xlKVj1AwcU9zSRThGzXziCggfqLt+VNayVBOX2BrE7fkStWGDBMve/5
sj0HkfIhEfDsirkTjhypBg4Hrd4rZ+ZW4ggeSpPV3qkMDWblTE2sPEFCVMUqtUJYhKxZFoKiVeez
xjbqIUYuqIqGvQKDup0AouQERW1vIEm32uHiLWCNcdDUx3yYGor+7slNT8mVJvlWVw2skSeTG4bJ
Ep6KCFW44Ud6biPbb7XYuQE8caPseiieNwIP7iu0fWteB8GWUNy8hAzV3BR3aagQsFXuAnxpdED0
IZ3+nYGBCB6oKZLMtLxTlsehCNwCzwVWhyKMI4olajSEYYuFDzuyjnNoyHHpzy3leeYP3F7I6Hvp
RKQ/9Ea+wSriYKIBn2mWBq70UGBPuI3F0KOQPrrGtF/x6pg2eNQx9VVWZQb39eOb3LpAV27AKCZh
d1m9GHgXKES7guk6SFsuQcGIU7lnk3M/GGKGjwTaRhxm3mEmkg2r5Ohmd16hJjBqOlGD0W0dNiSx
XHAq67bGCvzLCoxiaXsQMKmSgtJEkamVe7fM/TeNqgMrvqyTE9EhWhbdblvSPOziH9HspvLsepyz
zzGuX+ao+1TlfniDJA6/CLPI7D4gAbZDiTZB06+jYakcZrht66Vm1l/G7g0gG3bYszgbnzjy173m
k26Ob5IUvXHJ4aWYgWeQ8ch/kL2ES8zPI12X81M7r6XJbuteo/racgjeUUbyl/wVTX3yh3IEUnfP
PshYR1vYWPE5ex/6/vOEyPgrBJUjvhuyH4sw18tvnLBaVjG39plOeskI2BHfDDIplVhMTWw23TaO
ljeDlTpGT3Dm9TE+T94tdVSaDkOtxaskgbnqfLCY2sEK2PY3ox2SnDHcthii/rEUdRtffltUcMNm
es2HFzEzBuY+eTs0HYOcAQ//wiTdwc5xLHfqX+I0MFVs+7QNqhKigYoai3dDkdv0bEIrdQhyQzHu
wtIQGb/K5/DGReOIi68oeHMvkBtg2v0ecS7yyhUjKfUJk6W0VSefsbb2KJURugbEkxcwDYxgNAJT
lT636Hkl1othYUvFhLj2bWE5MuHcmNGC9lLxosiBJ5hlbxsA0wvOboiOrOqKT4NiCDbQMRBA8mnN
OQ0RY9Oq87RD5rDsZPbCD//p/ws6tsLwcvU8jazL4dXVwS3/vNravg2+7f1cMSm4gCodeLi27rON
gRyTYH7QlKRgN4vLL8gJPg3gRXjZ3D5GM6YrNJIqxMuJS90wSJZ6zZum8rPR7HryBjkhz11giaTw
MQy/TfjdtwJ2lA6vcVW08cnQ5fZsffkBx8X9snd0GCaGbs9GRwG1piQ1kGI5RLKt4V9lVHBIAKKs
mu0NH0ze7ZUKTOp+nT55IDoFkWfQPfP4RdJpEaZETxU2Q6LZU2szagVm6KevQ70YnRS2cAwXtDeC
xz1Y4gsULn8Oh5CmylKvifnOyDp+H3ifvpcVUQaY1KjWxnivmyqcLfJE8kjDytncyuY4Kruh4yqY
C4p1U6K9ebSCfhCpLdvmnXodkoDxek5r7zGweCQwBKImsSAujsgNJzVPq5XIbWZZHK3PXCh1jvdP
2KSHd3hAj+8E2Gc2J92EKnVD71/ELdgpeHJ6UV66WItVppcOO//E4Cil3E26cgnd1Nv2XWYYibVQ
59eKpSYSpYwUblrWA0WTuj5Nyr74SSJxHbeDPlpquB3TbaYbA4p1DtrxQKfpbGU+/5HSYqkzysWQ
+dGDLKNRM66Cr1G71CqnnYVEwAWAUoEbYntqYdGtXHnVJPcZ5TiGlIJHqFAAi+dgfgdb6nxxzxcg
T15DAIA6nFFjj8bNKNiSQorxXPgP7SNPG63X4KUoS2vVC+ULg0qbTCa+K19ddWoa652od2Q21bLH
HCdi+s+5vV3Sxtmj/iPxNtg71yFrENYJmNjLhqd3hG0m8vkDPDPL6NDOltZe46JaIS4knKVh5EyT
4HpdY6aWmQ+k3yAoJ8FfUVMgb48fgiOFSqxYaIyD8M7tzzhCSBZ0KaiTkCRTGAwSdxinKZYwwtRW
cuydXLqs5dhUVXe+OSEYbElzn+R1woUckOTcFuuHpPebBsIvLvMTGXhr5p/7qNMHcxzPNUCFHeyZ
jaWSQt95QSm70rjjk3R84lq/3QNbQAPD80KAwOGNiWLeRMeEGxBIOy/8o0+vOeYdXk9fLVw/ssBX
6TXukvt6chkLvhPVGtcvkYBgr18qIgSjmQtKT5rdDyMrKfJsLKWvcnc+z/uVYH/JHFcDT0co5AwX
h1/1C4MABj9CeKbLn4lPRI/ksxmg4x4qar2GtqKmjUpl91NV7+dD1dyIajwa4skMYSq2UntEr2P4
5ODjcXFH7q0yVWhEYV3DzGEu4tyAR+1+ZqKTXpGrcW4sZUhqpdqSN3Opb4r/XwNotW1cz6YWa0bx
hdyVgmEyES/IrVk0b6MNREOMDJypdg5XuHo4Ni32sBNoXq8VuRwwyWmPJIVmaWUlRcYZed69xbBP
fINw8aaWmk45sNPc7eD+Kp7hMGtc57GuCOTkhpLB0gT7EEwtv7KyowMGKGtyjQRjivg42+mwXyNV
Od7iglJHdSzgCEbuyJ/Bc9qmI2vqa8EVxDguSYdlO0gNC2TMPskae+ic6oa+Vfp/uceE3LOpU55c
rHFdHIe37bREr3qX9YhTwnToL6H4KRQFdhuBil45xtrZH2nMrh7FgOyWmcN0LP/QCpBRb99nNOp/
3ufEHCARM9mY+BgMi9cr23Gxrlv5lkVX9Hv/anVBOMYOVv7PmvZYYfhQj8xISNdcgV2cTPR9MJ3g
OI0Y81taovJH6to7iDvjUDm5BH9hxWO5yrC9Pb8UyHJ16d/U/HYSSrLWVimTyG1PL/LS6zfnf2qH
oRLokVNVWfzhkZKJsYnjPF2y4ly9dqbCQThv2Jh1UgQ8N3BTpOlo2qd+x2CvUJghnF5XqXZHJjz1
LFMKFqv+aYpyJf9QjdcalYezvWXoefsVeBfZHZKMkCcE6llL4mKnTOwob+UnN6I6fBiYmCvEAxYM
32svYQckm2ozuGhIHdO9Y9Yb7WgN8E/SX+3ATU4YjePTTZhhhed/RCIwkwVDinkgaR/0GJmdxVIf
bXFsefOr8v9LNGWauQNzDwVpLcRK31z8gTX1XQ0GLksfq/VUgCjjwxeDV7AMYaeCFeo74jy9m5CO
5/R7v456nngdSyJIB1EcUMc0jqstC38fS6U0/woq6oltG4z5xMASj3+pgZcjwDQn9rN2DOKCPmXk
Tkn/w+arK+ppKWNiyY/KU9n9enoGr+oIFaM6/x1q+Ex116RhS60LbI62xbdn3W7vuO/CTHaF9e+u
58HP28mTaEdWdQwdrCKMJXp8xiSAScYlgI1xB/Ue/h2rnB3ojvV9qzVBy3PcZdlR2hvccw+vx4NV
Qwlra5EdtPeaLoTJQMIQdXj6yr579XempgL1/whmj3hX9pU2k0jcZeFsr+qpJ+LQ5tce9jIwIbFn
MFqMusgv5MXkXBnOLogICsKDvzf4N9YtA/aoyXHCLfOqs1VpIUB6lniCjqG/+bo9/aUUGIjP6t04
sxdp3nZMaI4B4Vk7iB1WBLaFjuOApWOsfgIFq39Osotb3svtXxKeNPC1bo46wCrAUnOdaDeM2Zw2
feLx3p5QwQFnpZs3tysZk8iYuwIm0v3tNVUVCcRB7vSSC9rMxbtyBPv2xVdeq4XUnR0Ucj9CczpS
7XqCPi2b7dpqNcFS4ienyvLTuJT5Jl469lPhdTcx751kk1uHF926/uuJnID74OtSA6zADulL0L3W
3qQXEiKo2t9wlFVxCi7nVAy64j5E3LEcj5i/E6rt9sVl8RsCFI+u8Lm5C00oJnq+ZgA2rhnJKVLk
6Eq15c9kKoPMdb5QzWrnCJE9+uXrCKWINJ/ATAcYo+DQNefv5osnZ9ONXPIt4jBX7abbx1sVtVqz
BSQmZHKyaLpCayATV2EV49H9c4CcAbQahmct7iBekISbarel9HUghNyl7VERs2q3NoADb2bf55xs
b2lY+GKfxHO8DjMNhtrD0ZVdEVQkih/GaOYHgtOBYywX/1KSOEvGtfIx810rjmiJox/qMuXgJx6q
Mb3C6ZEfuh6Z98UwKiSXrjaMma25+ZLYHXcwhI9Ulc4BdBHDpQaq3QdQcYdfzwvUuqSb3j5Wvimw
z6KhKwthUrdif5QSe9af5BsI9p/M68T+jnsAItrba0cOyoaRi6vprJfQPsjfvVwYkVGclkLMUtuy
Nkh0AMflZ65bMlbB7ZOY6sRbSQ+MyFobO++4CPH5bigZi+p/nRjdV2r6V05XDyjoTnvigHh4d0pu
bvUwC16g5rRW+zm69UlCnlMTVD7jk9O2oYXseM/wZ5KpdzP/fSClhDZj0QutRhfefTdWZjlupR1j
t9zDxaidqAB+9MqptPjif5IjWvktFCCOyBi4wdqCrlFAWfNCLKC+Ka9zLf3y8p+3PqcOcYcVSdL+
rv4IOqEtzFLrkTR2DsPbZyRLNbx1IRamrnuqOlLWQIjvh90HaoK0hhwe8dIpoaz2SU5Q4ev9O71M
T6BDlnqUGS0nRqVgfdn4079ofZWi6sb4kQ7j/Uk39ZAFBB1wMI2lElZtteDYeB+fhIoSvpviVccO
48qw61PKj0bchXX0MsCT/75vxiwWhEORc0LgyNEJRN6fHDAglRvib1HLplboeWV0LUYcuH8LaQX1
rdjajHMUehDy1vW2I9VKtY17VUlNBhsbHMdz+SdobzovPJFqcyfBXTCYTEGUFI+YuQTH7Z2XFlWW
7beAVjLWkmFNB2Z/ovSv6hocMpTO5y5ptcatH7QuNRyYv2EQuDpeJhNCWS/+KgKXtQ826Op4nvAS
nCV9Xqg98DV40tz7sDJg6hO+IoFyBrdbZXm4ZslVt/kNCZzr1VxUpwUR+/U3UKNz8JpYmH6x6qAn
o4MvZYvC1wf0QrdAJkgyQSn6gKB64OsjwxrVbGxs3DwlIwJJ0p+u/IhGXXWtylCpnDu9+FREYDya
a5ZJZKRpINkXEhgQXZLicuHSZSflqPkzRrSthJoTiafLWdoVe4mEeNT36AkB/QuT52b89h6NJmso
0BXDNrQ3UT/GPpTMOVfnwvILkMc/tFsz9BF5Oo0EwRFYocg760xFoS0lZ+BDDVXej/pMZsRONXFe
dGlyRqjzxPZSPoATz3rLlNgTMXzXKZIoJnDm3C17/zXuvGQvN3jAtyiQCYUWSFoIQMHef82nAYnb
vL9ynBR7UbfZbvJ89ZyF7L0Fm7UPunpJWcODIhGbs2oDJJWL6xcPhijBRrIcr+qUzc0QcaX9krL/
E7AsrPPm2CZhedqX210bgRAyDrAZkLwNADJ4Wn5WmP9MZ2wsf9YDZLhnsnrZP9laX3q2AFlb/iI0
MFv8ke/KoaDJbUmOcVfsBSUsJXE4lpFm0AUS3Lqa/wMvFPkGNaO/GST4zyNz3PF0ug5JUWpBfxW9
a08hl+igme4PO95N1ehGbMfM2lmrpXrc5MdFBZ8anlmnEjnUhiLjl3S1+HzvcVY6kXlRE7VtrAb1
ULCk0h6JnAgtecWd1aU6qlJTlHxNm6Wn0DzFOReRoxNyUj9/TXZNuLusbp75fZGak3T4s3B2qE+4
Iv9qbOl3Spc1NjkaHwenNtUwdmuUZYvmXgq+h8VrSd45BDF7vnUs7JzNTe/o1gtUUWyY3yrmlKJu
DPWPUrEWtw5wOjBPLhDm22tn0axi8GRe79bNk3+J3r6E+jmB1PZmhEzfElu6SKdc2cU5szKpI7et
Yf5/8g0qlr0QWprikzKPIoc9rZtyz+MMuofukqnYW7TdRbxZWbXBro50NMRDrXQiqVwUMStSUwrL
7gHW3yMnJ7PAMxXeX6/Tgnxsn9vpS6C08co+1ep9ipj9OIqsfoialTVpSPwFIzj2wedsNNkMHtNq
ZOVsECbjzYrUyxg6Di8o91P9fdUHdWeaV/jbuve0Gqs7BLCdIhHsoWhgbrcddb99VkgUxJ3FnDkd
Jcn+tlogZmO0STuZyWfx1XcO1yGuW3fBzeOzRTHHkixRK/z6tB6IyftLfv1jaXDMyc23MZMX7pXp
+6MRkyXdxXquT//K2u98p7A2fxfkArYy5GksBRfKsnfVMoEsjyDBNnZKWgUJzZv1T4xLiq0MstKR
48R5iisiN4DQU5V/zLiWMIY3ioK3Fm+JE/u/P74aZNJxyTl47HPbDk7e547MkeVk+PJqXnC2MbV6
1g82ldNJlSayrx/l2keKb6vVQuBeItNOtfrRiZGTkDNDEsGjj1zOUUQfYonfbcdcPh/nR24xmuDv
m82mW5x/bEALhFj6Wqj3/bCiGushPyaK7XmNsk9rn6xh0tS2BbRylAEHo1Fg/9i3/0faaDE3f96g
dz28x1hyR9ckPCvMFAdTFHN2eLUh3ZMsg8/CNVrv3QURPV1DVA2SBtvtwvubYTPrzk0DbdRwjRTZ
upUZlV1HHUaUCef2civCnrvuoxIrVEIS6YP/ocHCQquB6azhJOC3WvSX5s/I20ekMI70bWLrRzZj
tDXTC0fnmPHdxkyTlrmtTQQGRkPRoqyFPx1DY/556I9DwpO80x+FwhDWbmFonnW8hOPaxTiib229
lPrBGnACx30vG2D6ltq366m31tsLhx+FiyuJA8tmspJaWhaWP9Y6Nt76trY3QFjVLMSMrwPcdnNv
7sWaAwTMg4qDHf1esIIjlBHHcE+BXRBrSNobJ+NTwy9Vp/1bJ0gY2vVvqhS8VfjIacOXfSfPeKTl
Hsjo1bvvk3wgvMaeVy8KMPpEXTP3VUDarnksp/qMZzWswvpU1PG/j8MupiW0ynWv/RiFxQmyTuDW
NFAQMY1PGUwvt74FcIpqfh37ftprKHGBJrnVBCSIm2aMeMi9oCrqB98cGe65GaWrFp8MM4Q5OaSP
r8jH9o74Lwark+2e8E7xbZuuvF56PXnyGLrPdL5912aQimP1g5JplR3LQm3ZrKUqmUrbENof39YK
HcKYKffEdGM4rfY1kMW1IwgWmML4aqtarRkdhHGakzvIYWJoVaTXihJfTiMGX3alE9XdhIyn4mii
SIFMmZ3DTcDp5MevysGrCmChxD5abkdpVFQ497+fVcb3Iq7HgJJTozwVrZZs2T6lpwP+KsN8UuPs
RgvgVCwKCCzbBlKKYW8hEvOC8ZuSQ8TLwcJEqvT+yuo3yQhoHUkx3LLXQMPleK3csewPtT+NS19b
Zg4enEGon50ANzPFuYPTF6clj27RK7+Ln2pj0D4o+ZAmuie6arf5cHVSXlCNAj2y7AxamTJftD0V
VMvbwRsVEStHazXkP4LMvR696aAb3GA9Vmsc8/zP19DXNo91pPJUHngPftAM3uN3Irbs4iTbOtxc
rskr+QjdWLHdG0iEAgMi9D6x9a95Lt0csyLGcXYFs13CPaq79c0K771yaFA9gf9sqsA1UayrZSQM
Z3DtYecVKTMVcbj0J1Z2DpoxYeIKds+3Urmd5FuV3kYUs5JmXs8gsECgKiWMdA0LMWuJicf3OhDk
jUVWKDB4fiHrw0oeEHzPFegGT7EhwlOOfd60pkNtIW2GnjfE08eG7RItG4fPCsnhPe8fvXYC32tl
YayiJYfwsdvpTHwQgeD0sH3715dv1+Y3t/Jm7YA/9IDGUrWyu+FgbCcIihUucKgv+ZwkNW42afu9
i2haX0ccZXyZ0/11K1WwARvSskmwrCT05asBxqebyseJt/1SLZmC2wO+qYziE03ZgINX/GrFBiPd
LWg1x+okWygJ3HMblEQ3occqGm3ZNktHKRrjdWksCP8D8iI5ZEapIuTZfTWOKf9LhHYOIpsE/Mav
DGkCFelsRVGQnK+Y6KlW2oTgYkqqFXOGv2KpPzJT7Qb2KPkolE/J9fY4KBC3jRBlC0eH9ixa5YmR
jKahQzlRs1yZocXqp9UksPPh96aPdMPFXSJ3ZB0/5kv6cmnInSgScdBSVfqIqitoLWn4/o+8S7+p
VgKNmTGPWj5ni7gv8+oZ4CKlQTKSwLFcr4HgemEiAbnhoCjVWGs/hClk9TFf7R1v9LNB0Usj449C
KeGMkxKTLXWor0qQILzDptOzrdyiRPPrjQqLzTg49hYLlgjWjTSAKy8BWeSSZmr8NzQ0OZJmRvw7
jMnE1Ju9GiB+1OxKGzgZ4zqvQVx3u/ekJacut0I5tB3XK3+Dov00TtU1w0v/lK/0zqy5JdAGCEwK
KexqXw9JKVrkz31gdzkF63DqCc8J6ks2KL58XeiKw3LR/rkLUUDWDA++GbvWqrd3QzzoCfrwRxoJ
Z3m/U2EivFaPfHZ6adAfH/VQbdw0YQwt3NEiUm5lDH0BiZ2t2PmLxVMyzPeThsE7Pr5oF5MiO1ys
skUDR5Hzgd7op1sbRUOMLU+gzFBrMecBZPlFVJCtKx9kTXytVb6IiirFPpVxJ3J+rT6iFWNEdhNi
JqS7Do0dy2cH/GVxrFmxPfq7hvNQRAasBH0YeEZGhRCnfYRqZOl6enOescgGmBp2UQb+QzXijwOs
G73mkLyhO3JgRMUcVVDwtyVdhK4TsP8nkuQ9KA7/s+2hhe/7b+xxmdcz0Bj0eQwWy+fM/+TX+cwr
0nG/04D7cFpYrbJnHcROHC7bJW2+5xY1BHOBm4gm7t5rQv5QOz/8niiwi3JRTOY1HQYLByvGsXQK
VGlTr3/eq7yJjQ21VKZyXX4MRp3bDNs1ekAh57nyvtEp28051b5/kxPbh40oQApohfez72UZZO9A
WTMC168h0ICUn4wDbapP8h1SSOCXs22zPp9fEsiBt1czrBVo7ahmpF80DDAyeRsu8uGnAfewcnqk
qyvIqnEHNNs3xwm//j+CHdWNuld+olwa++OFu+gl37hYQQsqHAGckaxf7MLnQx2vZCYuleBH6sUl
U7kyf0h5FRc9QDUhgO4Ke0JcjGyPHRNgDpKlYDUdkzqTac26Fjg0L01PCwYXjNxZpJqT867qE4ra
VSn/lPm4eRgAKZ2rwQQQNjmJmLRYZ5tQUO/UrlVeew7iTmR7hY7AR/gXiyzcYsMGCqt7gWo27MgJ
xM20ahtbgXhARYqyhkGEv8YipHLRM0HY3TkW/J0AlUbwK3yAFja6PHcKniwIJRKP8zHfm6cIHYih
AaQyk2L0V5rYkTatnLFnCXKYbUSeRqCrNpSOgSI8setljjDDfp0dGTgoogudXLFiJAHx+/7miy/u
q0FFq/BF7Zk/BpXNAFkJEWwpqWizU5pZhasnJQC0yF1DFNqwNbL61W3W5ac4wE8O1racSvNT7RQa
W1sXd2Lef++HBiW6LUv7XogGMUMoNWSzHpmkj/et1ZH1vCZWRbV9OMso4BOMkX8oD3MxCRhSwVtS
jyCNVI2lDMD3z2coP7Ew2orPssm3GhpVBZUubj9wp01ndldzGW+nmhAH2ouvnX3/FXTBG10XTL58
RDkldnVi8w+CMv+r+SX30kD4hYXji5JS2VsGl+0/CBs3cnx5OU5LLLVKL8xpFeljHrdl+MJH+IXG
oj/6y69s61ntjGv/1+U5zrk4kKrf4EVBSvTAQM2QOsHH/ntPUca4zZstxipRv6F8JLk5kpZie5iq
fi6chIjGTd0dws5wYpiD6b5Rmxybfs4ZJGsedMqJzs9St2zHFUizG9L8ZsXZ8Vuqn18wbLvLxoSh
6iU6Xc6SKnR92euyv1/gXT3TyO6DxWjJ7VDcJZjVk7/U3V78CD9wZ4w4uD3T7v+Zc+Ms+TnH4F1F
bADtDf8Od1eur2B8V2DAP486Ec7gzxqd+cqfNPqeBqArJfHDzcstZ0g4XMQj58LZf4sWYEkMlIBo
TdGYpQuZATmYSnCmHJ0yU+zn1uE37ocCMbNt1tetjLy/jGFMC9oiv99mB3g+9w+S0IsqFO9lWsff
ZZKNz1lEhDN8ByuCJlnRmevbKSSLFoBeUnglITIKePbccs32DTxm+ttQdRxeWWGlMhNuiLYKYw+L
PzAj/RxKK0YjjP5kXfzSU8dU3qQFH+kuX+/K2n2fkSC03+/e6Oiz961qT8j/pXRnBoKErn1VOHph
8LAPlgUxKx7H1o1uuF5YrTcoVyGYfMN/fwsfsiI2nRHJIevWUrDls9H4vXRATbTceHYrAZEiKyNy
J0WauD7svH7JJu5NM4GtXPxzKd2YAmstLTReWgPYmbkQ/yKhQB2kJmD7NHHRWofiULeF/nKZ/UuD
fe/0PrduiU9kdH+QZnaIG2l15cQafPwbo7iH6i7h/CPIzd4B1qriez9y4wto6mqM61jv3tSmn+vO
0N8ObhPCp5D4Qaw2Ibw0YKG5TQZWBoaYDbr9K4WBFIKakj/s9TA5df7i3rwwRbBwOUmOTWUH22OP
qeBWxjw4hvwkYKXqh2y7Zy+jVkqgkTuOAV5RDhwTVLW1kDub+5qX/ymnzQDmZa1gBnaAJi7tQaCi
9q4Ge/yTbJQ8doaShIYrwBu9aVM64wE2fB+SvU/uhXSh5TD80d7HSUeTtKiN5+m9X9IUg39PQGje
gNhDUW8sjXNe1f/HMG+MH4VgFV60LlenrPBz/wFM1X40NDL1rl3O0tMFXlyRtR8tWh0IFTi4PiOX
VO43OpjKjqkgO9ui6mhQqEQ6/1mv7rSlHmW1l4Lm17KLJRCJHa9S7Aq1W8r/ZFs98w2DO8kjbu5I
dAtWJvcYE2jO7/+6DQyGeeE0Ln3hFeA6gTg0V5+4WNNsmXqp7NixkkNsPTZ2fcg8XiYSEW/6cTlY
Wf4ZN6s9jjA/MEJunlSFGhqv3tpMVDyACtHYj83O9wMCg0aE91mfGUn++qCzCgiFSOM5gpdsOYwV
FNWwDitIhygU/nF46XlNeA1dp+WF/Qllvd+9ZRlQcz7ZeQNXCr3ltgZyR2IloCMjUlT3eOXu7cMK
3Bp1logsxbAvFma5chlwog/njLuy3bgfpBQNJidUkfjCykHZDy0ZlLpb6Rjl5CEXOzMyWdyqCJRq
OX5WdCbBuS3l7C2NRKkXcGjDJDfTnAUgMvt69NO9MEkCRgJrPIr8kkuRx3cS9apfkURoYPlWbDd7
+7R9Oc/6W6Nd6Z3tdQ7wt44eIfPRJWIQ6sgn82lLTbTqwRhs55G8TqNBufx5JvNv+AhLm1XZeD6W
qrN7PVHUmcJoCXtgUdG+oQXTZUYITrU9AneRjvHQnr3xVuStexcxh2cE/10cnNX1TdXrqXbypntk
AXA6X4HdFVyfNWKh5whA8WIhBteEznb742pQcvS8TmWM35YeHkh3K+ZG+832QN4LbnwXOzbhk4RZ
HWKBJqZ9MIomS7vaG7B4TEtKifTpYuSp8ESzqmlQz63AjqdE+qcJpg7/cqYTZL2meJHIg2ZYM9Aj
2q0Ug7FT4EPlagiv+cXZfFT2+6MfbmhygK63a62A/aqiwjh/pkwWr4312CoHgcqIp9n50jjh9bD4
cnMPQWiB6aP+7incq0aNooDjYTcc7SYTti9Sd77Y97lwIc7VBPnAN3UJbGFapE2U85dig1ep4ohX
Vv5uabp21ep4tP2+PoPuXqXrQK6LqKpZZWdkHvPRfk04v5p/r/FRxnyYRh4c9wYxHTo7EfVQK+nP
so9GJbLNSa4N3bT9r79r1F1+vkQAJiVSV61R009ivrYIYCIjBF1520fQflEMP9Q0hibv9RakFlw2
1q7ehcG5kd2RMhRiAkMhmELGDKeAC0Eoht5un+0J1y8gD0/xckzM4Vk2sDjQsOql2LFSBAg3XezN
76/2VplZS4T1B92YpfbJOERxukqCxnTCVJget0HczUi2QtfosdUfm5JdldSZNDFRlLERxS9qSldO
XJEuvfM6GTUaJTrgQshqZZCmfJ50vo0EXB/BF3RtI0rzn4uDF7X68atzMh9lT6nfFtFGwxLpGtcX
F7+FypolrG3E8yh42SbPidOVr+Bpldsjzf9kWd1ULGOAc3U7dBJ2uOv2DhcJjdeN1nGyq2pOwCQL
74G6smdiOhkmbl8YVHwD1cpDd5zdYKZl2PLmS+HuWl37A9Ldh9GVe1ph1ySMpLdmgUfg3KnZv85q
DC45WcGc9NtQQRUsTDC7K4kTNMFaAVPXXyAaVGKe6PyAoxa2vuipwWUhuoVkIlg45uD1fLkCntRM
28Bl24sxaYEMB5Wr2NEhD11F9eGIAJI6HL3KVfELjkxn1qSfRhyUDlTO3jCQfP7BZ2XbHT9MzsSk
XEmjdrkdgxTpGr+keILCSqiZj37jf9rgPIvrstvCoQWLrASi4Wyb6sOU12KjTdwidKGksBL+qPUp
Le3RTUyCRcvoiksX0ChFJLWsXEs6o8PsL7MQhZmfgymD7adZh+CH2Z8/LkOSZsQeEf0GvQw3QrOR
Bt4TVGP5e6CIAP9X4zqLW/Uys8Zal5ifouAQzj70W04jSkTa7D2UcOJzCeqXjorVU/60vnODselh
HOA2ygVj/hr0e2GcG3sGqp8v7JcV4Euu9wIWUDK/cKnpeSNRPKs+N0Io0sf7IT8K7eHMw9gkqU06
P6ubvlKqrePZtfL9yUYfwjg//Z9q+WkGbuyMY3LJsf3Ou2Sh6nFOvclOnonD41YNX+aHUun2gIjJ
mNZFLE9O8hKLoxrnX6FUpSg8okY26IT24vc7DWWMqSdpl5InC4/dOO7VuY5BPixvzmau7Duoc1jh
EjQbmmIRZofZTOpt2Op917KRAWJqRnr2cqHUCyGd9UajzLJnGkx3qCiz5iNsmhmgEADJ6/zsIOh/
BMtneYgtxUKEUBaGVXdsYHlN4ho99ozYajh3XzLVPMmVECR0UTCLV1sgV57TswqJmQJTn1wsAKUO
mKCoQciyEeEi5aWJX4NbKxY2KMi8q3WXLzS50J5K43pQSjAuoHcFBx5YjHyv47mPWgdNEtxj/Qvg
3JrZuLOaWzcOZnckxoWBdolekYRBCFrxU5skuGBI4VQ5jC9gxTjknKGjkddEWKOeFeoOldfuCjhC
NxGmqQumo+yRc+ojRhbzzGPMH7Z5f2vN3S2I2ivLJIrgu0bU6doZE5LcQubbWykIWiW8W/jnM6Fp
hDmLYWfqemqeePdR3EXt+SExEaKturyk3zI5JBzmuXemlKr67OeLVkWcg2rRY96uLdUP+n4Tb4Dg
QaVk0n9StUaLPb8e2o+m2c63m2arqDhkxhpvtqx293S2oZZ6ak8YkNGOKT69RQTeFXddV1hr0JiX
sTtDytBr7oCqd4BRCPxpOjZFQvu5+HUpnvC+UbD+oNqgx6+21vpuJg2z9PY6el2e3Mm9FJzIJVkx
QvC3WliJtwdjdz21JswInovPd1ERuYvzh9oWHhum2BZKPaoMTcNlpkKazqVDM9/ESZzzNjQLdCdH
eo0QdSijM/E+c3nLiOoSLPzW5+5ojLlm6lwadD0TDE9ddC3TIZ8YYIkW3jpcmxCBy2Lahfyq/M1D
tZ4MEyX0hKDcoDzjG7fFd3rMJD9yuv2FK7XoQdrwhxglhlLAif5o1XoXa+0fgI1b+m3BXc3UGcgc
p1zNDPY91tHn5lXRrNYNJClA54DLmDs44aXvurdwNINRnJ/2rGsAJobuLwnxrVTd5pGq7D9ODTeJ
phrVKeuc73AcxPPvtDFbwu56MCrgmG/k0ReqViyic3Sn4ys07v1ndX4gXp5cp72wp/XWy4p/apbZ
H2h8q60ADr5BCclHFdkWpShT2r1ubwBdjcV0fwVT/2aWCV0IHvH/D9C86HUxeS4CEFeRX8pW2IA7
tQNz4H4tPkV7d5k6oG8+aPmNPLzID1K9HxcbesbtlcbbGB4Xka3XGY2NOqG0PmSLV0eu7alZT5oQ
EzsSKLjA51Y8TDICU2UPjadyrIF/WEEv8j2ToAsNcNOPsNqCgnrbQ5owS/LmaTpdOM7m3+FRFstz
jCwYeO+o7gRHE1g4sWunX1/FJ0WIPs/bxbQWb7fyOnQBAJ3xuqjh9N5Bqwko4XqBAzfyOCWj7Kwd
H93Jq13ZVd2jjnTyFzzcg1CtJKN0j5s3HGRVc7IDWd+Sdg01+AiEx7kXaa49b05V1xEC8SlwZqdL
oXTBUzOvIuABs5Ljf1Rr8IQG57AwF+bQkND+A/WaGOizbkDh+LYQwbMLDoyZyOpzqixBVtbOPQR3
X01Vg0PQDnEwVh+zd8J4L4NaKfHvRoUn2E/0InH966xLSpFVmwQoyrkKkwFvC6qYJtV4krYcVrv1
2O4b9eLJRYMz/JrpQKwG7pWeL0dubK8tBcwulXyAVscGoGQzJMUklJUTWY2dEdaA7BT6ui4KTSMi
uW4uNc2MlsVZmPIBE+2MilA6fQjS1oj1fNOzGmzgBp3msNREsM8pSGwC9nAFDGYq7fB4Q/yey+cI
qywnSnrD4PTmhLCS4g4hv6sjMcvrYzcObmSUV0VnVGUpDLwWar9Na2C+lwHY8aS4spudhfmETqGK
cOiFbsYOkvMMuqETABiEc680/fu0zxwkc3eNTNhC1wY3UV5ErD0/X6L06EIz++6K8F+2Lqw9CTo8
aU8oCzop/XWwiLn2lqKDGzwBTT/HW/rQqfqrO4fuJwn8Q6x3XR7BOqedV6Y/K+PfkAbUf+pWFEJ5
lXaHHd/R2vhuDyJud595Vxe5qs1Xufo/XoqGlOFhn/k/Ne0UJiP8Mv1itV7UktQHIZxcjgkFjEkL
7gW8WD/masF/q09fwX1Cvtm6inv4Y1qb7q4E+ctApeJ05ubPMcyZ9R1twAloewPrcMEuJFqz1iJf
mjPhuneuzNtdfuFlFfZetawEK6/yy+75DXMvXIHi5AoKgoL+lN2vreRZJ+v+jo5Y5ZVa8lStjvWS
JR6pA6AD5cDWQrZ0dTL0kP3IjyDQc4ieKtS2oKwbyUeOIiG1KTOPWfUtEUZpJp/b9nlmXS4w8BIY
8iOzLoL80BPQMlab7nkJeqgeAJbfRaQe+BfGPpY1HYF6f3ykRQ7yTqjGNBnlhnUASQ0YlTlQvfRK
AGln8JVNRFDOTjiFm82oAeR7BZFUnnd8y6zQCtqpDFRie2bbxDCLKmLXy+IgjsKiWolwDVGrInGE
szeKR7WuSci8scxKsEkhTqE+qJgNLAiGTBOAO1FJjz1koD3aPXmcwluS2PEVV7BmXfGdr/qXcncH
g3n7YWIZseFR02oiEllxIp7rmPxswvQzIgTJUDcH30bj8bBt4m0BGoIeXP70NZfeJ9sXnYqKvpSF
QpusCb9e+t4DXmDPkQzbglVbLvy+z9AzubJ9/3xDLv90oHSXFV4++83pPNSFiEKJonzzq/KN70eY
Qs/p/HjAZdOIi+sleJUkHgrcBZAtUjFRI3nk8ZF6cBb9de+CTJSp8ttv1DeM6ZEGSbzEN3ldn0DM
MRTHB7m79scb+IIGo3fSRoxc5l7pJyUauqHu+cQM/csTij7N5ZksjZDAZGGKoV+PoNwx1nKb9q23
xZVM82sPU2kaoGrQc70OCg3V9jlLyr1ozCxeeoWU4et9UqtP5OCAXTfhB1046eHFEMX9SWm5+Xt6
EjbacD0P0d+xOwx4a2o2D9D4Y0r6hVInyERdl8CNeUkM8ntBSB5Ldwga+fPa7Sr37cuU+MW95xGA
8siQ/sz7MM+LkZqpExe6sALeXndDn4RIMsUUuYnbMb4JiOJpRe2TReHdbb1a5AT04EHcEW/5JELq
n95F2ytpJzrDW0kJUhvQsy3z8W2GFrTF/70MveEpFRvOif2H57Z6g9CM8WDgd294Bz3hHhq71NT2
cKaIZEOsHOY9KaFxESazlQyBQnKZL1nLqL/b6L6VWnH9c0X/ZxaGRdH8GtYHXPsLfbwwH9/bCLyn
sOYg75DV1zIs89n4Z4oge9KiwCptaVDRdyOzcPYPplu2ydR+XFYKUmPpKzeGabOLVc4OX/v6jP64
w8bIPVGWl1q+1mUx3ILoFVb3TJnWxnOxxWohSbdn0uSh2dVjQkYWRYeLgvtjsN020KJsXznrFqbR
rFsrJwcU31wxtGe4T2yhVCqAlpUjt+3c+GwijfCMhbZna/t8tgYXoHsAqFtN9bZJ4NmZ0suCt+0X
oLCHozn4lkMOJT7PExta7i8LjmilFYf4/qOZnPmjMFLj5vPsSIAX/6I+E3O19XP56Y0KVajDUIPa
Yxd7pz24Jl/HgZuqKZlBFX3O1dLUXUOeRQH0i5H7gjHTL8nnD/1D92hd0dgMkJRMwEHKll4PgA0o
P7JKMXnkhVEKdJpix/VE/nufadQHrEIdtBQA9khZAHijgC3BtqQNVHHV+1lOodvswYz/+73+wmAg
IMXL2FpOrr3NFKy94Smar9rsR/hCmUct344R1DnWHhZ8BBLDoOO952y2SOiSPic/JyTmnwhX7pbI
Tx5Y+00+f+LaW3dQs5VIYvzM5nb1Q3pHbB/v6LV7SiGMLAV6T9oBMV48nwvZ3+PDB0LKOFNuSSlI
z3axtzpUC2cE/pCmZx0Ou5omGbery6x5hN32nK9BSyCpaTlDP1WDQn8AnIIgTjIiwNdZvAlAYeDi
E6Z0HO+ssvYx9KSyw5ItxDCmeqFcN/CMWloKv5JSf7lSCc3XiikhJC71fbRlCwHE+XXVjFCiB4UL
4KRhpexGGDQ+mtbHgd4K0igCe0nxvQMdAqnnYGaEjEH1/iwdMYKRvpDlStGJwgGiIjUo5TL+Z1T+
SlfW9xCtE+D4HxH7f3p69G3Zb3WgSo/GWn+VeJrPNe7NNG38vIxcKuc2bB7dXMcOMnDtUkXRnewi
tPQOu9PUKiNloZZwUGiV8VD1dDQQIL3Nut6t+ZVMKsvjykg1vd1KUa5QzSbX8WQlx9f8pwepbWIl
ZxpkzR5YYKaGNB52qHM19xPmxqKb6oah/5Q+TuOyhSl/kEEBni/Z+qWuyXoSDdAqQJpWY8cq5kQT
/mFM+DU+LvX0zX3vtf31+/Y2jY1W8UQDp2PN9brfsfoNddXFFtIA/MyyyAejYjaDTXt2o+wqM61L
R0qNwBX2L1aScXu6AomzuCXZ9MutpHhngj//oAiV9kJtIhg3DqYCWlRr72UX/VnWOp6h5P9RPTQn
1PZaZdZfsjE5cEekOaw17bTmGyQOo+oDjhrwbDjEqP6QZz+BZfDqgDa5EFtYrOASqaNkT+OozOsQ
rUndOLXvZrxacIEpci9zMeJlyI2qlFdK08KCV/3VO4SFbheE0gLPB5dsWeJBD2EeMbnySIPGsqBH
WjojXDHp3TB6bsV0FaslaKRwwG+M53CdjJ3t+1ZdhlIpIzpNgWTtmwG25d/lFlliOBeD4HHuZAsN
XG3wWzOnnupRIIsPOfbkJSX6T3anjHsu0r15jMSEYiTbU7C7WsKtzGyoOwW+GfsFi8oHW+OwnSbg
9CsrnctKJPlGF+Qvu9t4QVGbJz6hisN4Dy3P6+/6ltQepy7ubGbdgrj7pgopmaUoD9Py5WNEITcW
jZ6wq6WJ9Zq/rFJgp7hxLh0bdcLiQ8WjGlcA/MD4NsxEwqQl9QBOWwrMaqC5irFs9UtyQ286/pMK
KRz7dZiIhBfFhZLhkjuUmS50yWKbkO1gf9OK326c9eB3MAui6j5Te7owBOX3v5CYafSqyNtf5rjC
5MLtwIydUsvIrZvwzqOaLBzrt4Z3GLBClBbPBmGXP5Cx8pULdc25uKouijPKF70KwNmCbAxzbS4G
7HAWA/gF0zwClfEuIs4VMqTiPlt02O6OpCT1Cz4ULx0Q+7/Z2HAaCScoNcAcHAjDDkn9tXmh+oIE
mml+2S76dO3St0c2XXosJRNPb6AdfJVd3SwWBuNrY5ylALljK0438YqkIf7xdPA05PRtJxne2kvM
x+WR0b22WZN1N8+NxQ5eegH+YD91judtrKaO8sor0eEdZfta4TBTdRBdIWjibRivsExoyvbGG54h
tlRDZ+bDe4T3AXtpiWxZACmmIbvcetZ5WYYHF1vvgAcboOvtHCyCcrU8q0rY3kCz4k3Wsd5FuP93
un2tl+i55QeT9T9PiVV/DO3IQhNj9Opy6xz8ZesYiWgaHI7yOV1/O86uDDAuM5qab8RggFCc5IpY
Hszc8FgmhyvTvLDexzHNik/3gvTLHMBTM2dnMdFR4mHqiyOLhITSc3oUuf4la967eT1gmjeL0YGU
fM0uDjSCvgVLZx5c31/CIqJeglY+y9oHKJq2drwysKVtsAW9WLJyUvllmhxpPOXpMRYkb3jiuMDg
g0VtkbuFxoNEXjGHtmGvJoDhgAV33Lr01OdMUc2CG7jvMNGdYfnAoTU187Jq/LYvooAMRoqAntfH
lIAr0RJNbFquYh/QkKhTMtC3Q8zr1TlsiRGCZXX9zEITDzSFY7x3LkZNfXtMU3VxYdZ8bweRIKNq
7FdSmm1+z96ntu0sipjW2nezGavmmjMVyLXrwWNkJkH4y8qGt/Jyk2NAdcJI3s9THh8ehiZKH3lb
WLFs8En2O8lqF22gWez/Q0Ovb6c0jeXfzPCMZJM3qwo1PJV3UGuFlmQ+c+FbFXXybu9OVG01LeDM
gWjD8NpHKEMBcaY7wLYfNLJf9aXwGLKsPwlWDptTQjgav1+HbZtEmcPJceTP7p+wCkiiTtsYK23m
KVBIw9O3iwkttEaUiv2TN3MBMQL1LPsDhpSLXWYHc2oyJypuPKS1SnxSav5EPk50cMNe+fj/fd+y
thOhLSyUB1BHtMXXGuxslUMGGr/w1MZHly2+WinqE7bxKJ73qllWoHh3nOwFia4uwh8cxAEMevEX
Pq/+Pk8gm+u2ikAOv/zD3P1otOxIwTFocMVuIs+ccUl1AbkJXjkecNwDwXYtJMiZa8q9MLoJXZgL
Ex7RtzyAOt5ssql30eBUBsIcFtEhXbR0/Z4vG30CO1fFi0xvTxi/awjwqgVTCuqjTV1mzD451bgv
44BNYeOnUmNxhBul5w6R+rUS3HjSD8SU7XfHAC7Jkhy/srMlFPBXv6PcazFAIAXq3Tw/JTsyyGDf
8let8XSGLH45TPdNFALPPGeL+Teqh0zygE+Of2JsGZDqsKIOr8qiv+Cv6o7snNs6SVwVkmfjZpQg
btIvl71+goWUFZqsgtoWxcCQTGjlOKHnM+O/bKj9gE/drk6kKJZLVm10hTSm6mafpkM6/t2vgQgO
c7C3xrpSt79sUOg1Y3kUP4N7mdAXE4hHKzp790XluTbjOoxMDUbQbgpZckOc2AqJkLP4kHSrZi/O
d6XhUBE/zqz4OiXhqh3biTR4F9uf5/WtR94oi0aOXsq/f0Up817QXWAxB4WPPjmyK+5MLcaP2yY3
9mfa8USnuKUqrZxHv/d6ITjbvqqn35GLSAosOnJJ/yAmf1klWnDApAyOU5Fb0nzA+Ig/2AHyDx20
LwvWx0cOHBJrSb9LBapLBiv+Flk+wOGkIzCSMkA3tmha7DTI4W+p5ebfEoZ3+BIkG6E1hn7GkvKp
TznmMHJiYeaZ3ASGvE9Q8nQFLdCishFo+bOQm0BWS/B36fmeJ0Qjvq2SqitVf5vZErsisdAPUwtO
toBpVg7iMO94YqjH+ulQqJCqLvuqYOOROWUIthcPFtnNtOrYoolQ7q3V/p3JUZOPciEM1gCHLy/x
HrCO5M4c9MQ5gfPtJa93N/6z64YlCpJRDVQSKmRD+lyh7Hvy/T9c/9/xNbTZ7cInRRqg3cyaQX9p
7h+ADMop9C0nXzuDMQqXRgfUJskdhuYOnqq+R+YrpyEPY28HKDQosnRaKbclpEyeLrxWZtIbDksk
tlIm1TzBwW/WBEEf1rOjyhcOrKwNMClYH/fYpdv1zkAtRDyjGDzdy2BQtgafNT8Qgh7RkqEI+q12
ekuD8D3nGlxgOIbC1nf6DaTX9qU2FV14XN71j8TMa5r6IG0/HKNcVBX3bMUuyQi21Uhq/WPwyLrI
J3dSQ1AHL24yQ2ZADEG3PcYDTyNGBrKcSt38B/lboQT919A4tCWfriMdSJWB0ePHSPeCN+Vf6i8k
3xM4BoCPxLlm9It2ZpwXgbBqmoGL4obg4izU7FjpXKiX8LK2Ao1lcW+00/l7Kzg2gQpXmoyPFgZt
cJqF+BfU280EzBXI5avjtztw/55sgB0QOII1NoYR2m3rnDC7LGmZwlS8/oEA+koR/Jmg/9SQFuTm
DPrteMKWSxd88z/w8rXw2e853klWwyXZ0NuBguOMceBdws5i+hFtyLbbg5QZAVqygwjyRpoJaK51
G4ioC/otJDFvh+LI1LnKF+MXEQTf8/TxzSZzOKxrPxW+n/Zc1nUM92Aoeftv1lY2kY9h5DJNoW6X
JNTJ7Sc5A/hIe4evkjew0odI98+b5bNxRWdvAQFo1bexZrbt21tJ5+zNeD49ZZju8kcryBklpA2N
z+xm6MW4fvph1hdaCwc0U9YvhU5eQZvyhg0UJLzypebJa5V1zPR68JsJy2AsBWo6nSsK0+hvBrOh
wvtEyuGdwro6DFHxjPRlwHsM78a7zor+G11rolh3f+YAa2+BPLRUcbY2Kt5tfKqxZ8xGetGN0Le2
cbQn3nDbUBIEUOG0SCvE1O13MOQKwV1W0wHrmklDl53aHB6UK+CdgDJWMTX+rkTlTNZWSBhV3JR+
S+M/KMOjXmvjPbYgV9PEcJO8KWGLFGgUCyGHu3ENKZoBYf8Irbn9ze3S0V/JWd3877JfKNBB/IFN
4KYWzgpFIkFK+SQ+hPLL/vtsDNwHSGybHmwJqQ9dJGEDGMChYq0gcjENSjQwpoOnq2UCtWfaPLph
0YlCChcYImXpsnX+SiVugzdvLd2QhL3fTOLD0A68REz93y+mBFpboaoyYYLnpYyD1yd1nnobJbfU
ybrD4wbWpCzi3w2ZRH6ONOoC8iexDqRw8BLliYzvWhgYi/DTaKaWdnoQE5p6/Opcm8PryN2coJz5
QhjeMWX1cqsEqX99AAIKGrRfV32BufMoWa9PtLtK9mjTGw+qlJpXroXrvoylAB9g7Mx5+0puW56n
SDS0rletL486Vx5mX3aICJZPWk1dnQ3lPe84WKp+Kz0CfR/kiYC6mb59nV6Zfmn8HoFP5Fxj13wS
ZYvNZ4sgcsXb/DCbOxmgxew56yfxePR2S5HhR+x8ACp2VYar/LK+QDug7+4CjiR1JMkSow65PXNi
1ObNkmvfbI2gIf+3J0RWt3zlUe4DRwIzmRREiXVCsVioFdlUVjBsoMtW9xu23qkZloqOA9YvPSEZ
vAPadbIkQ9buCLwgzDe8COykaPo8dN1O99O/YmZ/Afi/3FKEZSm7UJt65Gkw81D9bLvClWJ7Izjq
fWbCW27NHwn7VzVJgfSz8pNkJ4beU1iJMswCB4S4llaeM4XpFh6mc03cPDSs9bhkaI84W6oiDBaf
c1cORW94Pn2NsQTpLN4XP7M7aHKBoh653Rdz4kaO6sF1MTwRnPujlpz/jd81gdeq7Y/aTeGJtvFi
04YAGD3rz08iDuxWGNjY+B+SJUXEdcgPDDFpnAk7KI9Djqfi6VhDuGf7ss1vt7dkEkvMzjv36sfw
9kcYUtzxtpnBJd/tm+U1jPwfjo1MffgIVsG3DSIu7H6toaIQQZukr52/buA0kXjSD+RUbby9FUEO
rIUliVrIlEFKYMxxUecbufVjiwsSaRzyOthZUnFAn/bW9Fb8cJ1Xi6PJsWjAiWmnlz7OUDzfLmmt
Wpt+Njmz/5X/7mBsIOnl9219X70Mj+RgY/P61Bd1w7aAS8HJfgHvKIXi6jfFiSMXZWzbZJ3Xs8bP
qq02a64oF04Ut1H8FcrfT4OpY8yCriLge7aKeraDBs5QONQ1mTQaNxVTjghuk+4Ldc+WPZqLGIMf
jDtXzXWga0sif7gZENkkFnyRsURhOoQ/Mo8fdCSmV+s89APfSFMVaBDALzKXiQ7bkCAt9AE3VV/q
j1KxQ9yqYHSa26jv5Sq/TiPEaaCldC1KBj8Z+lNLpcqWLh8Tg4zvyOs3KOXHpcZQQ/fSazNTBSSI
0Mq+93LMH993WIOlNsfJ9vhMHHV/OjkV7V9bvZuIiMyi4whPnZQzy0ubF+TlwXwHBTMobSgAuiKn
pRYKfFUy0MLmpaqGyXPvHbbAx2FLksSbZiBmYiFQ86XuoxXpqvZMEOQ3espDvNH2QX0Q/C+HvlLi
2CteTMZnl04UL62jodxGk84ubnGtnw+Pl/iiaMMdgfQqVyLplZd6HkYNsz4kx6eF/Oa6Sm9K8mIj
8J5SBB/X+2rtB/IGxiPYXpKozeTTKxaAQ2GN+HHvblCZD1L4R7rr1R5Rh8l73ryekPLsuIKzzVIZ
LMwRWu5nVPNLGdEg/5/ki4UGlGhBQ7tsi3uiTPYzzowYsxsAKqiav7Iu5WyaycscTIst+aaUD7uC
D/eYfpa1m05bochIO1ib7LlOqi3OJENczljcyJU/sVlftvxbH3h4iXQThebSWDzr7Y8AI4HXFvTh
cwyFYi/AePs2yzRwjuwej+3oW/hh7vYmGXvID7Y7UUR8cAr24iIN4znVltrXuSHp9p1v3xA8BS1N
1YC90xwl4jSlOEugeICuwhjnxIWZMyNgAY8hWQqjXqxc89RMS1B7hGlLrga5Zm6asTznA60AuYYC
6eqoCJzYxYoUaMaJvVPgrhY7uVD6Vh9+fSbI1nNGGHuBQPHa4UmhTGpHkxnVPU3FNzifIpOPpqBi
Ugn6ZdMilVQTbqSUruon9XhrdDY8YzSMt7xKvLbmhWQkpXsClXURy8NK+kq5Ps+sIV7FQzHy9X03
dXmy/pC+Oio1QpeFCMYtHcLyKhFS7xvy9n/pNY7B3A39gU8nC2VbS1Dedar/43pwgDQd1jthpD+C
2UPwv65UrHcMQR3smNYbJUw62JUDof5Tc3D/gW7f+6xbqYdoozpkDNlPGhoLzRMBniNWKKKFo8lx
jrDjfNvfdwGSlafCR4Xx6iwYrNY6kECWjA00pd1IXUHLBK+h9yj+XOw2LN8tUj/VHTS6CZM8/Hkx
unwaSGfTFcT1LHONI1jtK/ymVJcyKp9zvK2V/2Z/11F4U5oCkXnAa+VaDytNHVGAtou5wF7QODB/
T6QsJ8PUsUXBOPQCNtU8/Au7FW/6eU4CHcLDXIxnuA8dmHwN5PNTD4j3UCJENehrgHnn20XlPRri
eq9Xh0P43ZH1K7mQ9CHierp5122zoSsKdYJVFrAsGx1cKrA+otPqzjR+uY4+9S86OhRHwYDCzZ4F
V1Bj6ORDWiS/w3j/n5FO3Y51cw4n/rzUzFVaRFo50NP/pX+DGfbPfYpr1L4o4aHEwQZp5fNsx4mJ
xvLgDVzUaaGAuOSM5/SKLHy29zKYqQ5Fr9zaF7hPjbdxRlbIY8tJ0ixDuThNOlbC8nPnyZ9yjbFg
PO1nXQuQZeLC89qLNMiIJRw9Zx+hEIsyoqkr5yJvsJGAObEJrgLB+hh28+2zTMxtRzmttDzqqucl
39HArT2jLG1QWIGThSH/wl58/nHPNtrFstT2KgrV9UG01mvt6mgSIXmO4lAbsitXMhKC7yM+dYEy
saVHqNJNMam7hmev9jW9GSCqFQGymmO/JNe1GX+vAlx/VWuzLU9MbQOafrvVY5TjotLflbnVrWNY
8zmx7HMBlt39jRPAw2CXL9FojKDd9npF2oWnAV1MhChfMC0fqlTsBxQeGC2reSjbQqvXVWdP+E60
yYY1tFWgV0FaW/5Finu1ORZlFIzLbHr/6nkJcc2qpc/cb6VN9lrxOTcN02Mbciatsz5UiqKsHns3
s8Ajh99pq2P9PwL5VhHR+/TrhHE1yrW4eHKBGzF3lgCr3QenOWT/v9sNWHPa6TJWgd+ZkYj+WFHe
9VqnRgK0ynVGt8cKcC0VSXV0LNVCXHNK/esdVqyeRTpzoqaL9f9XVoRiWEcqw39wWu8ZVHM2jHdl
c/lA0oJevqOV3BJzMQ89svfE2T3oIzaZsRgPDgtmT3pl5a+SKCrzrC0iQRyMwqzgYAyTgI+xa0eT
i365RjjI583PjCJahA+xo4V4g29q+zcEZWFxpyo4Z5udV8xaEVmDj583x8c9v6tmjOJsdkh12reV
DbgU13cedPa1ISUsBvgNr8YtdhK2pcpCcs5mmfTdzyRCJWuuzUq0OskpKqv4hez/kgIUYHD1p1ib
RtXgdforzr6LYsH9rHxaZufQtK3HR/xlay03fxascutjWcwXo7pCCvuZJ6z0cMgIFt/SuwtkpTRX
2ASA/1ih4Dc1NvBLlKzqL0b/Ti2uhQ5jplg2KhdcW5IG2bfmBZjXJo9J2cKtOo61DqsJ/+bZDo5s
EjtCv3UHNeYwqY3L4oRrWMziECCHBtwKZ9ZQtxrJfFKb5nkiFyvTP8T4eNJ0ii69h3/vcs9p0/oz
MkLM5+yJkeA4y/P6ZxvO2Bdf+MvDrxkyFEZ/eNjy3NICGE4nD9eZfQFNwYb/J1rWnr6v4kpVtkKg
Hwt1Zd62EykqTTtPjAEyZFpBKz1+rKpuKR5DSWijx3AdmHMkI27jIe5BYUXFOpv/ZLMMEZLs5j73
HmeZ/s7RMWJ+LDALkli52WZtqknPn25YJ2pf9DNQ7gL6yHlDOupiu5ViAGkyTU+wJSYBBuwpq+9G
RDJx7T2FqW/bjx2067C4cc9NHCaaAFB4yAwgOZT+XJ8IAGnnGaP8q3voH+5YP+0D85mL/wuftHjW
0c/A8EI388KA4PGH+8MPw6xlv4Yx5GFlbcNpOe1O4ySqKw1kDpmMldBEHo16yEanqb3UkAo/8xED
UTt47qxuLAsZtSnbDokyDKlNm+04fRt5CwlKAxmZAT+2wA3jJPdM3+SKs10KNpdR7mPu2GaNYI81
Epsxsn3YXqoMXNHB1sMny0gMWaZV3Y7Deqdsw51cUrsYxUlgomChlWrFkARkOFxP/Ha5Lk+E3Duv
KTQbAJLvNv0iX5KrPrc6GPg1s+u2apYc2cnfcL3RYblywP98BTETco/ISuiOEffDR8F5L0sZyqP6
uDZPLu2kC6hGWFw5T2/syrsiwANCZ7lTsxeiNeFLaaMd7QQ9Wnmkf9hmvcaeGjeUwrIXfbaYi+qY
r23eepxk5wGRiSGVeZPYFrrcKAKwrOcq3/iDZ26ldieg9QySXo9+palEEtAdeuQUZTPun3RsoOQo
udgsYWS17dXQZd2b8qLEXEr9TwiUKJWhh/G98hcOVwYgTn1yzQ8Z+7Bf7fG3aRBxpiNtv+tgQ9NZ
uIUJCwdRI9IXES7/YHWUHV+4ll8nzLgCQMxMztK/DefUkGqlgDb6tGnVx7A6DXKtKaKabVgaL0lc
biM0pVLpLERZ4z/8Mttdjl+dcIGP+Xz885IQUJmeU1/q7mQfijmZG2uK5YkEVNXC6mRd6PE+ZUQ5
1qt29EV0Mpbkl5rrRPu5mZAe6bUrkDt4b2jy1/xQmDRcPFToAASnvYKKK0sI9DHUPdtGeH5hjIxU
teQvSr3Kwo8j55rjie/V9YE02bH7ZjskmRCToRy7wWg5c/xa+jIZWN1716nq+19+MN7BX9HsVtR1
LAd3v7kNFuyzETI6cFlilamv+dfZr69xpgHFM5bgtqKmI+lj+E/Vsli5l9EL5RFUjXKaG+Z8uX/y
I3A5R1V95+3ZGiMq0gwoLpbYQqPKMBkThoVXYCKBgCbw0HYyXjGjw2f54YUHPCFl8l5lRopH/1Y6
YuRdxHMT4eXLI/3xQfmT0mWW21PabpoFZZAJ4ko9YcFiAeLNHuyCavj4oWx7cDmKpcwTZFbkE+92
CZc3FTEuMe8szTkzXUTR6w1U6XSMERh3GDIxMw5Wjzfl7HkeDaE5HhNLsDglMiXPjOtp2eyFNJVM
a9znyzgOazZtIitKhIjzfY7xtGg6CZt89ziRxusDM4/ZYheGROgZJV5kYlbehtsMsrbLACTyKm95
JxZraINhvHJnAaVgrPCBsFLN2Uyi2zfdWrZna/2YSQ6zr9rHSBbYomL8pc1l9ck4DiZ5AIk4fe4y
xZartI6H6Dk/CLRhg/DtruUxcfegd6jI0gS27stSs6OCcro1kGSLHyODdUlSAIaWrnfVDzPlbxcC
1d8m5WMdLAhcpClUq7nJg1K7VHW+xTctUBCsbDJ11X28hr8EjDGCpXmz9y7TGdAO8lwtfDQlLccx
xhYgRastxi++pXIrG5xQUvz0HegsNS2GgAZXx9gqyvOzPm8t4xS6w4Hn4vrBBuaJQHNM184kvRM2
QIL4hxZUnsfCwhgKZBq39bE+T4t7sRxhXX86VydIr2xDNqPkTBNFDHYOstR1WSTL/gBBYoSXRgSd
k4/ZOh2Zw+XozsS/makyZ8VMfzLqxYbyrkTIItxOuewn0JThOwXMgqYsLzf0UGdMFocWCIZenfDa
RxNye+od9qemVmUfdFuklAYyX3oKzNKToh/EkwgD/zygFMidxYgbeeu2Tuog9LiOukT+EPUtlyhA
4xtDabnhPv5tU0bViSBHaStjUzkZB1VpVhHrSU/Sp7nOcz0u1q2vz9yX06SjNRPnGwEvf+zc2HyE
bsDe22ZiytaPs6LWuaVbwk588heHLUBx0KH2ic2QDlvrCak0JJPTlaJ2VFvOnHWWkR8MV/0V7VDH
MuejjjQURAbRXG7UUYu6BW5FOG1lq6pqgAB33VoqPHMSZdQoYkDhrz87Y7uVICb1AAzb8rZQ5ECR
becp5laIDVEFsN1xX0gnr1hRFTApk/GsQGAH8jRQkdMdiT2WssQ7Fb0Tjymz8ZSDIMHWdD4A99mr
e4EY+OUoNEoP9FB4U541e6WgMKSS3Ej7DhH3/N0Np3XI8LTnLNdV4Ji74yr45FkGJKOuDAng1PsP
a93EsxVSTBmQmMqvvvXwtZgjuvgdF8fD/ppH73QwJK1CfR2m7W/s+26Ty9AOqEpCukL5+3KEfGSD
edXKwsB+j6fCIrxlgJSE/WNd99iVt6xgvpp36w1w4J6HtEp7F/sWT6YmMh6aVcp+WmLbdfOGtytW
cT18aNlGnD72qsW+z12IMweQC885dGURltiVyoDBZkt0aYsACI/SH31QRwmgZ6VN6iOYiEdiEY60
VWf/BxV1pfhx6/2WXMLVMekjBfq+ErDQG5VOgyc1E9twK7494u/4iCZw/TAufB/tiQjdg6QQbtbw
P4KyAPt7eHI7+8NJ4/UBm7EBlp/z4En8nIIZ7ms8p4mkhKD4UQ5t1zDl4pCOWskNKH9tymWWDilH
8hdkfz6gj/sLJpsM9cp0d0iI9ybOV3H7dR3EADYHvVoC+ejujra2fG4Cas8W8/Bmngk4ziIsOnJl
MCc1Bf7NOU+yzijZAfCbbCwNVNn7hu/UPYqVo4fXLtUli92A8UTJuSuBZh1TMqUXX1fP2wktIUry
7QOzSfR54f6p9NQ8eqkAWA+BpzjyQEFsBk/bmxVZoaD6cAkWLNiThud5Dnyvtp6cKQspZr6xGmHm
gpg8iKZPgF4C6UABmMkY1NK7muYCNfGQKYL4EsyO8yiZq7BAm9mh5TcfxfstCwf4YHdfejiaZdqH
YCOV6NK2lGyqDyXETaFqD0GEy22Exv197FD7yM34qwxVXL1VFBtXoRd0sJOFJV1SnJQE5bS2GSoF
nhZO4r5kv1v0l0Ry6Gqyrrwe24Fg4V37N5Z0D0mEF+xbv/xbYl0kv+oINrOZoj2mNYdgkYSGJmm5
3Bkjattc7rzVRjWTl4lKwoG8xMv+DQkUY7eHwIZDaz7dMj34y+q+IHVJ0mfGajiHC4G65o3lVWTt
xbYRK6mYpIRPnBDUFxkAk/FN0fEW5/u2WJjp7YVxiXP7zizZmcL2X1FFZF01Eg73MR+GGCq677Y6
qd8hW+rTUn1wCGc8ciN1D2jtUkAed+0AtHW9/5+cSBfdiiDHSMhBhrpxKXJJmOL+JZXGilPG+Fyu
DVqOW0bJgp4eg8BsrR+gj40qr/r4YfimluNY1Fjz56I5gi37gSfKbSrV6/6gZUGepRt3b1dZJPwP
jkYzRoWKytbNzeqYXxvso9rk3tQGoZYteNy1nsRXO8PB1sjGMnpcc41sCQgZ52A8j3hq5L5Jn3YJ
Kp1YJqmoeXK1+fsMZudne1Wi7+8pJmqA/DsBCvZpRp1laR/dNYGQk6HAexB0suDz9baDRekAHDHv
bXl3+6wc9eGeaCl+B2h1g3sB7+cH/Tl/Q28pU/eLxczE2Sr9WoAqzLdFCUpjohP4erYl1NirC3KM
pMQ2O1kxPDQrJGkQ39e6vDs9vCkXPX0M4XVwF3cygeEdpkkYpUkhjPNtJnGsnUb9TFEBuB9BhTQC
tbDTyTbMUFQaWxgiUTtzsGFgtFPVdMPRMYw0HPGInSBD6maOJYbXY6sNNyzAmM+EkHlmQHtojLQE
AoRgj3qzL57+oOY4UXoDyMThWmiHfzIThidUnUeqchIdnIiBNywoy7tDJ0fdFW07PkOj54YMOXBA
Z0LNhbQa/MmnZeYDR+F7SxfA0+fDPp3rrJVaBFR4s++LbtY/9jauNnap68C7ZH4zyYzDLs5yS2RQ
6a3emFvEjPD/3ap7g6tgF5iX4A5a37Vs1+Y02hz/H+FPfi+vdhicgKLA36L7IlWoJAs2JgrRkAPh
QycO3c2r0/cbhydqNe04apO8WeeUbXCS9aPupX6IaRwIlOVWUxaAM9ZWJDsZxWLnjQ99jGnEt5eb
JFrOOT08w1tgEvjRNjOorOVadN3uSM6J5DQzB+zFz5SEfrccZVPRdiHGTnS/L+GQStI+FCJkCHbv
of73FwbnStc/GxZkJkrUlc3ZSp6VaCuNEZN/GmVmehppD9ZTCR081CXL6y4TrLHP0JLwmnzdc9hH
PwUO7eizazLKhcpsyanhepSie6j4DhSw0soOezMzRUgaBHcKEGLqfwKVCJ9qh5JPYnB8wXKvX26J
49NkM9RBT2WpUWGiw3I08Xk7FsR2NUIdm4Dam4BTK2EABGYcrcr4Phw1JE6NHF46nwM6SIheaSqh
1+ExMdj50Fb+nCmALut8WldFqeLuD9MI2f5TXJ9HtMy/PPMq4tif55am2yLvKrm4NC3iA7dS7upa
nNtc0cRzSoVSaHnn+R6a7OVQPhgk3zRizpBGewQY82SYvyCaiMMhO2rN587lSoYo/ASlvlwTK0uN
lpZkTnDuWv3r0cnCa3u7cI0qQw8Z1dBlSdyRsiMMWYs04tnxV87z7PTGNTP1wzkRbsN2owd0KrTV
GoEpwGwG0ipIbg1IWPQNtd8WBDOe7V/SEreAir+wX92v8G7bYEHPA8ggCi2Io+XQjfhRDTDwLAN3
q4PK04F+7JWihS2Mkn3XGLmTSdYOMA+DfVmVzWJrBs188IwviEucSzZiAk1s9Ew9kdl2Wvkop/xY
mnNgeTXomZyym0lF+KwHZNZ0XZa6M15+O5dnyzOGxe1hcuihFFoGAhX6k225JXpBS/+NgW0AFsw1
K4ypdD06U1IJzjgmP7WUwT2pHf7DCFTtEVrkjfVqhhIXhIlopzUxp7pWayo/ZwjhihsP/4mqjjIU
WU2o4R/oJLQPxtD8lLZynHXX4iArGGQ+EwoohKj0y68YXMbXR/HVTru/sE+CZYFxcjAwXcZyg4Mj
HDvdgMDtpp4jaWSFUMlGUAWXj78L5B5RHzij70DqXLulmxfi+6Ra05IVzvEs7GDkeJkwSqdBBtkq
Z18QHFfZ052pHBgMll6zqeclOY6DGVl9Px5w+OBqdg3BhSCGQ1TTgwV2PtoRryX3Qn9Y+VMh+wBi
RuWreAqj0zA7oBJKnGHwev8NX28gaz/khxUHhhQ3nAZJBw7HvlmpIKnLZ0NpFBvQ7XK0LIx7tFm5
lVbp0t+45MDc7JKgw7+spcbwi1gq5JVM+rRsSAxZo7kFpGw7TECicOtTUsbEq1uySfHgbKU4+7XV
tsbeiELz1UXpfRQ2CHXI0E3Y8X19s01SuZQ3//AKWP+9qNbOCVNbqz8LOI1xTqHs3ncfJ3+dANvx
pu4iTdsx1cxCndkNNfUTlXPs27i+ZOYmAHRZVAKrZjsYfq8TZOina/BlWKDNEL/J5lQF3XtvYyp4
i9tGGG14vFBQhKoAu87ev61K8JXvSiqpFSA6dN0pfq4niVqhVFSaGisxZeAZUL57d2VMFpSlABL0
MwmPeWnc+cfYODgD5Ucxyd+WpbG9VWz/loQVi2MwPsjaOPLYGr91YAI67N8ut5151/5I/2/+QT9H
Hk4weLcc9cMjySFvBIFI1hH1X63YPApNyqgVy3dRphpVxQQaBOfyjFZnSDKIKbJQwzorznD+AYWU
UHuXnAWMwHhBa8zodbJwqG71AcURdkJdMnhrWYmZNlkV/qk90vPjISCpvh0k0Lf4OkUxYtqDlH5Q
s9vysf7YtOT8mugwIS2gtBzLpSUSRmnl/6iz8UEPkjVSWqpySijfS3Z0h4AlfNZaKnRwqt+RlPTs
LTa2dDdExQH0mSjYPQM7wdZXQli/OYRyD91tEltx0j2nfs7PLcTkrEjhBubIM0S7HkD9dGs4v9fK
rBLGeCoxSiON7DIE6QjFYuggGz5XI+qvWlCUzdPyt+ECRsNKXSUPCdB/CccVZi/NEx0M49BwbST4
5gYJORrSWI5dyelz+AvyCWFbk9CYLH/11hzK8mFJRTKMGZdqB9LkUis+AOaRCIEuvFt3LTIj+SqZ
hUMf7gKA8IXZDEgVR9emJNY8CHNyfTw96eHIYtDOoJaMY00UFC6n5Q3LkPNh+1prNlxrhB4jZqXa
Xaim0w7z46MMEvRW+yqlqLXRRT8GIV2Kq6KJbE4sMbrBGLj17oA5ycmefD1t3jk7iSz4bu4NCbAH
Y4MV5TH5uMh57hqE6u30zk9NfH23lwhLquc2GIUc5jrWf9ZGi84LoOV+yUaTw56evp0G63vcHVZg
ZIHDgDhZLFlBRPfhB4s6eUYVc8uPUjIfYX1XXDz15Iwn34p7SBsoyS4vkBIsnxRHFz5RDE2MlK3N
92ItrxUNU8jKb1rAJnAfFPZmaaNW0AC7fagU0mScwUL9XoZh+yLmAWXxqviVSchiKPWI/j7Pj76k
HWtyX+VhdcbIa6vkNdQoz0S1go13wo+BRbRnNtoxQR8WOS8ZnrTdk5mJhfAz703uy1FvdwXq9JB+
A2wh1yDMYA/DYMh7PH7hTOr3pQLzpsiZCCaLR4ooG6wIlnzxokked9asB7TWO81zBWjk4etSVJL8
/LHvvhq3Eu46jlORG9cbG23AD/vcD/gYQNYQRR/ksM2+WeWe9Jn2he2/Nb/QsqFCZGyUX62AT+2g
xqXZdymle4rCnA5nRyOpRIuGoyvGuHftkZ3zIyKJdtGC8eqZydLnEFFPpXJjEjgPqkt9Z0HgHozV
2xJHGjPLBylyMyYzuiRalrHz+wKhSHbDUEnGTPoR4prf9TQQIW676/ubtubpn72Q5RKNulhn0ATi
uJZSEQxk+oHZe6vtDB0vQjVuAq3rPg35DvP+bQAX/3WPr9fx1JD4/Miz2y+v7Miaf4CLDnuzdRpT
+qm/EgJUeSS7m+4EcUmcybEKZpcRRvQhwZnRLIPSOTz9TKQBVtVfaSSbT2T1aMI0GClNAFIVWJ0Z
7y+5yFt2+RCXVVPJZgQ7H9dW64BUa7Ieyn1H+e3u+AnwHJKQDfRJaKpR4q380hBVqKRExQzw5CbZ
7i05GkWBXC/fXa4nCBPOzaGuKbjI9ujibnHkOpgdcWySTwHWIl+65weQX6JAffq/4j4tST9Xqkkc
aqMMoaeLmqTVs2ziR0azw5fCxJ8olOX4022KK05e5CqrGTtqiJLNk7lzr24rAZe2DZWnQUB9AKTO
G4QoH5cLa3OF7AIpsBCMdlNCb4Rshngv9OqqBh2q3zrt4+EBfgQSZvp1JHXb+rkn9ByLJ0nADrjM
/cFRP1mki3X3Rtgrg8x/zShPRAGSF0ARMqzSZUE6SywPINQoj977TfaUeZGLE7M7f98dWOo/ZQ2+
Xn0P7vRsEn2FTAXQg1biUvafWoQqWuzT/Bz0BC46KruWPz6kJiVzAylyLF38Kc8mP2BQRd0foemc
d+j0AiZdltJQu9KMFoeYVTvGZMxE5GFpHIYUTI9vzvYnMVCdN7WeSC5nB4K4tjepW4B2DLhUkP5C
hUvzGdgITc1pusGJm259aNx6yNYBA+LvbPNjw39kOB1TfTvxEcrUuk4mTElkXIRAL9F0oemEX5SC
wFJXash57h3xOBCDYnvhjnE67Plw67w83zJi9pBZv8Jxh+ch1sbMjqZg8SLWjuHvOr9AWIFa9OK2
MkI2hpSRAO9tHkW0QRAZDK2F5gyTkpss0zTN229POHyb5Yq91t3VMCm2KJvGs9KLvSVeHfiBMM52
akDLt4kje0fG7/9jQoChMVxTYu9Zp07pt0RyhWPMY//e5CpOzzo184mk1kHaALplZfgr10wDD7ob
PZwB8QNh2cDqmZUAKBgGxKjcSJBYzYCGYYF1i+dxZnsHcSOKWTfbFIOgk/xclZPKKzm8lj/3iu+T
SiKCchgf15a6J9N0r5xgstGrjQjU/+iKV0O+ZM4+l3WdFApNHWDkpAmRlJFFhm0vL1CjwTxEzbn7
aHopHhOjB15jmrNkVsk3YC0EOPWxx6faGyDmxBEPytMSWbL2WCreZ2s8hs8Y5evnKr7cUCCBpAbl
pp1fz4i33/LaMI+qPwjrx+aM2LDHBtzFnGnyCce0b0gcz8K1xacEQpWan0S5m1exp7RRYOTjKWNS
UqhepcWS6Rpamdcupio1omGz/D+wwy/vROU93VKoD1FYgBzgFXbbWY2JKt9W99bJrxvpYZHz9/fj
6cSYTpIyPDDluVMa5mUuzAJkrqyHpdiG9ZWKTTa0wwclMgb0QyiLGy+BeTI9ERkZrlT8j9aMKE2t
ZZgHN9gEAgD3d6Vg6jWBFqcL4I4grvXEnGGI5wy5ngjVh8q/9dQaCh2roZ4qpf5HiBko11Fe3nyF
9qFh/AnrdjAlCpNamDZIyyq7Xra+CK9e8S8g9at2pHGgh0rKXoof/1nUpzZ3M7bZnSsxE+KHbazL
plvUqVEsST51fD5dl/XnoQs+OhCCmkw2Vb8goPzQAxuBwOzpHhWuvyxpATR9dEjb6Bt8C6OtJTJ5
yCuu3A6zZM6lrSW31r6HrmgiC5aOznh501EPIdDvfv7iUCnltx43nCmk/ULdM0rOPclvJ+97DkR8
euni4KBPIg2qnd9QdMcwmRUvsJfXNfyOXobWVaNLphDgjchR1ctlpUxJx3KW0xy2Fr3ikY2dYutY
16CeitZlhzEWY4abWjAXSI37VSDmyKoedzlsXVTpyux6i1F4aMs8ldAo4ltlAQ3JuGLW/gdWzuyi
S6ffSb0g+wi0FItBsOll6YUtyLia3SRRhubxLp0+gWf9oy2Oe6cxhbIjLD6z6DLFNCKj70CXZT0X
TepD3py6c2cIeAbDBX4sF1HJT3FrorJOkIzrq0HyWw6xbD6kKpGOyhK+JW7ylpfQTW6HIyWlHvSv
O605iY3mBQg0ajt2MVQB2REFSdrOncbFE/2AIkhuL6vWTNl9hTYKoI+o5gmlC+2EQozA33L6F6yr
OIgWtTjo+RoslUNupHwcuHfYlgqrgdj0ZOku6qO8J5pb16dZFcJhaltHanGaL+cOCT8xA+OVPJni
sUv3cnjoc6lRGrLaJL92/x+G3EfPb2Ab7EfsG/STFTXP781Yl8GRJzqXBBOiixtdt/8GYlbPhtR/
Wfu8YbxtaZZ0cWkWN0f8gGAqvsBBR7FJqjRd867FHtRVKMY5SrYnx1C6yiX6ROiVmY7gGpD5DIGn
YY23w5r58kh+4gVNGAmfKQLqnGQwRGyNGWL9sfbcT2iNAtP8jO0GrVuO/jzjY51915o2rKoErzF1
bzSKiAVWJAOG03TWxKCmwaEvWLCLJrnAm3mWOVDqbrpc3LWptfwzNVI4K8TuZJbgkUw4UyT0wNiS
NvrSaCqrbC7n36ZMAqgAVAdUN1cNRxXoTfahXgynTSHOQQgVFiusq9XT2+o35dRBYowUHt8kfXac
hz/e62/i6P+vrkFXbDWQUj+0I6/gpw+fHRTrFJmDuQ8llFmpvVNa+D0q7RbJClKxACaejYFf8RM5
9narB76QiU5fAhN41AMsipgR8IOtG1vJHTV72TRW34zW69IY1COH3Hp6+weyqqRuKyiXXIfHJe91
3We887F3UvBsjUKJ6jJ/QYWev1xVstuDFFPRy7zXsAvEfZgo5n4MVki7GakuyqN+jSLIDxm8fTFk
uuTfhkJB4CpqiMad3fAW8QlPaHn+udt2Khsw8PSFFaBM1YS8aXwzBcuRBQRq31hsuBKyTz58+1Y9
Y/K6l+8NJd0l/39AEHSCdj+27spaPYvZdHSI6w5lXcJDmL76atnkZ7ZaCUWtA5IIu8pinjvEAox/
89iKjDgTwi9ZASMaU/pp7S9DMdukSkrO/BVbhJE/VIlEs7wJTTHCTJFJLl6L7wzuEGLJJs1or0P/
j0nb+Oz+ll5Q1nA7ppItXWkSVNaqzRzSdfMMQhYJ5vps5f9agng0OorRDAoQphUBF2ZqN/hn5Ej4
6aXq/Pq3FKTNs37Cd0ma2xdxnlTJ71hPXnibV6NpR+u2n4DpRv8kmYtPcbi3a9GZYLMnEsFhAKAc
eTeGzc0atmdcThWEly1eCl3psuOpaVvuMGs7aYJyt0MZ/iHI10z3eY2zl+LNFzCTmWSBag0Y+abW
IhijdTKP5MHSJFGwEWWKAt6sRfOlghE1gJrcQYykAXnKCcP9hfNh9QRowNHRoWAtG21dV1/aBCNy
WB4d2115VVShHZtlVzripD8cwlqXeihxmkasDe7+bOhgZ9WhObiQQORs6i3RjDNG3CauG/MNGa9q
W1JBZC2MeAQD9dpzVTVfgZD59bUhGiBR0c94OirIuQfivzCRZ3T+eYVbj3eMMmV0JlhqRSB+yyL4
iDP/T1nroO00l31VptnNdL5sxpB5aQ7RkycMMK3MXDcm8QKL0O+yyV8wkkYv2ybiqKvahfXjdhhQ
IEG++pOKCP49QCcJvUqV5EmD/MEPJUKfqDw7vd/x98pp37FupdKAga2liAguD6DUFmhGYdMbCqJH
lZQMb7pzKgvJrVwRPVTosAHLvOPxGMsvvSIG/jUylqnXD0WjnvhTtfimUxVbjDH/9/gCeXowLL0A
+Lhu9NMb7NR+uJKahHBuTpJisxh88tN5qlx5gL9IXuE+059sXoFjEpVxKKgqL8awtgygnfRKfrNa
+mN5BQ6JF95HoRDncQ5FvV3mjy5a4aH1Iadqin3VzuRUhshi7qcpoBMfCx7YpmGhLR1ftuI33cvY
Ir6m0NSCIDM4LwkR88fmQwafxUlK1L6JMkDxvcgua5yIRFWkR//w9xvkFCnO3YTZ2AmDAkRuUAge
9N4+g1Nq+JPmzBUO6Jsu0Aotbt8LMmBXuRyqFYaNoUo8ORS4uEa9eDRcNDTNQbz8minAbye6KCaG
Bi9a3SB0d7Q078OhjC6BL5+WdqfEduFlL16I+gCifF21aJ0ih4ZfeV7VD/BKyuqAobY4oqwkn/0+
rngdRWYUUPY88963Mp0nUsIm0SuhmvSZqI0ObpL3w+3sDvRZNgug+XT3Xy34mbEWXVD/qAzLLGxO
5Si++I9YfeX0Ece7p/qdX4+pDNdPHOyw027uBZ8yRoqDyf06ldvxtbT1rc2AOF4CzPyC7mEef0/U
gs7jTY8/sAgr1r2sbhBZJVdZ/fliEC2hddRBl0PjfrBVJTA1zXB5Oq/629lJAs8jM+E2f65jhQgk
p1heUBC1vnadC7Ofga3sh6Ub5gqvoRbf7VAxMV/CCp2J3HwgZkZlMNU3PVoqb4McqQ7s0nbWkBrI
UhpmKaIOYYTR2z8kEmsTfZiey2Qz2M0PEMl+O3zq2TdOKSCE/XD3w1JPBSlwD+XhfQ3RbzNUgXtf
/mINutDXl961jhAmVklNvbnSSSUJM4tvucQF8o4dnURBQN31kOCxGFA6r+NXA8YgJ6fQX4sPEwKW
E8DI8+imyIs3YhAMit8VUuOzkzXfCimq5fUppIKxxva4ZTUup+nMkY8rrkKJkawUwy2qTl88z2Nc
ejDSkYWZIAhKgDeXyjgwCXdPAVjh/D+n0MFLVBc4Zk/lVmnk0sSwusf+1nhIgAynse8F6N8eyZKA
dxqmNyphpemnDT40Cbp2DpOdlLjnwqgjQjRVHpCEV5nQBd3ZZiKqEkJHrx7yMTSic4R5JXRH8aYH
Gx8cZiE0CwF0pf3soUaaEwZV3RUikqjJn3JLO2CkejtlCwyDi+LNE/TMy6hOfHoKDiir+s7nzDm6
6ceElwdhx/Xygq4rrhm6YsQOewsxly2LvMnc66d2TQJLswXs57L5YhlM7xBXDsxrvxfucAAmSIRB
WCiE8Xd4zQ6Ln/SFZWY+2yYiUcd86C2zdf5HVsRTcXxchXae36QUYgtlAVzUFF4ySfeV0NDENHFM
CICm7aYFCjL6qN0TAEu9M4VnGHgF7bCLwGYYuxfPEWgsyvpY80q+/H1dvt9899NPsPBjnXvUSu9W
BxMB2qKYcRWotHS0wRly64M1TUDoarII+UdI5/CVh1/rpdN39cFDjETKH2eD4VFRx69HTkT4TbJP
2jmcD5NdBofX23Hcfg8XPcnJ9ZztmVUQNppvFvVjE2tOrw+YcLkJM3KV4NDeU9l6YCS2czYHIu/S
H4Y8YBEbDquuh79cFcDtIbbEsiR5yWSEvLBRwCd85GU2SlnGQbVOxlxFwmtdno5loauYeUIDGjhp
8G6TGXOVAuhzo9vzX59X46Rwh5+MIGM+V37O5dZkmh2AOavwG1jS6breULAabHbMLZJeM8t/Rv0h
Xv6hvnP0kCzX30Knz2R/AbeUuYbSBADVUXxndoq0apK5baourv4n7ByZtDcfRIopT3Fc+0H1OF9J
ako4YxLpIc3HTahGd53GY97WN2hpOeUcnRWpab3X3zGP4R3q2qicqxAP4QDKuJfz8OS96sFXQkyk
g7xjcn2saJK86B64yxoQZY0JCdLJmQ6xUfaR73PeIa4qkjSOpi+XW5VQgIHLYSGEm88Dx3VFOUe2
EM/QW8eHozdFqHuLCpTkB1dGTx0/qiADHR8s2JJfPIj6wxAgTvDOpJJi+fDTvMbqCNonKrqus+1x
aoEUjswcrYz4GFX3UdVIOpMj7MmfhP8LKd3UqLp4g8ukiZ/oMtYAmhxF7k9oLC3w5AvPxOFBxl/g
HW+sW9NlG++TXvkaXYC2tXrHSJbrYfTWm9C/tKXc891udIIxMp2ZkYjpBEVxlCkP266xS7MCHpcL
YcLH6pwhAD8oSfdS1P30fgzDp5CKJsKFjnh5lJJJ60ucOzKJ6LTMOz3sQwMOcrpPMzrqHXulKhlH
uFKcejQ7NDOWYAwUdIRkX7ngSkh7RvL1ma5/C4i/EstkfwQl2vxWqoyLtKCm34MPKVdL9NY5K1aT
owxe8yv52RRtT31gk52+c5wunB0N1+AVUDRZYrRrfa2AC97JPsTqO0oLfHe5JgwJ99R/8EOUgNC3
+Y8bErASSTuPiLI13mqW12zG2YDfvj3LsOm9nDxUwNj+vL6+QxeMOV6l/9VQFH1Y6SUThRJJumhi
jHEOPEbhbf7qBcUTZtNWDGJGNyslNoAtTVR61B02rieg+zE4EeG/54WL2MaoCjUyDUVcYbsV00lg
5TNsyH6HWQYZCXcMT/pSFH6J7nI6FrtO9D67ET1J2QnsikVpY+ZmuLDVKidWQzPHhnBhxMy5LxsE
xtJ6j95fN7Wl5mRzGdkW12lBHhVUGXuUV+MJkKkjnMYc0WYv+jjc7HbIV1ot6aLZEp9HHLCvu3uI
geVpP2fu/XXinUrsIeTBRz1bdeiquMnvXKxbUxw/4rOb/RQqc2IegmBcSll+hwpS6e52CUyOydg7
/ALJpiX/1247qtrMZsNJU7rB8mxyxHMM0oHUHkayGx4CAEI+aOoSk263WFt2J71xVtOyay4Ea35b
KRVwRBFOs06KX7VTZ7jg6uyRS0OjudJ4NEeyjE5GCkDOXQXTSZFZJyU+/XAwgi/hRtgcvmwK/mUm
evG4HVX8IwzatOHag+aMNO/vyQ2bkEsrXXtIUavGJoFMvPaKQjurhjG+8l+g25b9QpDuHp8ukA40
xMo6E3NSAuWTApl0prwUL5X1SkbCtI3I5zLBit3D5Ujbl4qZdadvLwUMN2nMknmxMcSjgq4lDaOn
M4kFGf2foiawC7U6ip8rIODuaQLLcUPqUwflbkAD40JToLNNiqttG3pvlpYmDf9HSE6v0dXXpojD
KeEmMTbDx44EWTX/ij1jYOMAEtLT3HwZ5Kl8EdHpzK2NvfOtTxDFcx0xIsnRdDgi0bkE63WDVpEg
iaAhgOlGRTBjGx9ABhX5K4rfev2JrVeNtHU75iJNS3kb1J7WVL3BFUkwRXfGd0EJHRWwDkEL8yDE
4hx9xqi7Q4tnAIQqaTHkgzIbrj/ifgInE/CnsSRKqKbnCyslOoHJVSRUqnq8nnQgYhzhKkWluV2V
xmQAfW+ysYiIcpGEWVchF2iO74xaWjIsTSKKR1DHuNwXB5BDCyo0v7GiRm4XJZVcJ5SUmYq1lARB
YpmSbeb3iLUwMsRm9uOmnkq5x+7zazgKqUpR7QbjEhYy4IHaBPjFMcINHHajOmHCPZiJfMelifvd
wADyIuIpfIYMC520V5KXIyGsbVFFOnj24T5mR5FDKWUFRw4smf8nFDWsGA5JX9E09ZE8pEfWGgRP
ApQzFE6EU43+MSTW/yuECGUNh3tEW/pbFkD7Qwu7E0AMyDRUd/csXzURLou2E3s/BFKFOnh2Sqiw
ZIjT+0XfB/QLM0meuVw/cIUro2oTSXAbzbSeNB2aMfdGzi06VbWX55v6Gu7lna40nHET/vPSCB6U
d4U8dmPbk6VNmufaDKaWHXg7ItaqM/Egw9WaPCoor/0sCwoMypWKoyhTgffVAz8CRT4s0f4uCKDL
qCGzUor0QysphrPLHs/+KCODsdi86pBsmr8sAU2rPBIuWicsy7WbyLhBaziYvPDOdaYEDykpTpC4
025hX2FMdn+FhM4iAfskTVskWuisKyt3FjZS7WzZ6NlFim4m9uRbSeo3DQHsl9f/SSAip3ceXX7F
qewiIRZP6nIHXRMAvuiaEuKeBEn91iMl8O4ne6TV0mTqjpWU8VmDeZZF4C98DdtiYQBidTdtXiag
wur3rKHWGtNvC6lzlgwZsVw/f2of1gcspMAAFo3SkES/Uvkj0Kf2u0xlMy3sm3av/DLOgbgEOfTn
d8vjITKIih9T1rPD1T6XVzDJ2SLx/jGvDrETuz7CtKTkFnlLSkjOJRZlgmUk52dlml5PvGA+niUn
xbUaHcXt6q/OX8wvj2SSZVFlBIAV8Ab2xZERUSy9U5oMx9X1Z5LK1545Vdh/BaS0GNlexoo5lbPm
sDCUGgnONkmssbYLaPXW02/mjVN6liiOKd4FuGsKCcdPC50Wpr4maN4ky62TOpswqL5bxhnC6zx1
6EPkwTV74ZQ45TU2Cn4pVUr8xNdPjxgsIgem9EQJZIoJdzr0CokwZcBwwWJuAanhL8ZTihh1eM8n
al32+EVwYScQlDCNSKooF/N+w47v4Lp7cDdmQrV3NnjCiY115y7K6pdm80/IUtayDr68IdDNg9q5
yJUcMtpjahpODZ2Kq6QI/lxzqDvIzWiwJxMR9HUKsa+60Vp8pDRU0838cuDm9D7xMDTJRguAdCd+
GHUbkql51VThOXGgij7lIYjOFM8up37fhaN/q9us4QPtmPzoC/YyE7vJUv8YsrOJlkT1Ce4LRn9Y
G2molwpo1S0bmj7B3tOKavUCGN3PzHxiaQbY/miwrlsxUSn0NYWF46zSb9F+0mU9vwjRVdxyggsT
tCPfHEA0iaRXrk4abWNsslJDm5gZQgDj92GquIhG3GWKghysYqqxVGyklzNwWt/uwHYH4QrXLGmA
1GW2fPwdK5GUgGbvQKhYTVoHK3UWEUobsj71EXA9vWqkhZUPvI39T1vwGBkiEt00uSGN/o9T1Hrc
dA49h4rPSyle2bEhb6oA/VFibfA1KCFv8P7zQqGwP19yMJYpOTICnigtU8M5HV9myeYlmFMe4CFf
D/2Oeree4sGfIVMyEMdbx9iQUwzxYvAiHYzHrpvz3O7DUiTEzsvVtMq8ocsWi4VDDEDHaUYL+p2J
POL2dpx839iqFBnESimHF6MU47fh43uhBzClEJldmVLY2G4Y1Mjb88sls1RlfR5esGl/91li/2mz
zM3ECJocxACwThH4y+vEfcSSfsOjyejO/W5FtkBgs5p93I9y+tWxUUw9OcoyNukJPWkgwMj0vyAS
iHAGnZf8WQrvy6UJsVnynliGYcWqU06Vp3fZx1gVrC33BlmgluPEdIsjq7r+U9MHBeiMOgco2tcs
45x+5WfdKMibgtznz3qQxztst8fAMPwDy1IIn15yu6MtnI9W748a8eFuuTkJ1uzT5QDzveMi75TP
gxKc1h1bD5iBJO4KK9XW9I6ToO4j61cGqV2PZIiJ8fJBmoaBKvnCi7YhRq3d7CZ4h0CVVDSBr1nJ
vRHf15nhvXsz5Ah6Ew9hsLAucuOQvNHN4IWgHNxUWQdsUqfkRj9b+UbVW85gDwtdg49xirWhvYjf
5bllWTNDDZ+AVQpZjb169yOTGtC2+HnviVOr57e0zJIZJXAdo/+ZpsYcqgy5won/WSQ8rMe25Jof
F+cM1KUOlmmRT1oJC+7kAVvZcfVxlC/LlBib80pPgCmN+oyHjik+olHFCHIIg8THR1O2mxKHPQAE
vBResr+5MDhGhpE0xztnKQK3zAr76zCkU7kF4tE/tOceHPP0E+s88c+YcFKkLYCjmweRQloqoEQw
IR/wCwFYG/2FxHc6HG3WyChHYy99PTH+QFd/xOQHe1nsJ+OTlI3j6KaJUMc5OP9gZi+YKco6Jv23
vZ/gEa14cU86IhwWo1K4QItJF72iHL5VdpWuixATuTmaXTpoRJariQbp2is2F+2DEUWNs/gRvG6Q
01UBS4/Vn8rlDfPUNWIyOYpMJbqba2DRoXQuu+IGqXRMW1jREcfHn/g4X0TPga+pmKa+sjjGE+Q1
tbMwBdmCHVAAJjOKLqNQacQnvh0L1+iHcObnnkyDQvDn2rAfJvm/BZGD3yb2hL/WlRiD2AjeqakO
XQXFv3fwvdcYpdT4jWkxwiOSuDoxjBY/jMotEs3DfxxZGQp2XhcHkVg0YAqhLrqZmKp1RJvj+I+g
x+pdxFdPqCIWFFTvS1iQlkbKccIs/gDZ8EkT59ik0CLafq/rFZihKW7yXvEN5e5kSMKK2bQT90ny
2DVZdhybYu1DFiybzxjpDlfkIRimw/nO/E6MRd3EAUI6tXv6NjRILWnAfCcNq8Vrdw/oMxMsFM6W
GY/bzWH64czC7rIh9ur+wqlRU5ememe7pUz304NHJ1fPf/yDot4iWFEC4uC8Jw6XVydfqMgz3yil
oMFemwbAgSc3kbr4jOG44HoCEMMKPCJcWfsoKqY3jqwSUJc4KuQEpp6UKT5fcrk4gZNd65nxRsnA
aI9WkdOnODdKqxYxzPhsEdE4ba2gscdHNd5isFr6ZBosYZmVjsFrU6SwzrQqHg5n+BCiSCA2LapA
P6AdCsHq9Qhwh7ReWMIzqKNadkd5x7bYto2SVpfek3nlolVzD2KXcab3hibn7Mdgj1r1fWNWep5Y
nE/IKO3hZVVRzGWa9rkt9r4bC7UJ4JMGS6yims/xPoEqtBGUzqlFX0FiydKWHMgHfcKykpmcvDo7
xxYkq4u+/5T6yOVeALVv4KCvzQ8nykyiovuKQTiXRmHbL99cvbxm3dwJLbX4fHt97JvZA9/2G/4v
+dTAkfK+gaPebELRidUp8FudxI4SJ4H2OH8EpXz5n3vd25+8OLLsnCnxcyqynCpMqUypzaA74mcM
16WE4akgs9+zDnvoi4GnJGzzQVJQnRuJeAOTluFohLOtWlIBBrIeybv85CB8X3ilHVroWXd9za5q
P93VSygtN1/FTGlMbyPB15xXGDHtlC6X/QXS/KEtJcJYi9UkZ0bWDrANidgiZzYzUMghR8gl7cCF
hHcE/LpGAJzbox7PLKTN/BEXm9LHWtG3GIKnr9YRuY6woOwmx3upbNEqObB//YVguEbv8QvTTy//
qUu6nfquDk32n9JYXSkSJEcncb18EuMK5CYz82hYvIIL6G8aAOxZ4KtHB5ZkJT7QlA4wA127x9bE
wKHDl2HAiNOSmtBtlyqzQduNGn7+bielFs1PyYYxQBBgl8UTv4mE5HGxjAIxhRPjjqXErC3CTFLO
Nuw/lxOqxD8Yfsz2MpkU/cXvHhmLtqLOq2Kmrj3sEaIoMUiFbiy3eoQ/U/BgaoZV+D8le+o56m9r
YJaQViOv/WUzQyHTenIPZ4Zb5vzZsmZsj3S99AXFIM7h+OwIQg8GlRmYqjXe7BiD6nfKyYfhGSj5
JoBMiZUBuS1NtBiWseUyDYQJD85liTb6lh8MRbaYa+chI+EdLNpzEgQzDzzkagAvtiJjX/E3VACv
DUYevn41a9cEn/+cGZ8kjKbQUMygmXX2vaOI6Q5E7YV427snAYtsYGWM2/gCfcaHvAsWHJLakghx
Qaa+Drs+Dm+nC5HZNf0hSrn0oLPy56ShaVzKnnU6lwa6Jcf9Vn6S6/DmRIyHtYa5EigCmb+JJnx5
KgVeGQnmGPllGKxcDiBReaWRD/U+iGXwtGXuZqYTa0gJzBSajEuC60uirPWOnwz62bpGJwsbVUmO
9x0GnzK45gBtFr1401RHg2fFoixrwM5LJ/S7xJ+LHMU73CWnzIdc7re22mTpRucSdD0HE5zCiCpG
47p5WPXIFzjYW/cLSaK2L3qKoSCwgOJXZ1wyYU9E+BUseZm90i9LOF4II0tsNGfpdqtMC80PYUNy
FqaVTQM32jQ2ssHbXQgHr849En995XVXSzI3QjruqIj8tjfnsIc3XMNJmhbP+hvcZJQQDljyId09
EFLQhou3rD+SUQ4ohIXAKIWvEMLAYCM33IC/6Lu7uJ1ZDic/4XQ+j6Wr+uxWBdGCXloFq2PWxc13
d4e6k5qElD/EZ7x377c8y01sWCOTjaCWcxOaFEPou8TI5NVdQmezbc20NqEiTnyO4QkX+wMfUa6O
F0dCm4zVH0Zd6sg7XbILJGCDC+cqdEdH281ej5pR+klVJgQkBQnkJ6oK6WZHp5hCV/57+59j4oML
ZEOrHEEDrl5sKs6KMStF9HPx2AG6Mz0/4JZ46TjY2F6+XQifrs4I2P57Zdj5wLMz9O74IWBbJI1k
53h3+rZHurO8HhDF0eMLBksHybkf2zaVYk9Z0wi5Z6WNq8nJ2KRAEVVZTIJbvh4Jm8H1cUTwPQrL
Gbw6Y9ldQmCHOQZQhltQL+isFtK9BUuzcaHXsiajfz1fr9DCusqikf/HCZzuCoz64xwetqGXnHrY
6WUoSltYn5JWBidkObgRaQyGyOwgcEMasNs+GZXclEQvqd10CJHiSup32/E6fkuI2LCR4BxbGYAH
/E/4UrPOZmpy5xZij0tXJJbNb870Bt88+3WeqJipyZ4Ze3ktOicptsK/cYA0afPO/SfNtH+RLpy/
2KLT2EzCNhSwXSWeqbodSIpa+L0I0XAg1MEUzmqTYfnJBEcjWSprOaHgLyj3TjqyzUo7Uy1Qk4v7
KIGhgf8V1D3pe8as4kFyLn/YGwku8A0myfSAMtzy4qQ1hHnFo053HTW5jCje63eH3DFIOWWK+CBu
btsfWF2P7hxnL9Nj30jZfnz7hBO5USqLMMN85e5u67kv7xndZIjTZejjIjZCHcAHkNGsxhmJBl5q
JYTyheYyCrXVgkiUjwDnyRvtIS0UsJ79mncDSjnNN2pTIANNXBHlX1+aTeADA0ZfPifXjG95kwD+
EPBdvQHpbkCOv0yfH1HjNwNs7gvcIY8b7mHU4GOZhDb1YxwVNONw7MDyHN3JT+x9GG1GlgxB9Fzv
NAplJF7x1XlvvuKX6CRE+W9g8jkDhXT05XCf+I/qoHMaGViKyxt5f2CYvI/MNrlplafzkAuwQQUA
GxYfnc2B5ng8Mo1+vHl2LTG7pphmaSdqtoK1tMJHHwkyTgC7wHczgKuWCG6/+37yv44hGhT2q02R
CaaqzAW147mFCewr5UcSy79kleCxKbisGIkSpL/rcmFUQRX0lBrO0j9eVsPER8HZksi+IW7ShC4/
b7t99d69yG2i5KdJx/2D35Pezs6Efbmf82gHMUKIJlyWSKz7UgWAf9qctmcjrIaBuv7ML6DVZ7qx
Yfa3GnowVayMoAP5Xr5ZoKLXeDDzV6UfnoaAsGUv+WGMxUMY20CEnrBjDAMxF88oGBLKq+iwqDBb
AchfthbGT7GHAGz8yTOp9znvh8qHc+CiPeSBun/skND3lKKj6brqmlI5OKjyPkKKtapYw3G6Sht4
dCKepNfHWo7lz2166l9iu98JdW46oHPXve8aRfNsp9j0wXvTnODOmfWPAhMmdbtSniSVx0Qgk/+L
7g/JNK8kIzv7CiEI24cj1JCgv1Kq38vQoILgvmZINxLSBU2/nFcYDOCTKV5IE9+QjuJwdhXg8I3m
bbqdYuSeEuflnuVcgYOIqWRZzJFWcXxI3HHwfW4DJyNXJ1sN2tu+oqtH4OPYtJiQfaKmdk4f7Gr7
Je17sZUrwK+ZEmZcHSKRQk5Uio15cHP6v3mOzNl8DfEEg+0u2XHHKCOX2hmKWVFp7BotP3ISBzET
BIZpZCuXOzkHuJT0OLOpEY/Y/vqoX7zWB7CKXLx+Cqf2AiVviMMw5SWXvHT3nJxuMUDxDZOLMUuZ
YRAMt3jp0gCesNB/XoMInK3mo1a6+p0NihYke4z4wEABQK5nnyRgYJibs1QD31UP77h1OeJpRwYs
I8SDln/lXYSCgLHn/mTtXaN2fQ36Gb3ZcqDtg+YpR1XLc7tcSC5JH0cji+5WYs0Xx8aZW5/Btay+
hHWRIYv+I/kU7Prwpfy2KC+jao6qv1vhzt0Q+IEmx2l9mtuu2bVmR9fHYSyjlRbFNDFKfqphrngv
1q+FrYOf/isQGcearpXopDyc73DQf7pebVPUT6Ob2MEFl0lT5ArLps/jTuLQ7A6XrE1vlwb2HRHi
mXX4I3P9qyQWXAJnEsvlX5CvJYbo82bLmCrOonusNliVcHWW3iirFKI4lhlJkYRm9HKg9miZ9PXi
o3K3IPGB4RdWEL4zDUpi04/+lBlcc2gM9TeSvnGeZxHYPUUjnlrlxNY7laKVXBUO66m3ZUi0Vbfn
Bi21DGKpa/RpfQHxQyfDDseTSjUqJPxLXFVEEcV/mt0TH/cwaki95KPaa3oGkubt45IFhWqjNJUB
2GU3vkD0tyliPzortRVqSClw3w9Mxq7cQ8n3J4LIzDAe77FTlop4HffCfquyrtqSiAeHKw+Bg9rS
2VTZCq0A2ijljYUQO4VrVBMl2fBOg0dUTosimtcYGghy+y/3GP3ahdbtByRd9+qTpycz2Xx7JR1E
3/Xva05pZwvKu7VFtMD+L6qurPtEuRQp5TREshrtenKMchS1UUjlh3/ncjlIqF2SfwCjRi8vNlUE
2N+gsRo5eyRfMJmrmzpJZYtONP+Gk7dEZ/+qyeYiu82CspVzEr8yuq1sJgAdzGTMvlOAzDURccn2
MBEPcuuRcP3yVIanwCk2h3MJQfGJ3n/GW415ZGSgu3KPFg9l2mvtL21PUVTf7FRe1ThhShf4WbRn
wFKz1N8pqG3ET6xSA0PYZv69O6vxHBHE2CsVOrUnEE8w5o95VzGpEDkngMM8HAXUwikEGyQEhUWG
rBTbF8SpliWjCFKm+YErK2R+/F83wx6lAWyOmgmgwzt8qUVw9kENv5Jw5X02qUF153j2mzQ0B8M8
G15S0ZvkKzdj4xGpOMHRgvBF1yOHPj8xuH5qNLT7bnSBO5vmBGmkw83VwomwhAHTQcUmVVh7b7+7
lXwUmwKAxWQbtgBLeeDp4Ce4mhNQynfnhoq9gIA4uMQggoynm53kLCQMawO82+dtd56lhmokHT9h
IBoiW7w6oC3BycCd3iJY19mltCgp8yI/gmrA4cJaGBNSShIpw4+9ksXjxCNgL/Is04ZB1GTccMFJ
jUYXG/wTfUSTmm321Ku1WNRg5VMnT/QTZkYcKR3jkhWhJRytfrltO6hKWmHzaq6QGyLoja409yZw
UM7jv66r+9+YDSj346n584dgqFxO06UjVaY5H66Z2ZsLmyEswnAbos1bdigv7n+m0rQqK38wbu4e
/n2MmtlttsUctShcyr7A2DvG/VR0gDRgezHOQPjtMfD3Aer9D0j6rF+A8pJZEsk+wrmnN+zdyF7p
aTmXvLSs7y5H6rxujbBvHQHSmIH1EOMB5BcreBXyUdlNcajUjVxf4OOrCZ+o5eZ7igrb5PKhZvkc
vv4YWgLBsFdfVMbkEed3IUr7y43Mnl55Y2j/H0kiQYoASSiu0LjtMT4E9WYGPd3HmJzt/wrEYCrL
BpIO51ZpDr+h+K1weVdzxYldkFfeZULRvxlxcz02oqHbKcYdpNKyXXDjsHmgIwCZ5MPcVj+GPJXd
V8r/ocKeY2o/41UlkvY3km4m91TnlruMTNhjhYrJ/aesiPCzkBPb4oGwYiceoP/yzAqQjGWSglfl
X8rb60yiiASAq60/r73yLuekkFaeq4N4y8WwUc+utyScuBqYyC8Oieg4y3MBc8vss0zjMqCYoJCZ
2BfUuKT9yX4SH4ytJ5wWI7Yg+8QuDufE8MIgEMnpHcT1Qw8DLkhrT7hSPxb2KYDbqa8q/lWVtOUQ
IyfDVxYHhZc2NlHxxeS8HAjOFbW12HQI8wa3hA1sIjpLMKp2YVCtmGwWt3mrHQDx1OJobo20FZqP
jFAYBHRpBOaNHtE7PxxSMguprv99eVJ0cBJO2FuGfHcZNDKVeGLfdS6AevYTn6VqOute6yDyp5ej
s0xa1DF6FvBD3GXeN4yfe4CDI8ku4L55ScQYrW2bIzlk8hBUf/NRnDn55ST/EvcXATsh75jD0zWm
XgdV8adZPTDnWCibildGfMDq/PBoiRgGw6Tt08ZYDH9W1mnQ159WsBnoNp6aU0Zvik4gpyZPWTMB
RPGZ1a8qEv6Qzsk6nchIr1v18Zxj8gDDBnr0YVV5fEV7K7IYNBWKjVTSnnBsBLF7bNbjLYCbIMsb
jjSlZt/3oIQCAD/RCln/4OyL/j2QarKOgdqQM8Y/9nUEmxtFGKlNTiMzb/B83aflZgGif+e/9jmJ
2CmCqcm9Wm6dJF86ZNLAJsLxCpZAGYgebUfUIMkjGIJBDfgvRXJ8bwyXzzwyUNt6poTDFPkB55Hx
IF5snwChy9MwX57OTIMPAVaB3N0b233DDB8qPME6H14BRUPDeW5qgAaeQWm58VdoxRa/KksE6RST
hjKd9DZh6BSm9B8b+d/7osuugR7qbNfHfE/TguMTXjoF8zUeRuMxXzFtJ299JLuGPOnV4uZSQFfO
VPQLzVj0vG4MCIfJCs9IVsk7WZEvtpqmMPFR8kCfVGpI6s0P1WNTv6INZqKzaH2NxvJ4FLFXjaXp
GVw8l4HbuhqIbVicxcQhkcz3UZdwH5SY6dQctl7bAXIti6z2baHAxLlnRnQOsjG/qBiD+X0b5tox
cYfMS5JXF5/a0/pZ9C6eWxC6UfERyXRT+tShZuLHA98ip4NuyoCWNMglGHjgwpz+K1Z36KynV6Vp
VViy48KZViuJonN0lM9xQBJDFg6RZmg10Km8MJwkos1QCD7IcnqHUfvSo2fz0h/Q/5UfA9Vt8Vrn
MGP9KeICcfMWgxiqDCUsZUaKyGH54z7VeIWZP8HLuL0tFV+KvqlbOXyT0CC0euqtbIbCHGeinNcV
RFH4RHbSeiLoNiY91qsYEvsZ7bE+hT7J8MSh5lVKTJnFsTaslfS4laBRSkJJsYsm88l0SDWHW//n
Yz7So0s7KkpcPXGELDx4gWNAQIJd0MPccI1AKK4Tr8UgP1/+r8FYxdYvcoxtHpHCV1hodb8cYIPQ
aD7gWF32i1HOD/viE95RpcnA/FzDuGsT/PtJ2teoCVCvcUtz559/N8c67/W98rF5GDn0UWWDIanE
wYzzJuf2BBInFreK2DcnfynR9w4XqrBgK/yKjP+4gdWuToJ2TX3QPCvhn+hAVtIfNsLSRsTt3k4f
GzuLErf3WH/k3MU0XmdDsiwCayMDOdBUBd300y92IYXCeNhDBSTB2Sa1VD242G7X8qewb9CIqwHD
P9QayyCUyhB6ESjcbUTJ/FXf7N3/YIKMMepukKOE2hJhD9x0guc7yv/EDhMTsnPru+gm+aw3quje
MO8IAdIcE9R0dcjAR0lHVnWW7zWiJbflDBcIWYKg6npQfzY27zfv2gk8A+qlcUsOhanbOYn0Mf+g
NZcDtbzsNYu7lcoYCV5VRZCp7LJ41SdkirH/GXVXeILxpqGiBiblOSwBOCFOjo06bzpy3U88RaIX
6u4xZTR+IypXuFPlVdslCXnGEwswTTjno1hMywfI5PLLvWswRtwqmEySiTMiSd9hUqirXSTb52ex
047UKrZUzO0UFEsNLtAzgyR+ph2o22ZSl81okicjrFbV/U0Bkx1N2L3np0IARKH36SRwDJNZVgxJ
7waArYMb9ZmR9gDNfHekNDM6puxgLh86t1EA6MfTogdOxDYAbBjC+VUNxnjA0b6yY1riK1vNjCHp
JdFR2uPwJ2k5wvM4TkiUwstspybvNRXA4aNxHBArsRK7iOTwPKPFc/W7B6X3nU9SGCbXbyfVNJU9
O1FPEWzGi95Wkj7NL4elFwtwxxf389yt+gOp4Xh4ksyUzOlb4bD0veHdxzEGgQemOhjDrJi705Wq
vY86HkvoodX080L9xWRd264u0Q0FJ+MlI96b/PZ3FXnWKFTWMPCFB0O7hySJS4+ToKX+at8n9oZp
dfX0+lzM5dTHAFMjr6D5RFi6QtOUYz8dELm9PXekCO/ECplLaNTYabxhXGf9A0pqeurQ+wnyh22k
p6jX0Mk77ZX0YcTeMfFCIwGE+1Dqenh1Pt72YbkRz3B28QRTPcKJBRgJ2UHw0ZDv2YrA4zwS8woc
SSoy49AWLScuUHxyFQtPTc2pY/k7ofCSqtuGQI8lJ+fHlbtC3tWmuTimIhAG1dO9REYuzXlr9fL0
fNafjDtVl4rXG8WiTAjYaKQQTLjn28BpWM+sr47F4Fl+jg6ZfS0fMA1Hjltx3Q/be3m8XtR/KaEC
+F0viVN4uPZmNw9MrkeJiu8zgzEA6NhiGGzbUvF5pQV9LYmcisB3srcRrLLsyd9lNZU4U6fByXHn
dS/xs9e83bDiYsUipHP16f72PU9tZIWn3sRteB1MN50e9W8mggKDwGbimIaKgKg4zkqLgPTgq3yn
SZYDxPzmu/VPR9EoaI+odaJ/EnyyNCep7WovZd4qJklI1nT2ZdKYOFya2Vz2qamXtzwZvOYTQW4C
VzrVfPM01X4w/YFvxz/1/dOAO7tmR04XYn/hb08VR5yJNUGQVx+d3rLG80Ng9Ikc2jD2yGCBcXcW
hMJTBHKn1Ds46wxtEA6g67ds2lmZJ3W1vt6JPnCyW4YlAEIrG6yKjiIFOShl2O8tVfv+0ea0ITOG
t5+XPKJ02UjdON5RGMNI3Kei1lKNcMTD1YMittmZ8+BhoxnvlNLyunmQtrrD+bnsQxDMW7XxsV9B
fTY5ECh6mvORHWHOXGByGTbRUKvxxhHBVwvwqw5o56Slao+li+RB8amAEbkkzSXeR88o7MmoQELC
62TgaqNZNAk9taplfs9rX4t6m2LYV8xdmUaOvxtwZWhBYdTSMFu2qiQ6OtP63yUt4qM/ehRZXOwn
XvM6MzNnTAfOnhHqcf1XTo6D2Zi1i8wToJVRphNYL2li43Z8diyrrdGXedKJi7f00tukfL9kIwzE
+lQmj3GXfks3fxqfwf/PcRLxz1cOeUp9gZLAy9yqqKq3W8AaLyIiR0XIDaAbPXwrHxdZ3Simc+Pa
gAy0GDrCP6HH2PAaXotc9GquuIhJh1qoGd3W6T8PyBbmbsZK0TrgeVdo+2I5GvkQRd53y2RY1QmG
EROtqvrsmRefn4OdYCTxcgMOeKP1PZyR0uKvnGNjx/5mVQP8zt25ZBQNmf4spOi/o0ZoukoSJ919
YzRBwvVbEyCnGdGn0uU9pyfQbr9uZCEl2lRqKfCUXzctE0QDWd2J0HgA1p6S1YS4K+VzS9J399S9
W2PLNpiN8qdsbdi9aQZHYBg6FQIDK7zCB2iMRedfZsgX4uFGoqPRUO0FmqBuZvv9sPQ02FVp1R8w
0d7qNcMobRtepD277VfU8HCeFYSGO4SqXWeTKiOdLH+HZ+AjxhiiQ9yS7gNxa/jk5hL7h0TPzl16
GLghZwOw2SCOspY/2ngNWlwSKDAmU0ydBhP32Xb9V54WI3hAu6h3B/zVQxJ3VSs9N5mTQgTSAXV4
e8QyaM4ODkAO8KKjz0XP/HLqorbo9icfy5MINxZL7zjkjFwJ/aydV8Ic2WwfQ5sEwlPiEtZ4gFol
OXF8ybIAUhetn9aRoONlTwLw3yvh/LxQ69zXEzZIgqLAnzplUG30V4dwOSTwvLGNSrKSV8y+eB+X
YqtWt1/WCOJWbDHGPuwUFWFXOJNf39UT6nsF0X5XJfIoKh4R+XXIz2EOh+XH7ceg2F/hw3J7Toh1
5XTuYiKYPV0TkHN9CWZy+wY78SZOMEHzpdTewf3prDlz1qIcBMf/v94xONSRKASXXoTNWIUtyCX8
joTuHKboS22HeztVpMTAE0U0r85Do7xOJ82wxkItWsqvt3cwium9+BkH6Iex5p3nIDplj75EJ9XS
cSjoAOaFPuN+m+daCanKHslwWeBvRhdRBsiAdj3v7YZQmiuzpjoncp5sVYsEP/Dhlo1nATdyoJoy
XlyrmjeJVKGe1TOCsEJG7PF0p/DCHcxSI16iUt+CBLteg58XL0lwN4NkzoJefXm6Xu/iJe9UFoyt
TR75yI092JkFidBOYJYQRVoTiNlHOoWaArcyYHkXQp2XzcZ7pw4miZjHqXyF2H5yQCf44uAzb/vn
AlsvxXtOsmexZ5efxYy3lTy1lQ11Npa+ITIPViU2zlpJhg3cfq2U46Q0tpze5vll54GFRjQ8Kxs0
44Lt7oj2Ygcjz8pabrjteK2BiN2hMxCfA2kPMqu0w0kBLSj/bz5Q1c5/DKP9DK7nVqdPSEy5yFCP
7JKHfWEHy/GH3ykWJNC2B9LFZ3ZfSAHdZ+iIjwxjqLXhW1LMYkDbFxUeYP2kpW40QQQHBdyqaPyc
H97uZcudDsnqep2GLWvd0wENtVAzh+FChVRAQ8PGHxvkTj5YD14Sa2YvMOSbpbz4ywE+0BP+9iCn
7+1U4Vw9nPPAd6K8WSNVXj1BgUhpv86z2X3byyi9t/Rv36wJGbAplPefcn19kU1vpYSoWdquOZrW
ofzj9z/Q2H7zZU+BANT6jii2jt0jwA7d/xhI7pp38BmDx/Oxvjisoq4gx31KuX191P4UDwTqmtQp
W0fE3AISrD05IPtHMaUow7QSDoU5fNeJlvHq3qkflXi9Qkz2fRzVvCutmBwhOvA8JkCuaLtU6Eap
z/buwSx9LA/QKDrE4mjtFlQ1f17sFlfE6GH8Sl8GM9c/F474dOLJCgi5QimYrhmP3F1UbBykSgCq
DqJEyHq7WmA9hJZ34+gLwynNZRBM8vpjjA5NLCgh0JVId1EUs36JwkYUwWQiSCQdDHV58BIDLVwo
xmteh1P4r2ISuBiv5t86L6RYwMVV50qnmpQIAURMwoeWNefV1q8HDHs65qP/w+UvOPEFfn0CwJ++
dyC0xaUHMx2fxJBqaNrmolmOiVG43tdKSXJ8S08yJmSWvJ8USXBTGJAO4I0I3m57J3SRir8US478
4Q5fJuUS6bOmnGlCxbA9zkpMsWV/qgiSsxuL3hzJfz/qCc1RN/x+jehqtJvNzKcHgNMCdR/pSA3E
ES2LBkSz9rF32+I80a/0EBa58c+LjFsI0NHPHX2frQQuCYbvAxidkEoZegZOt9A7k0RgEG0HSQqt
QZrGBQ7tWtBjM+lg0kQJvBlpF+ePt7tPs0hqILzcBXRhJ5cWEVSaEEkwVqDPSlwo33n43dUo92uO
+yBEJ/E0pSh6UV3heOxChEZwjb/kcaEQOj1YtnllOR/j+ckgxKPVoW0hjWkXNCODhW28smt6R8lI
v3EzRlS+ytbaxiLTXq8kZyUQEKx7kg6WUoUShDE1DQVkubEdXZfl5gBahrSq6HOL/lhwHten0lDu
NEtrIfjGQIaeOmJPdOex8sBXksUuMH3erNjBvtRR4Ey5qaArA82pI91q//wpfI92KuYOpgIQ9LrS
fpl9GOjNQ+Fl3DEI+WhE0O+bi6V9YYXKsnTXpHGUjytTNJ0UUpgegKrCnUMgtUlJqPgYvMwm2TOB
Na5WWL5l88NzLj4UIrKM3jVCmcvwxdarJ1NV8lsSAsDyKFrP/7wtnuo0rwQA6FQ3Wu8//AI8i1BB
s++mcNQeTw4L9zKPhJxP7+Q9V9GVNGC7wYrVW6cwTPuJKCB95jPl97AMIW2fpECxUhBy6fwUzPnL
cT2NsPj0bPTICRjIxaVjEU936YTt2YNsOftvUgzKlikikyT1xfOAsBx7vn6qjjm32lR3DkOvhb/4
RgEnKKBeklVRvvfHaEr4Dr5I88KuHBKN5ZhO7Xkmc+pj8ZGM4Q/oAaNt69XMI1URFgwhfHdcVWRK
njM8RrL08lAZyoucCCPhETYb7FSz16BeB9OsYaQO9VYbyqC1x1mGdC+TtTgDU2ymbFFBnTjnFLBd
/EZYwWroD7om65Ps3pbyG0zf4/9cCyBfjmwFczB4nsKi8HyY7N9VnFU+mLxGnEhKolPMQmVFSAHh
ytYNCcI1FJ29jrzlaTIJItev27F4i5drvnLqFJgpsx/tZrT2jgrnlUpTBI0qLXudivWbZeo/xbHo
1e6eJIt/E4VQH69hEddNpS42dmsuAygM54nKLB8iT5R0nrrQziuWUPtQU9PI0zl5Jpov5HCM1HCW
Eu7+v20TY9NbYE2/KEhYss91r7C1/ZliCEVXrX3lcJNLAwCM9Kd3rXkGwKtusbFdQxctO7YzoOQg
GbQEC8GSMqrU9cIKx8q3yLzEw+Ad5hvrFb2sCSWMN/VGWVaQpcY+U8Xez8dROw3jvWVEss8Xv0Wp
XVmjLxuHdTrAXLXMF+iz0k9xnwc55IbEPk/ESwCD6R79MP4ndwrMlCvJ6GaddxKzjE4KvHsrhRY0
j0ObFscBilYyfhTI1dFXaRNufRHOI4MkOiiGcC3MqetPeImKvO5APEIXPMbsLfgZuA4+/RM1RLlW
n9rHw0jNeb6M8+uSDiJGvnHvg0VIWqHLJwqW1KBHsS6mW8CR2LQ6B7DS1ld/jb9VidqxT2dpbfuX
NHZ7oDSNHL4tjpafEiupVU0sRl2apSnW+OxVspExK2VZQ9knkamgpJfb4hjPbB7RbO8RoBO0nON1
PoH3mKjmfC7K7QCJUe/KW970CtN2nJPBljxNoYWy8PSHW7P0r25RYGgMmbZqvqfSdgcCbvNcxYfc
kl+wiyj9mMdE7v2tatd5wqAnV3936UloUzIthsPvrkwZc29rkTP4w+xq2TKvYf8Y0Z9wS0gBt5H8
hy+zgnNvp3wnkkVZOz468Rjef+Rt+2l8BqFfJP2lcMId5SdkrG3M8aYG15jy2bLpc6679T6A6NqH
iXb3Q7V5I4jYWdwOo4B4hFBAxFqobWrnpEzYNwbsD5U4IuYMULvzhb/cckDb1gHmddQr0bwqTMul
Fdl5MiPfP0PJIe2MOlLz4CvUmxrYk77E/5hhUvx1hH/16wdPsMNDpl65YhsYfepB3dNAMwcYd1zs
RRDF10oE88yu4zRtHvXf5DTOrwjfCNV+FqfBq/xGYQjFJcEUFPW9Qbj1/De0A+COHxSDTshGAIc4
WcDvPFWr51k76UW/cMFwrZv5g3bTflUS4E74Ukot6ajLpaJKmgU1ECit0VTND/Ube59xe63WfF9w
aIBKD63CoOTHSuAU986GDBzU5KnEYDLR6aGyedFDksnDqE3LrvJDHusDGttRicxiuZMcjh8rz2gq
XdQODIqeDp6YZYfZBF6qsta5dwwOQ5tTLAM7kqT0nirFkzxs9p8ZI0ZgqAobZ8zNq3/+k94I0x/E
r/CNNoyD97SdlsZi052CMqubyCnsddOQ0yOPQn7hucwCs5NxYs+V28D/6unE4NycnreivdVF8G2q
0l4EW47yjNrbLQgphmyzDSMOSdAs6YPf8uh6NvGT9CDKk0oodCehQ7Tn6XzUfvGPJFMvLeScDT0l
qKChTiIKe6YnpalLuDSS9HTyPLUmTlgEMy8KrkQzmlDZYuej0tbdHcjiooA4UlXeyLMII5L2nrDI
ge3AhVJAuxZ/2otmBJVZBinXUBvNiwq3cWNzj5vM5uaK3+O3UV+ePVuUaixZn+KV5+bCsti6esfW
p+DRxYYVylAKvam5Ym+KpD9bNkiS9Yd/NYqM2bwDyS/UbYCagN0WHb6EMl/pYkz5bwOUwdN8/kmW
D/vOuk4QZCCsfaQBA+FKvshd05/rtQktw7JN+OZwO88+/OIsV2/dhtbNU43zjcvLxJ1lw+GzN/7l
eMXISgQzHV27fkZHnq98jM82mLuWQ00kOscaVxFjgRPGjpOJQJ/yIA1+nnyuG4GYJbG0RmREoD/7
akVZAbiVYARzGdKVgtp1Ajy9vYEMxQvDdsu+o7XsAgTGv7oLV4GphlfQAHW2GfVtkGFX6Ie0sE/X
2KOgH9eg7LgCuA0/KH8NdpyzsSpVBV+Q9lTRdOm87AuD4ESYOliYRM5NVjLOkYjYaNFZ3TcxOoa1
DYaZ2bcmRgpvTDL69j0qwi+safqr3L0t3pE4i1cKLW0fWkcde1YAnm+TYMAAXygFVfOmXHrppBcd
AoDkiajvdrtfsyjG4gFJn13oQWKl4nfHnkvJt93SVyYHW2bOHpAncqvSKA5LrbilMiN2k1JvQQZC
TvwjiwLC9+4KNZvMcoscGQSHNo6f2kVuZuhgeIow4I6WeiZogOM+aMktlIF0xCtSJU9taw5unwqF
2BqSHKXhOWqG6qOUH+5Eg5pEY8xNopQL6aYNDF2EEerFT1F+syT9OEXZL/HgAP8NLQsjXu0EX8ri
oYq29KZ0BcxoWWjPm3DxQbcH6LmeJGog9NTjN+OGABjyyXY7J+hK+O2ZRAuoH4ZK03hBs3nyw13S
GvwCmJAgHfrHBUftYmHvWvGXuMb3GcLQsjjHa9wzkniGh85GtjKr1ONpFdl+7AhpMpeW9HKY59Bb
WZS6D+AxmsELsa3t6Ex6bQgb4uuYpVYc4Kd5QhovyZZ1JxQYtEiuNhb3o5dEZKxQ8/0e1F1QrHmc
B0QLeEM9gDArTkYeTAWZzRLSpTobevAegy9Eaqlj39KYsO01ZHsa4kInxw0YeNPYs0BEYqM/YMRw
sx3rXr9Y96U1AmaamfXwCbDCGFzL0yVn4WtrTXvt0NiR0/K21q6ZsVSRXxwdXcYq4H8g7icbkFQj
Az1wsRVxp0j55eM1XFjXrzGA727E1Zn0m7gUQ+uOZsM2Zcw4euvM9uL+7sORgklCZL/tapbAbnsX
cQeB+wgqe1JoWDOC8hhuPNQhLIwaFS38LYs06bWYe5AXtaQ5xjv42Ua/FqBKN7PDAx0mvcPrALTB
SXVsETmf77jfuXntqjpRGfIXZYsXBHD98Me+E1nSWIsbA6v8xphXgfVA04iOXlz1EOnZcKDbwbRw
LznZ2zEGziKwyQMpRlXnY0Y+ZdRhGAan9jl4xltztdSMQmoVORYnEtkp9OmfOSIIyZzbDOrJNlU3
2b1KxaGhBJSX/pTSCA4ukNu7yYmaCTZK3zAwmWCz8XNic/r9oxjIyjHJIf7XDchTjZqwuO+1ypks
qig5UqGRPkraC3EdeR3Qsp8dO1KEadUiJQKYNEzms2xxgeVDUR9XnLbxUiQJoy2bCplvtYh1rYLW
zezt+Wo37l0+Z4k6MY8FwCHkEmV3ikRePkFdwJCr8MmqReEU4wbFEvf7DXOnLOgsqGL+EQsQU18l
Neb7Xb0vyN+e4ZfgSjvoqhrVPHGbyKjk+l6bbakwNCWDy8t0UvTCRvS0OYpjwc9MbszhN9U6yTRS
J8b9k11O/gnBxckW90rIi4IalmKH9gU8p/MD1KnEQ9fiLRuCECX3qFWrjdUg/EIZoWuGH0wnf2Dd
xy1nmKUXHd93fBjWCt0h2klYceeawQar3irpMwR93kAsKOf7FVeAieWVoihk1Py1icfGiUKjMoKn
61OlT/CWMRgHmESWnYcTmaMNAR+4PWOE+tsJHSt/DITJgJEzgOaICUscK8LFzPs9utWvJrYtrNAu
nrXIMj8nGr0p01S4H1IUfQxPEO/CjGPBi5Tdr7HTr2rTEy8ui+JkEUGAayGGf1cGkxmUmLSdu6v0
ZvLzsnysLpm8FRETTx5DazD/KUhLO74VFEQhpyoinTCaLre5/1OQb8KrmOA2fNaaRmgYZHQ0+fF/
jy2/K4EMYwZ6e/7z4mLz18nSS6kaLsrqF7UTx/YgXZ08DzkGwr1LQmka9zXc9K2uuPWrePbg896+
uAkeeyH/55aItq09njVtjBbXQbFmVa1Te+5+CNE3bSg/TLBVJjXiVPK7e0Y6zURVIrmwI4ApwYcp
I5izuqW9I5z6M6P4pamYsl6rvqIV6gvzlaFX/t5ocRHWSVuEo+Ow3qTmNwEJkFC01kPqhkSmlgJb
JjgDHbZw3uckT3WCN6X6rQyf9zWlasLtmFbE9z09adXcteQny75h1p5GW6Sa/55ntFa9HQhe7mzT
fR7EEptvND2AuZDggreaf9bGhngr2k5N+8KwD4QYqsqzoVpY6UPrwRmLkogu0HwlGxnzCn6tkBc3
1MB9PZ5QBtiOQ/Iwa2Obe6slTxksT0mLn40M8lBMVfsOXacwgdN5EHJiYYfUije2wpKIO38BEaHx
mNzIBZ/gp/znDHvC1HUAAmNmZonRrD8ZZ9Er8DqEyigf6n57ROVHDJj2DdavJYpvNJRhGICynWJX
aKKV92uznCrp7KjKZulzBdcnJdFPCEfAxvg3Az9QnSTX6x3k3UH0mzj6rAo86zumAKAbg8Qrpt8g
CzYIw7e4XXCyUzlM+7qjQkIMsiIhTRxutcCphIENO8OkzEL52/8pkVAmeVLnTjXLLs+U+OSmsmC/
lrPsKoY+bg5C3uvSV6PdSb1ZFyeGPMbT47v6Zv92y1aijEMOde9qWTRu24pAsWxXPjEkrLqXK1Ou
ufx6ym5P0j2CxFP2F3uxuuLYi2nAIpQssPnrArKr5sCgKobh0+ovQfQo/qZKJEYJpHuU7GYVOxdo
c9FmUR1+BX9VAo29OFGwUKHBujd2MgIkTEIOyYTS26ItL6Hy3oZnztusJeL9AOyHDwerNa6wtnxW
tIsIldP4qEWeGckLMG3Q6mlfR1ct9BnBpeLkd3w2pm+WX54y84EF6p0CWKE9FsqwBPLoycLq77o+
L3fkiIGd4VybLmXtDCEYTawCjg54kHv/xeFkU/+O43lbqV4H/g9G0E5ju2fUOLrASo+pFYDqMO2D
ezYuyTxXd2Uno6Se0+0Bb6zUpRXpmZfZHu1X1JP0CP98VNUteGPQXJ9PXLwqZQbkdeWT8tGgot6H
kk3DoO+vcClmnQQMM0pqai6FfWsdu17cV2hYO7/YZ6B/HOYBCyJUxWDgMCOPWByQVKpthR2GxyeU
zOdIXJpM73Bxzj9Bn8onRVjKCSSBCboPlFjy2K5kLybQ5CsZ10PEnRcOI7D2Wkix34UB/CAIxXd6
0gaChb/WSLU2uE8Vg0f5k9BQDTTV/tAmif8pzu8XRwavvC5JiusnNz91AqpyJpEEATfxmOuiHVrL
xQ7MfFRkNGXBn1hCDowqMoa2sdifMhGkf1GfudFv+faEhm7RiWf6YQIoYDL10x3ntOlqj2wffc8V
F0WmXcaZNxINIB0AMbiVMzkqmIBWAhsYOGR8DBqlFPeJMiJtRl3iBLYrVZqA2WhLoshf3Q5tfYae
XFyfqsHSLrI9mZzeJ/mbt88H2e4dr7kHO0uGLwEpV9ynTHlN0Xl6J20V9AGwFP6L+mXj6RGIEiUd
upr/8RxTLIYR++VOCtMM4DYf5v3YwoNGdGtJ78JnmnlUOJ1aK6xxSgeMiF0wFG1g6icbfTrbHFdH
8oZ8JXULxNaJvRiq4yuFW50dEOgExtrCrYp9EhL/Xj57xd8WsoTqj4o+eyP9Jrjrluqg8E4W00ez
9GA6b48vLDdJpEDC1Nh03epAk1yu0piI/6ehXLR5RCQ9LUpkgmrHvbAPcD5bu7Iq7uunLYwwZM0c
u02CWbihQ22Bvy3YQKzKhBS5Xg9w2WQJlYtD0rY6YlqjZ1eMfhNf4Lrr+HUJELlp2pN7S5MWpN3S
SXktHWMrGMAOHZpoyST+doWTpyosgX4L21DnKkv8jNka3X5DUad2oQ7FuYZKRqONyMNLbjillLzs
ckXrJ32cBFH9r7RclJ4lyUv1HXXeiSLQzf3HYXr2JtqwZsSXGQ2rx4AuI7phGI4kPX9DWs1V+fi5
IB4dWmtjcPoFimvOANcuUgNnd6TDVaNDbh/ciJnH3uAWczgqURblXXrCpJCabsHk9LiiPZABfv98
o+gW9i4cYXViLabpeAko217nCTNe2OQYEf3WOz70TEtu9pTMD12nFhgB3nAXchvlodQ7jr9S/ocZ
tjpKio3fpnfeCy5s6pTMuQHMplsnQVw3MfIynytre7QNXWQFAZvEt5izs1t+xuRdIka7/a/STuKA
oxmsjpooxGnfn6FyePHnVVI7w0GN7LiQPnfaxbbVf0HHq4dlgH4/PuimsbcBNMS/Muy02xvWm3PM
K72zTFEX0IGXSFH1GxoGe8GRDAOuN1Wwujgh68XiBzpxvC5eP1KajQD3Us+OgflFbc86jmDzhQGI
CFgHgZDr/+NkXR2rIJmMbZJB5b/4nB1a39MsQhmiiFSD8iSXRoJTRP17XMCS76JPVAFDSgX0/OHc
DssDq4VpesW0BxJVkwrqC9Dncqcm6T7/46LTWM2t8TTsiLInoKNhoxyO51XJV+YZgsIGRBfMIqtp
rj18CFYlLT4JtoJrMdog4zkE36a6X5jbG3D6UoIgj/EOUZ/Dryap/4rY6iLrrPiNaojihPGo8te0
1fus12amRysh3dpIINllox8W0YCHNfDI3CNa5d0MAcFSA7zbmQxL5AlfVspMyTrCcTTmwBOlhtoy
nt/HjswiM+xpwz0eN9CfcbuHaHDGpsJQF+OTHblkuZKVfkc1Ahkta20r1YdEvsZdtPWHq9Rx/Qk7
FjZppKJpBK5hJd9VsplLDlgEUdiIaHQb35x43Sg2c+DzKI9u50dbCL78lR/yyyCF2SNA57Opyo1H
vBGFOqXYG61W4BIvT41Mt5PK9hVKM/eq35VNFZ51JtY4IFBUMjB1iwbJ9OA98NF5uRbIHhTH9OGi
3kR3U5HvG5kaNRAhS2JD4Pr/mQsGpVaUazPIbpFUw9lQ8goaZSmlv+UZbmFzSoxPbznrfmGrisA5
ogtn5jw/gvgquWwP3u4x41dvxNZmuXTJjiF7m5FCSh3J8vJh+ZaB/rzn6NadNuSUVOAtJ79vjdy8
Y7WVUmYNDs+Cmf9VbFNRkVLUCwIbZcVqCQ1iQj2+BHE5W9yZs9+VIBIxPkz5672Bm5lnb4gKJjGQ
d6+2ejJhKT+w0erolFdZnRpzjntrIHrCNQb92GyNW3nqDOhgPcC5QsMV7v8GPzWZ7YQUlZDSPHSg
PRnh31SZQ5Z+fdlqyT3X+OfBYosvZpplmPxBwyYDep5qyImI6WPjc4Sdbqxjfj/JBSzacdaK9ybF
hfYXzK1ZmTEJDKiEqJ2qJcWZJUegv4ZKsbzYKZsxGEDjkAPeJtvL1qpa4g4slbXRq6chTh3GEhoH
+3aWfy3EPj7amEPtEYDrb59xH6enoKbp2ni/er/KRCVNJ+QWcrv26U6R9b0LMpKUe9xIL7DPIunx
kh2dh+jhtsP2OWkSBYNmNGUbFL2gZ26OS05SiH8h/N1/Du2ERFgwAZiGAzmMdFvfEiLtKbLEqZNg
DbqD3rQcsdXa/WlO16tVIj3ENoLPGgAtlCeiHitpC3FWbYUlK8UElKzm/XXwWJrU8idWz5Z1ugxj
HTOdXkPWEB/OGd6Vcv6BR57H+obwTDWdYlPF8P1aeF67W7WGciPaUtkPtpHvAMY8bPkn+XOC6U+p
iFHY2fVSwjgBiNGw6GCo0YbObDK5VWNMw8TN0yJ+TywE9/ftvtlQty5mc/IuC5cjJ8CHf3nSVsvB
aYRZ7JRFdhUxPiZxEGvMFgf2PaFDdr77L1g2sW4BrzzPuQnnRblYwNWjhJfMIfUA9CDq3Xb4wr4f
PcItRec1Mizy6RFWLRfy2T9mC8+MJ0NdSZTxx9d6Sy5FP4M8m6ZbtIYXs0RKQCQaVD9Dh6nY3ema
Wy7Qk3A/5VuLxslJvHNbnqzZUN/YcK1pFcLnjKoKCpG+IzHhFBcLvAOsx4L7+103b2wyETXo2dMe
Sj0sB2BsaycgyTSAryClwfoO1yMcABvSN60fIrlu+p16ehFlUgQlHnpJwtlTNW6QjNkAbN5L0Do1
6nC1+kXztfxDF7ubdf48L8qgZLCdO09MbpunKrqCME8S6kpR/fFHqjv2IC88Hv2dBRL2C9e2K+7K
iilpIGIKCXZMkrA0DuEgq4oWRIbCX00owxXjhMu6vcmC9o6CX1O/JQt80UzQIPf2bEbTP1siYIny
pb+l2zAm94mUwOf7GaC4S4E5y/2yiI9696n7JT0Q5oG+NtJeqH32A/u6qeGmCUfKotNskD9DJYr2
RaIUmEIeD6p1n/8bLRoPVGvhbFKGs+CQopHGXbFT185tiKwEEz2quMB8G9XftNbrFlqN+wH4n/bN
+r6P0DR+78cGY37cEH2r1RNs4hezymoEsuDOUHN7hfN2OX5XC20iCibIqZCq45WoZ1XIkIgfnwAg
+h2upSNk4qA6JOErXAAUzaEkEEtybTVxyaiYBCjUGsIP4N49qbgZVffWy1HX/Z49zUtTpIMQhp/6
lRpk+UkSDB6WCOuvTEkmxDfG99nop6eKYFWtLVNk9lyPATy06ExszvsXf5KC3VZ2ICJ31gkXMLog
AJqZhbWz/EQ1VtP0swEleZuFQ0UHuOS63fWJAuqB38mxxfcke7hmj/C42feUuVKrm+0iBx0c5zU7
zorYBcdLfj+J6r9Ae90c8rij84176LpBMMP57wQqBnx27f/9fPvXyCIDcEKav/F3dh0sEgnWNIfD
IXpJl8cuAZqCEvMpFAYZtEOUtlgDanLq7Y2R6fMfIgk0gL43ojkY44PnL2+Hn9xeNp5pvX2TTp0/
ycmytKAXPMf6E5zlU7MOYhA9D4b0TvCmzHKHs7MMc9s92ka4WQGMUzZutVNrX/ug88EdawkrS53U
fJkSjpeWxI2kkMRhepSSvQY+THH/hkbaTEn6x1hQb/1Pm7YsGVNtplVEKtjUsHtQCbyry9IXnMuS
Q80Vl0Eo8qnQo2fMqjUgYUG+pIH5QPR/wS5wK4vpdVlscGUwfUCXsOpUaj7TzCjcFE2aRPYHMxt+
5q3JhfPhNyeK3UtpEJjd6PRqRsuUVDLV/MJyyH0hfhQKFnPx8J3bus5VLAUdx1Vxi2mjRXqRTnkW
o4h4lOulgMCiNPUFvjUzUg+s8OAaFrhAvl6tYto20TP3PqvCSx7OeKjkWAcyqi8KsETvJ3oSx6PQ
Nw4jzm7w6UJJS02nZfJLrZeuQKWLQQk23IgwFSBSQitadqvWItxiO7fTzGURI4vn0Wlv34vOyu/S
/T7hm812CiUTheuxEjDADuPvplCyLnjNAnY3S83H3XMd8J8WhxA6Uq3rEyh6PA3oQw/VulzcA4dm
V9Ghs1tf6pTESmydzjaegDgvRHCqvX8KzYvz1Xbfj0eX3M01KEzxOhA4wAO9CFTqfNgtL7WfUwMR
7AesE3fU+Bz9jmzv3EZ5OF9GEz9nxvz47csPKe1X/BTaI7GML/MBz/iXx4rpv1u14F+tNjKx7tzE
v1oB9uxrK5HWlPTzrXgC2NzD8NbX59JzxMIvZZYKdpovkkRFPt5qiu+y/a7WHolnL25azGAKQBz6
Ur96xgsL2fm2leE/BHHtHEVhvE7X1GnK2F7Udk65mknQn78e/N6LzpDgyNvjopA+PO1z50isSe6Z
gteQYAF83q9qQX8CofNQKzRZzC+EVBd8QUsliUe6Hc9gv22Wjy6aM1gTqtQCBeMKV5gHJwA+SQIn
m3RXc4josYF2zyLQsNRs2f0uswlkWmv2oCAMQ5kPXQ1uIv5KB6DlnXPjwu/0jT/R6oqP1EQvjhN3
dFEPHhQPDOYO0UErN0wfBCsYzAMF2UEFd34JJofetnzg3Kzk83r5Lv5DBMN9+hlFrUX5E+9SyVDX
7qh45AbeQ1iv45W/VQib0SyX0qLRShlCDIAOBAWwpf44tgf/rzhWCHNa0YjK3eaTZJCRm9JuMBRK
nd74s0pqw/1eJmXmjj6Jk/r3kz5nMNpIQmavYh50ewqzL1cVz+aGoINSdG6EgZnm4OjLpyxlhpNr
v1Y/aoB7NEmFfXl2KXoeC02gduliVPkgnDT4sNiit9DHPVdyKkdeE7bpMSp4SEsZ8Z7bmGyVdALA
wRpBQFHXUXJJVZyq5UtLdLP81IhVNZBHfo8NYK0oe32Ps+BrAf8BiBaM1I8KEL6N6jcPkW1H9/xZ
L9m15/gVFCYa4OqobZpSyRH8OOuMR/fIvJrV+KAJ2vCLVOKCf2ePHBAi7CtIQY+BB3sBs6ZFS4z5
SfBgdGrAr4uaHf0S2P6e9U6m5pHCyd241stDZ3etzkg8ArOjEB+/CzpXS4QoraOIPUV4XZga2DZp
hNNZjcttpZR1ag+2C7MsadJCIGTJOhOPSPFzNsUSLCoe7LtZYRisytyNTONrLIo+1jCUrAjOSZ2a
UsqIFfLOcudpavEO7iO+KUp6s9Ro0mJPqdLogwm7uN94f95rwADMoOtuKA/9t1bUEw3yJ+3SNQhi
ck5EBwTcddXX2WiCc1ZJN6IcNa8TocGR1exmX0aFF7UrSkLeoKmVqLW/swPZ9PJ4IvnCGdbbqw25
akyOTpBUrOEVxhcF2BW7H4KH8KkZf4+OfCGLKGJ/sRvm2lBRPof6SQesZSIGckmDge6toqZXsmmm
JBw27Vn414AGdjBCnOYZoOkIzbgc0I6j6sZXm/uyC/o9NwnUiePbCR7w/qASjZgbojIKYW3pR1zJ
A0OVo71nR+/cpW9ByewNP9Fp4h0MVsVC1FGZ8AJCLSS87AKI/ot1dn8gAzNTmaCkXCLjQlE/cv6K
Nev6pobcGd5PmrxsZDVwaUIcf9kuqsRAviJwXBVI7qxdXje1oJ87srtROJwwpxvpc79kAnIJTXkH
qoaMIq6RL48Gvzla1V7WqSjRkJ4FW70B6Zr32eWAaYAmB6fGNsbMDqti5euO2hcvAupfAVf0BODu
MrufxAyWEO7RMQ/yn+/H/UN1hm5cCstA/rPrNVKqGLKoelexDnwyPSjxfst5w7W9CKm+Det6V7Ax
LvIaVNNhC3DN+N+giEs0uSZQcWqDJkPMDCgMp2S82xurgkSFNfkXhfUPhhNZqH/XqqRitDLYjf5n
rljFhaEg0MrfmRj02qC80bQBS8N8f31wgmdc7inSSFhWqKuyooK/EP1T9jgsELt5i/ZGwiJpZ1QO
sPm4tg8yr7NkiltZkftWtrvsGiJBPkHSkoL6t7TuVf+/NjFA9ViYwRSi7g6qWFPaPxiyJH5euMPs
qK6THMzR5MXGKJkR3ekpvgxiFZhmDaNBE4NbngaDpaSoy7zj/r4leXHTjetNtpMSkrpoE/rQhkzr
S0bBBESMmHB/amsEmIepMZKvZAdieU0CfONSqLSTB1zovln+Hk8geqd5ZvTbijq8bET2dhok+cHX
prBOVe7hdd4bx3bPqh4dj+W4lbokLKb+/SGfaHGP0z2eRHL2jR+eL8P99KuIwOoDojpcPBs2GGmk
OYqwa8CSc0iS+LxAgVqONNW0fxo48hJ5FsRH26WWt62hp6p0UD9B7TWMosHzeRb8Y88SCac+xi7H
VQqk7Q44/EOWk3H3TMyex03WfpQ9zfzwX615JcyfEAUDh+ypnmWMjyLdIQcWMyKcBBtwQPTD8Ynd
iZgdD0uIz3UJauwQIJQtjgvZsq3XmmIVpuQfWQuG+Q7vhMddZ1/Z1amyFd9gbwCn4KzdkCzc/ZFj
G1Y9SCJAXYoImnmAczglISJDn/taIRr3DMPPBlp+p9dUw82SK8JSNDZuwfsw7oCmYgzTpjuusFvi
B9nKRhZtQTULpg8UANYNAErGq8jWv1c8c9SwqnwRe6AmUcTh5IgTBl9In0Q/S1iIgzE5sCRshvJo
75EtumAMDTumLp4maJIIp7trUsbnuDc/pC3jyRnucQdc3nFuFW5m90pfZQ/lOlRNXMzB/ti+9DaS
h3DbAt03ljlkZbXPkDVCwkAAb1OTrWM3Y3u9lvH7QUALEdonj4XqPVxBJCCWdj4S6OL0E98ZptNB
odAcamDIYS4EhGnU3X0zll17f0rUAhh/k0Cp5mQuDc/3KHWR+Up2aHG0+R29Ly5djrWZY9zxODi+
zK8qHJ0/4MJncpv+3SHACb0rZ1YdKl23LAsp4GMTwIpLWYpdt766WqdiMVAODZBqIGg2hKhsWNxF
ATesQcz/pLS/BfvSwAy4wJPf0vPGbJ/ohiqW+45yPOaGiR8THjHWAQobyg0Quxqta3ay2yhOaYAa
c9y4WdvvSl9R9EXzPuhq/FROY3mjQC1dYSdX/Z691F7xZb1i67F24IsyzDdoMyDjtJOqizwuyX9R
zlvSrOPG1iebdHPBm5TB+p/dW5eJuTWuAwdUA+vux+uImFtLkO1RnJZzXRdAqpEMFLa+Ouy4aW3W
chK0Co1BZtVWwfu4M5jmFedEvLnwRh92HUcPuzAkblvQ98YiBsET9pBvjUWZ7x3WJkeK2YCrQdBP
VHSP0dmip5RRFEhnRyRilWqse6Afe9zw9VqE16TxwCMHdJMnCu4L+BLzX6jkyCLHosSn/Isgghe4
zOt0wG2v62VERRUWrkK+4Yy1rprKQs+VTSv7zxpqSm9vCKtJDHcJGcG3i3oQ0lmvSSLHt3zpgl27
XYk7/W0gpEz56ZQr8BXRhi7QiMPFjPHtjVvfxCzc2/n+vIVTdz5RQbX6GakXcD2D4YruDpVG2Ke3
esABqgF39Ng3wEn2XR9gtkqozGKbvvrOoBZVbfvC+hHtPHah2BJUuGHoJK/j02kfVdA+W6Kb5jXU
M+l55H+XFFWZwCon5WI2TORrHiF4lxZFfIV6XRZvGjp2kJmYlYWeXGuJFG9TX9PoQBr3NETMTvEo
sKZEBJWvdZoPTurd9t9xEvkoHZ7ilMupMCUn3+hutsdkWhs4ZKI6pKxYtL9Naz9HD2YJuzMSugyW
Tsd2xCmVVccOPLPxmZPBpcXor6NDg+V2HjEDUpsus/jL/0ybC6beI9sViWLC3PFVPH1TqN1e1Hpf
UACiGsz2BTlbdLwoF9s7KJqhIHiB1wnEP3qhf6SZEGnsxd8b4+oFt4IykGCcHke9zzpwmv4c14Pq
zSiG0/x17MpfrSVS6bhR1xVh+vWr1QM0ZVZqv451m5R/z/HVU9GLi3jriITrm0Omv+XsyDQUl0lP
aLXQjnlgpWHIwapxvcXYfdWGS8hBcUi26/pV49HM7X5Y56DF9EmAzdj9VRa6dTkVZMQJlwPmO+HV
qrDGCyOUPr8VBxkNnzDnxaGPi3PQLBOupcq/Ls7PXbtlqOfp/Fw9MXnSAGcc0Ajdm732goSktQf6
JF5+gT4GlwOFNZ93D2p0ffH5PvUlU1B5Gs8Dytdyvmrtte7NDft6e6vh+DVj7IAFxQLjSKb/CkU+
IAAitC+PR08UJwH8Cl+O5gIXB3hwIHpvoepi12rdvoDLtXsxMOOEsbngFQZiwej44QnlN7WiLqaJ
xTkCd+LpO+WgFPKvLyV3WWjSpIU22QorX+A2DhXp3poU7zWyd5DOa0uz+BUPBLCOKjBM+7sjq78L
uIp5qFtEFzTrWE6uy+3IN/F6ljATnYIEWzbJT9UU5Ti9Ft2AaUes7eBX+m2MYO0Finhqt/U9rsJ+
yncKAD8iFI09aKDcLT2W9yTmtxuZsV+T3kn8IDT0rUq4WnnDZVhTPlkGCUQq4HOllYufWh0HBIkg
Zfb2iBgf008qJKwmfEZgycT7er91/czgj+49O7xvQKLXoyajK3DuSVki/6XeYvntD35G8vc+o+My
6jsuAg8WCywYsQYnY/pBPPPdxkrETLDDHZ1fqPsVYMqEVf9GJQPHB3gpth0SWo3NQD85xPknyOQK
oAmcQesvi1RYdl4li9CBi2O+FwbL/o+dl5t8FusC3N9EGZSUDHGAkGmdbSIVUKcP8gTx2nc9e77f
D0y8f9q6QIQj15K5H+eGBbU6eBO543v/pdKWJo8txkzo1pRVMD+/JEn1sEds6Z5Lk5BpniAeNIHn
3J9ubhGOqlANArS/33VNlWNPdHoMBxzhMqY0zo8f4Y7GzuAecUBOhosHzFYUB44enldcFkbHYeDs
IeiaNfAO7/YC4bJ9BBIsSOdfvEohfb54VbQRDiPjVdZVzGymB1qSc92GJ3daE/tmlVpi+mRt79XG
ug1AmDbc75iYd/Ev5uX79K1ngDOMY3cPatObJlwHRqCry1AHzibZgUReXOc92R19dWNeBvLDsaQU
OBzGu1kIamKRIfkse1+FXSauVRy1fQc47ZiaGgtggWpzXif9izv6UXSaqG6bE8l1DD9N6J0NCH3a
uSV8TQImcWkvh4mmsIBnOwKacvrz5g4LHfBYtOWbryfH+WPcsNYvQ7i7rQQOQngvaQMLpzcgqUzU
4tIQTLU002oBQZzMOJDNWUM+hvPGumgA/arPjXAjd1Cod5L/CFEUQNo0X8Ntx6ON7ht9zoVPXBh7
rqv5fgJcDERspPHBInFNmdTsq3es3gURXwvrjcEeJT2fCpUdo9xoRWbzUVsTfTJgOcvyVL2E51wx
m5d6QCDI06TM7kpKNYtKjzRKtOpIFlfJNHLMzn5CfXS4FypLd0WKxAHqXciDAcXk2nsTz6onp/f4
e9Y4SvPYMRsngoQBpuKT52Z4oW4m8rBCvCvDUv/XAo0pjEkqVDktDqjb6WZCX7sBTJw8E+pIeha3
00Nxewb7vNe5TdBDRv7jLA61pLrC1Mk+cbMdVLQM1cxj3AbvahpXF9dPsrHNg9TJntLC1RerQa6C
GwZFUIcqxJIyl2VvF/8QkkqOuGusQWft4nkE7e9E4ySaO36F1ZR7qOKYCsXcA3uG52aRFBh7jY48
iD905ptrm7eN0Srbfm0XHEyquyS/4oFh4Eg6uvVc4fnYo7wM2M1CD9m6THk7xFGwIoFMRcrzgrgK
5hItp1BGxAs/0JM6K9docJWJ4Uw64CrT8gLGSEgQfYIS6KP0wibzaW3aWXZa7nf3CSNSBQ5N3O8O
Ca+HidsU4PosPoMbpSGef1cRP3d1MuUKSuuzIf8aeBr/nBvkNcuCpT1lRrZmj6U82CbzbIuhnztc
GYWnraG2ZuutnVR8hMDHq2bqpHqGqdpYpNmUZBWjYgGztZTJsBwgYJBhqQQUztYJIhmUwqJOIXLK
zOE7dM3dOsZsAALGKfEAPxVaFPZqJpZjZMvEhaESUM2usrxmmKo+30DRzOilGF4ZIcC7AY7MbqfT
+6SMP3Qis40lC+56WhLP6zl37uxuCpuw+5rYDrFEVMRX7KuySNt3oG9sWlopQiM2x1ZLycPz8WCi
2UdtGtr6raR12INWLMfcgEaly5FrZVRkNtuRqJa0M3p2UdciZqRyWjLpx75bhQ4kCuR2AeK2Scjc
CJ/o9/31kvXDmnFysTmDy8p310b6rtXPdcMl0ivPCWOad/D4/rInHkZsznniWFmj7MQIgRf5ZuIr
udYoxC8FBrpSWIj0vL774NCt0D2mjZKZ72V2nUllnkQUcxoUDDhA78VE1t1XD08r6HeTPARQzLwI
xbOdCmVSpc4atZF3R7u73IiHdd8sSpon9HWEVuyF6x5qNlqrCNywDDHp7ZmK5MuPWZnMqJYPj5Oy
PpG8Puh5qX9fatmJ+qoRZ16fNhsxUlC0OKWyiHDKARn93uxVYhTZebyC0X5aeNazzFALaTavaFsH
vS6Tq4xoxOwJRIlgpZvow3hTbjHKpBgNQ4CQPA6HFHb7u2O68U1XEY3i1sWNzYIP/u2bJIvg25l7
LQh9w6oBDp+7voniW+uzDTyJXDnTCDqNl6NCv0woiQt/0iecMgjOVY2HARmC5Ypgtmek1WUQD3VQ
ZDtxi2/IER9qU1RyK2mRI0OXAujA7KZXRfgxY/3Ui/Rd6IH1wU2dpSDdRHviRpjz0mypNMRe1M7d
/O1wzx9+2QafpU9TFxkk1XfOVXyqJ665SE9niQw67IcJDebZ2DsgcmrcOdzjrMLybwo+qlGK5MRo
86pS5s7JKm0A7t2WkVtkdCVgwZhvXKExh1z+XIZZJc+uzbueAcuU+X6QJicDpNS18zy7Mv6xixpB
eFNEqo0Q3ZlYFOUN3LJsD+YcJuHxyy76f4DZa7sNhlLTnoPwXKrkPxeqG80VJVBUyadHxQnJ7ImB
3xDCrTa0tiXrkLF7mgNMcrsnGSRaUuZr9ra7Uprp3hiue6afc0ATACQ04rZAf0IWOSKr2LoLDM3n
1O0t2sx9+g96TZI1UKFcRmtjC/sAk4uIdI/njdEWAZAx6fC115d/X6nIUqNsu7jkuJUqAKWWtkPW
10j48oxsny+9/6/m4dvHrL0IUnSztA2B/KzQz2I53qTibv/T6ab2M4+r1q8/Yru+5EyhtdP+nQOl
/LLdAVrafVPZA6a8KBGysV6XBYAMGU46QLFN5q1URV1Cq/6GPqy3+TxRaP4JZwqiHORri27eraw4
iXXv+QpHvYi3h3UKwSCS8J7IZsC4UeRxK+/WGHGeFHPWiavfZI3L+w5KJeWHKj56orEeef35ZlkO
IUqZBC82OIrJEEhuIaH7TF9XaU4sfGFb0+vTumo6m3lsn0yFVS6VVgB6efh4rGqaEjPpU+pjdXAO
TT71F64AKTwCB+1tISkCNMsweFb450IY7TgXwhHhdZ/3qV5KW0Zf5AKnZ+5dpld+ku0wmE7ZsqHP
Frx/FPNmBHSqyP4QkpInpMFG3ibIpsWciW0n4E/PcUbp9Lq9lYzYFTIT43fnXSb3jg0S3DzQpt2f
OVTDmhkcIqhtRFBLhW1nLX9A5psDcZYh/zwfbBu15jEJSzmCeaJX4mDTL/OyOWy4rvgtJWeM0PSl
M3M2pfeVa+VCNbmMPHOemPQrfV6LdpGl7feVO0mJtsz6bnAq6tT7f2wiL38n+5/9/2yh7v2oeD4g
3v+mWLM0zpMm7te3nVpSHBYeFVJd47C5s/zB76WotN2aeA9LcHuEj+8LDUOHJKejew0/cqxmi/g+
X/UKiyKokEYkm6I6D4U5ORt8Px9GiFig+DVfeJ+/7s7zaZGXILo8pZKRUmfLRYgXG6I2NnjpRwT+
RDkNKAFYjp8nCmYIxJJ62dgcTFg9meWvSzGh7W44/GWryVVZrtACP3tDCT/3MUe65NETF6CB6Giy
Q2g9octOwgl/KUiP94e3KmYTCX8A1vcZz7WP66X/HK72DWz9DRFm1NetrjNddQYXqK7ziwrsXHSi
Xs+CU1TdM6/4rYDkU6geB621v3371E0UMUBYCttv3KaweylFz03W2Ub6HtteYcwlOM9OjyN4BRL3
FI9U4qtrfWwsKsc2CM6LxrLJoyKY1I+RFrBs5ESyyKasdXstMu5yQRbI+5XixXM3QkE2n4rAVyyJ
JkDImtGVm/vZTJzdsSD21stv0RjlVhbHrYe9mtI98aeOalbUND9Yif4xJaesiF1ltwCk8USglU/i
YRZ85PwkA2aXrEs1nLSjKp0EP1ugqtrMmBBmbL3UI6hkxjBW0arw4gsU7otNbcH7lKa76Rg9IfmS
uMU7JqLbC0D7rRbPJHLdNd+cPXbAyuK6I0iJsWKOCzNX19L+1YrPlXrI+lQR/VoRkmeUn2lXOXN3
pZBQgMPBlwxGzSbEk79jqooiaQnAz33lZk65ZA6FC4xD9oaEWJ23IhJuiUo9SKDCa0nmKx9JbA04
JeWdUsUWo4gRKs8omTqzxY/Il1BGuGNDeUPdBzb4k281pvS84XyxXc8oKqtM0wB7iSc6uXUuPC15
OXoi4WWCsZSMtYavtnpvGM2r+JS/nSCE0I+Nm1ghuMmqajP5RMdBk5iu5arWoRVbnj2xEJQ1hV/P
VHQgQKhpaRaawMLp+ZibavhI4P3vOz+VaW6oUoAOjSKkjP0zLTTfBokl9r6hPoj2Tld2LNqAWfeO
oYfBkblVIwb+T2ABBXi4E2hGeUXKydBIWK4Y8Gg9oiR4eDgGUF39o/WJMu2dl+RS+IeUdk5euiOg
dNZ9vycFlu77c0R9+nDIs1pJCuiccjyUwTORaaLwhMp9CcNoEuJXKg0TX4n0xoty61HxOur++XND
0XXhkNMj98uQPV/uR/sStnORuMhTs/UvohKk9rLJVYgiJQ9LQXZEGCGOoOsWdiJ3PY1cO1Zqb6n6
Rz5X8rfsNE1QGC14v5JU5HkA7jQR6pKU0UwOc5XKWLmMuOdaAm2FyGZqtxmO8BftJ+tPhFz44e/o
fTi49tCWhyaYF7SctbjGfmCG6wdw7fgW3tTbSKomq2b+unmFe+crZKF4EuFu2uDxwVwX3s+QDX9Z
nxLekgsLhmIr5M8eW69a+4i8kotzpi2ftr7jT/qdl66PPnsLIGt5Tp4cyq/cNjS3Jepo4Fxms5o+
9+PpdjuLhWhNCUlhFDL1npzI3ZfVmHWZBtvbhHWCWxttms+3NnrMBVop2z7pyTTr5Ldd2gSfFmNZ
A6fQlt1P4xpUe0bgpo8BO5pkVYiiNyrnMjxrgA4cA8qhc9gocZjsNClA+8MVviYQVqdSGPSFN/2P
9fqh9sbHkj1A/YxUHVnTgGKXVw9n028Sbfwf7wjZ9eI3iFni+M0+izUt7RmKMMpyh4uVhNvAJKmx
gpz7mUBTROCnWIfLZP7QmZLSHBzUSqBXhwRdrV8Uf4c01ApGG6qzMWb2bAThAF2UUQOCR94ch/CP
RFCyz36QFsCfGhLuevJOXdkONjAzbDlciC15zmU+Mqhsgu70F5SwVucDx5rmGm9XSf6/qwdDURhj
ZNDq9oLFawGz99SvA37fYtn3xnPCCA7fGKIOqEFWQAb99u15UzDzMyGNB7QEKekehjnzsW+q6uSF
kK50HoYV1XuYNYRNDJDYxrYqEvmc3j9o1NvMbjAbZm81dLXStByhjvdHxhEFKlCklevNpEBkjXd1
7+XmOWnMsSeWSeCIKOqeUbD5776q6h3Th9xh2t7h2nR444mX17bygETjb8dKEES4pO5c3h39d8yE
Jjfb+fHobX64Qy4mbXqPCD1yMY7GcxRbdZDJKOz9lfRUpR2wDqqRy9yZ4+8Fbul3poPXUlP5dgCh
WPyZ+mC6e3RVDIKC6AuWf8QbFQcFhazu0dq3FbgouaWmvjcWd+42AiFkPoFRaNrlLvXFia7/B4e0
iWAkuVq5UP30OqOs6fISJ6vxwu2S0zfO3E+9c0kF0mibDFEParMZdgSJFZVr/Wt/R5DFf2ALq18G
rWeukcS4pTZ5sxk0k2OtLRztbrndVLsl92dbuoYG9Sh5L3LktU/wxvB6FeZOxbvKHKJarXkAzrUm
g6G+7+FEYwxrSSFHBW39ut5IZHPB6jQGhYbS76LYQubpjeI9MX2KoswLCJvUxrSKTsS1w9hEsXEU
Ubqgb2OY1CTLoYdaEWuwIXMyzr5Hpq7tYoPthyVgZQylGteZZUDaIJR4Bq1WDr7f+/4HLKLeR0ik
TXn3e8pD8Kc3efVKZp/NbH7HU7aXPZHlM92TMre5ahRyJyOraDAYt51RR9sy6n0xHX8+BKyZFoC1
L0I2LRxtaoS4MKFEoPHiqu+usAQsmf7d2g1E5Nl0ap4J2l4G7maK0rBAXauEysSb+TIPuWFflXii
qx2/bay1lJBhUmMygfxjqcFoxBeJiDatN5kPNKyNZUFMkNLrGac/qdsT+qj+FcBYbdSHPt2DRyux
1L4yQ9CoZBhKxcygreOkh9Nrb4fxrxQVXj1JNCawNeuExpoqB3rhsdhInB0Th+yp2o/Npw3VTHJT
UEzf8NNknLNEOlNh5KoATR1hloySsx59ctZAU6M4KwqM4O0VzPTlYdvPY3J6MeR6difTCPzfdrEI
WDPthwqyD2MgO/BMSzviPdC/5gaBZ0OvM7XLML2tIN/d6MWUVcK3nx+F8UpCTlWOp1mfhGLLyZwK
rPNi25Dj9GxcYJh58UADuqKALxI0NHTL8iO0sabx/d0dVk8amq9LmdKtaZCd0lfHI1OaA6MMvS7X
8TQfcBZv30SckvOsAmkRLlMtsO0NwmiOW6F1b3jszrYC8ALN3Ziv24+Z6LwaIji6fGhkKkTjL4m9
hoRo2cmiLGDzbDotVj9YgjCn//SaJbFg7dCyTU83YiMBVPxxFkLRBotw3T842OWOk+uygoU/ue1T
TpuKZzi6dnS8336iq+iELPDot3O1pW93Gtlj/d/bn+M7tiTowMH1a6bT6qhW4aZXHv8IGU8CdhYU
a9rEWsdym+JJKI0Wxjw2qch522nRbPOCwjg6xdG8/QzaTgShzsZ/a9YBD7zQumncT7ApJlWlmTDD
VGgAqvkQnC0hnTYr330NuLvzHsoFZ/c6IzouiyagTTKT/kZ5Mwgn1D7OfpaYNfdJpkfwfkxfxoen
yZp0C8ojX4JlwZ9olBhxIKsc0Vxq1ca/fFw0V5D/BRQVXgvqUFfEposo7/zj8RiEsvhIh3lKdvGu
hTrL6ow6BNOpq5993pkMcQ9odP0+PrFDXS+PRhbyOPYWX0XSHGnSh9eyiDmeotCeOGhPfFnGTfl9
XQeYMHP6OERkgUCn/PsSe7jGgraLHaV4mjd8DVC5mfw4pTMIWF/K0pqE3NuEsH9kzPxI0eEb7D1C
hlkuZCYhh9ax3df6zKVv8gS9nA/uojbij+cnwCJKajxq2viXd7bEVNEDfpDvXVaEsmX/YxV3uaea
2XZbvkJsNBw00aJt/DhuEW/pVeQ4YzJv83Ct7XeNVXWXeNn0L3wdBFD4NKlV2BVWEmT6NSiuae39
/OxtQy6tESRTWDMst8mx3lLzDPCT2az1xqta9Hb2WCvP0bgusv+F2ffHxs7WmHjJKe5a/CZMLh0m
08OTwjGhNsdU1Lf8wS6FjYEtXuDk3kPwLpXtORJl4nlaLyzp1dhQ5+hRbjsQKQUb5BJj0lGyxykY
XJM1Zid10MGJAuxCV+uKh6fX5OpGuo6d22eeqtGvihCA/BfyDv4Qk3tpCvEE0WMBhzBIyu191caR
C8shDKHtvGPmHqvNvrkcRLBgt+BaLiJ61QvZUKPMqmhVsH450nKJHX4zmG44jS8+DboKHt8l0Aik
85YdCvAFU/kYIXYYA/Ir1wK7bIB2qz5mn2bExmCpc3cAdsshZkMn1By65rHJ1jIuGdaYFbwzlObu
zaIdceW/XD5vhO8qv8fTROk+IlmDRh5o/jNEIRJRC7qUD1F2APSLXLjvsWo08flHMEXImLyYl5is
CoExIg816XtuLiTQ2OlyqCWfo6vcwYHwEAPO3Z90wFM7y43DmIgi657mhVSwnVmn9KyB5biBtBPC
bFMx/6eYj1lzbm7IisvDB7tVj4g19ZaTAo9bwOEHAPWt0LZwf1ZaRLILv/PTNsmcgQoCTZPNLn08
vgsVYNVkoAXePNhToCz9QlRO1vwfvoRmAi1ApDdFb+7WZROffKrXp+c0CEGM+MfOIBMiKHemECc7
Pj6/umbnJ7H4mHL3QhqU1eVDrOUMvgdk5jTgmfWYXxBO5OlVKdWztVvVLFscc+BFYL8G1bYY3k7Y
9ZE8L7M3dFxBB04jsUTqtZ+kxZY7Nr9Sv/soXTVeu0hzm8nNAE2JtRJBPkACQ5IuHej97G+b0nUR
hJQKivfUd4SSSDqNss9/F4qrafPYRmygjvNVcAcK4pLBNXYAff83AT+7g0H6d4wneqi4/R5KpO3i
5QKir1ZsEC8eUAfWU2Aw84jEqY78uscEbDBRczORvT+41ECED7KHHDpY5OU9AgBoRiW29kXh+wNL
dKTvp2Woky2NeNktmCiJdrgqi17zJMXy0DJHYsQf24SH1Ho6GpoC+/zKWU86jbkFPaWaEeLWDm4Z
4zQfrotk1n8IeCCivUTChcJ+YEh2GX/dTdkT0uDkDlsleznlsi+YFnJUZmZw926scxP9zUuCCFec
0eSawXIrPKQ7JzJrcIKaitT1r05wJE+023uUre3zZSd9Yb1tggSBoNTy+/oxYF2JzOKh1KFfNbdr
gVHf/s9TJVnFY3dDhbSEJxKu6BCUWwpFEP7B+FHHE2ZZo0Ng+akMKR5hPslnmUJ05Qokd9uWSd9h
gvScONolSPcaPLPQMIrXQMnb3vBo/I0Hwa4D9+uiQU7oisL7Bdc5JkuoiFgUmtSi5GWoOuBCcGjn
/2xwuLewscov2PMdmYDs5D9cdJaqp5PD66sqHQpGp4KUZqoBehxbfBhqgE0wRzZywBRtb5sq3JXo
nS03dr/0fNVNxXBIKKa1PPtjY8acLbfxXBx1mXewdwW/G81IGhfCq6JEq7adDY3i9UXVsJaXBulA
zJVz6b8lYp9QOOh7cybuyC8427KoK8zk4RjgchUiwHMlhLH660oonPC9uKNHf2QWFkzADp/Ho/b+
R3aldji0t5vT9WpFMvnLIGV2BsJV/+92kE9b+0DxLZhf5YaHYtCsvMHyXSmVWx5tKUQIbTXBCuwW
R/OI4fnZcgI5fa6+pSTXrqL4N+4eAApB43nurTDGx88UTHV/lQpZJPjHDpFXNLcBcTWffXyJsBTl
AYx0xiUl7fMS9S8ApuS+rwFlrm+i4czS4Ze8HjDyesH88iDfK+1XHiRMvJDUJ7RSKLJmZ2hFybZb
pD4eJo2lWNq22Vqb5J55+zBmTtmBz6sEXrpiIpNwl67wofefSOhs1GCXAFIyDkiWzOqhzwcDEwaN
5Cq7jNQ3dm8cKZw3ArfD2mzXtvODOjhnRw7BHxY7Q76vwLXFpNm+G1db34qf2WrtopqNdMc0aJxV
lrkz0ZrHFKYkv6mryrOVt/k2HHGm2SY2wIHAnr8aP4Q7ewc0+ysN3j+t9HBCwhNtmnLpoW4KmewF
cl7iJWwpUp3nPb1r/JKEs7lOqYjdW5J422+onXbdnqdey1oyzBdijuE7ydcHbR5oX/Y9DnRT0hgZ
MmypEn9BJQpYHDtPxbxK8ij2Whv9E53QLTB8Rn3JtGF14Q9zhyjU4BLN+MSuRboVZomnjWp4qCpo
9FihDdNzNShNkDvc+Rrj50b6wfQviE1P9cMh8Dyaamh1jV3kfVyP/RXxc0whrSY+m0/uTY3/iNvi
MeoW+ldCD+NgThpnPDtDd6mDCllC68kiErT5qlGeBhhTcJ9kpvO/VoNYTPmfw3y/INNm6da35rSm
Pt/Ckprk7DfDHwiAzaWLRhYzMO1Lhmuw6EvviOP+rAh/bEo1eUZNgeqbIhav0+F2vzJWyz1Leici
l4w9xDKFB6DRpwjWC7Fk3FCV1+3j12mJJZDxjSwPW3O4EXZa1IaIU1RFJ1s+e+Qneho5Yg6ZSMrr
owE9/af590jjYIKtdMPy9b6y9AxozzQbO2i0lYRPcbiD0SHKR5OCyCLeXUAHl8o8shzY5vzMLdvz
q34QIkmnJPkD+jaQqoNZHamshe5LTUoJLN4M4Aym0pWs5CF5HqrKnL85t/1oA8qzISKTx/PScMcP
XLr1yb3Ll7R5mKAJ+6THPdz/FF9GzXBFXCOIVOvbzGkbLU6PqStpme3Qu1UUFl/K67ZAfUKSgdoi
WYX7RpuMuNw82kJiQpUz69bUPDiHMcD5Rx291kx8HE7D1jxPSNGkIhij4g8bDQHIo27JdDVTCoHB
0137w+U08yEc+JWhW5LBb+LMdER+kJ9pAFStxXtKVVF04rpN+41UmfIxLVrEN7CLzoHhXZiS41fQ
LgD0LvrQznRJts+DxBKoZrO+c96lzwACuFuC1NP1f/eG3r3mBXL4kbYOS4OS7WCcU/AO71RxhjwN
DepuLumBLm4nr0nisSx6QwqGSzPIpqGYbZAX5A25pVabar6teO6KvZ5PwrHVEpAwPHf9VIT6D3D1
TPUhQ+3iK6FP2Hu/6CvhEzlqydck8fhBl9L8uPqXl6zygrUMmMNQYb0Yt1E35wE2BKCT4bWT01ck
P03D7smiNnDzWQOqWqEBhxpVu2hhrgBNpuTqdIHd96In+ACp2iUyTMvcOMuxoD+t85Dc17Fr5tYS
AMLcjlHv0cpFdryeCJO0HEAabKe0fcp7WZR60/qnyQlzUmT9cNvsPRRNr02LV+F9gZwltof+AhPO
V1iuLvoujfXi4o8cSNIXSYiHuYdqe7Cc0MInOIhP1PTj7qHh0XQpbpkqKdJPV+VZFeoGvzfTIc9Z
+brT9uNtNhyka93Hl/0qpruLyjM3OA+ZcPSXqcX0cTHBnp1tlnnCHirmpZKSOcO0lI8Ohaaa5rvM
jhTn5zZ/3uLqjfnDL2wXr0y4w+gVe0VX7078i+XioYhMjCai+KiLIXhh2D1m6krKomRYQgwoauUC
W9xiZJVmAwDW8ow9EfJ66yk/kauVSQppPCUeUn6++YfozqcppHODrOe4a4Sd2lJcH26irbBVTWvr
sDn1UrSqDNHgp+1Skt7a6i7lam8Y45gkbg3TvZFaSoO9/WgQoRUwqiGrMcPJUz5GkeQXfc4L5TxY
sSvhI3NNfIQfId6nSLKS1uBc1B9HdkdmJZk0RekZdzNUt6boVGUo8NOU1jivxkKk6qzdsqY++nih
Y6KRhL20akwoR+u2B2tVqeZKElIrc7TXTtjIHSTIzmqvLupAOp7sFJoxmuURI7JVamiQVPbdZePn
g+3JjFRFJbENZec90uj3WTA+07YAO7Kw/l/I1dtWzo2wwA+e/Z7dAdKJuUWoDelpsCTXUDTTb8Wj
POOea6YYMI8EQ5bi4eeKNxTqtyh6I8lynjQLh30nCXQT1PsyTBvTY5Rg6kDrdiT6SpwvjS2HgR40
aTxl5bSwXj+ekGSXiql69vIjYidcqhhoCjUZh9jHUcGUQ0Jhq+fklS5k087k5zdr2aNBnGhNjgeM
ygbjdcsmBAoW6795FMqDCeTMa/m/mvu4rnfYXkmTrBxIIzX7zBuLeDyo61v5SEXRscd+3U99IFJj
nPv12KejYtxixdukNu0pcYaENk4R2DLOU4f/KWEmwVuyrwuTeARbZhUWs2gs+X1K1J0kD2nw7Xlr
zUX5Gqdrf32MBOsuhmaM9MPMIkNBIS52GdxXyY/PF1CF8/K6RFua2xw9giqbh7JqrhplMLuWxWuI
RM945hAhcJ6ltT4b31idfBhwWMTrsk0ZJ+oFEUIPWSlEaen5jw4JOAZGbYKP3sxYSmjTL7eRPwOz
miDTE6FsE/fv1vmqW8/2On3wy5CD3m702B4tA42o4ewx5oK9Q7uPXLJYwsz14l+N3IpcaxBxbh+j
LX2bNDDzXuhubEXpL7L0D5P5ZnxVY1WyVzj61YcOgIKxhH5D6Y9CqLUXmq8AY8TyOT/I2AeQJfyj
SgqgEFEGUgRK+gCUznzRDtFWoHb7tun0Cn5SGp4XllMFEG9bGLKFdhC1MWFo6uWjFxRcrS2MaCi2
LU22AmWDjFJ/Vt0o/dtMhA+lndKtKe52g0DkFfS62+lyT0EAUoafzQSdkH2mmf0nxnx3ASwxj8Bb
IlM9mxXMDuFsYevkLUBHSXPKOZ+c4l6L9Jj/vhCnqY3QJqF8QKmwvcJuG8j+e1NLbC9Bdjalsucz
Im8dfBi2BBMJ7ZmGbiScAxi+acvBlAMsSG6MqeQwbI2FUsk3FKhERLFu3Ud+ovmxgDjsW5EyQGAs
8qDq4YdzEJKVtLe7wc/Se8j5jstsiiPVFkEQoZeiRRx82M+6bjzI6cbf4JqdY/j9Y7vntUcF3wx7
A8X7z5j6/pji8gyhWNuURFHrA+c+bwUKERMA/b0xnUyCeeB9APcop23Fy9k5VJLALEquSj+tT1jN
0g/BRwjpCml0yAraM9lUoZ5CPobXF7x7Mq743l0lW80dKWwQmECU+tuyvqSKb9D41mle43R9DV1J
TTVTu7Ag4LofwF5E7aBeb0KfuTd8/PtMmKoOThtF2Z8Pa9ma2Eyst9TynqKfWx3wnVSWlvK5nWAN
vg5ECewWiy/E6f55Rb9tkOBoItxW00F5TCcbX9c/fRtD5S9jie1EluUeO+M4RXE6Xg77ve14kCTL
UBEpsMW49rC9ycOW72nghQo2P/moXgg8yoQI8uRuVOnAeJVNqtHqiz88LeMJI55INJ3AxaNzrYLI
5Z89wPpwuXYG8vI8EnnrPSiuosW8FBFn+Teibi4qVvg5I6Hz+00T+qDXklEfoulrHAiMOSFVAIWk
EbVN5r/VCHnR7t0r42s93Nsop5o3PAohdrgqLWnTYC5flwYwLtDDG89LYpFOaoPxFAth1ujtKz2e
1a5e9zPwzcFczF/PZRnBWiXrt3nby2PW0My1THFbQmB/QCodiW0b4eoSToSWKolGlj8uGFw0HIRJ
Hk0/VkMv+y9qalts3COb03zpMjn2VgMNAywt3C4pnG7ru/UfKmZr0VanTe0PeahQGj1DcoYZVEyV
5f3Z4z0yARvocoe9bEj7RnFtRzhljkeoQaTfMFU0K9SfP/uGjH+iY6GfiNjvVkQDzjZBBA6F4fMH
gxwU8TwlV0F25HVTbvDEzvGbYo1FkzhJlufYwFJqjC0DXCkzxvCMJrDeZ0k5Zna9dAx/NLCVLejQ
cK26al+1AJGimw2s0QN06OCqcNoJASQyM0NAgF2N8mXYID7XVvdEP5q7wL45lNrXqhbiakmTJYJp
8vgaYb4gUo16it/YyXak/WixQDLnCOCBZ0Am7DOCfDeH4LC+FomHh041if4rvX/NyhmU/AXS5wKs
LBwMPlzY4EYEFknFSgTn9c8T1+BF7FjFmbrY5GYByJWfvzoPL4Ply32dCBy3QJZB6Z6gNvH1EvHe
FySw5NW1LIN9iP/DI4udy79FDBtHICy7wVjmqQQ40zE03kC9Vka4lpdDulbpCtKRe5xrIMGGZW8G
mqJCG5N/3xEdjkkrC2ofGvUHWLdb18L6+Ved1UtQQxnkGnzT0kA4Vsml68jWQByodV8uNH373uxm
2q0mWOQPXUVAmHV77FvEZe5XrsSlxuR1whnwHBdBXD7j/EmMFiPVMa/liaqQjN7mwF+Rx8PadZq6
p0VI9vt5UvDU3VswFiB738R3K91m6xyyDlq1XQh6HhsapvGHKEyV44089OzWkBs3YjAgfOTRrxe8
mnXQhrQF/N1Tq2V4lA0Zkkg+w+/qUuC2QjdRyZlxggu/r5edXEr64ULV4ZG9LKhiWvPF5A4EmZfK
ew0mEvZDGFJwctOUfsLKYJgnLLDQBpjv3C7IfRHUG3YAkpT8TPvAOQRTrHQAzPHFpRuIi49AwhCu
A0Eu/rK1TKeA3Qze36KY5hu25sNSoTGaSTveSkFZGckk11eoOq2Fth7G8nP2i0kGX/Y5/ZranNue
XubsfNuujxcqu/Y0JVtoeKFl10GVwjEE/ROWT+zyzq7SbxAW8JFUBArBm9USbiHmJk6C4E/RyoSc
bHz/3kbhHevfi4emOABC8E1JQJhsBLhJNvym4HJBUyia9JbRAXSm5blXUqr9topeK0GTRv2+SJx6
LIWN1tHAFJubP5y3JobWcAjAZTz1sPkWXRkcRrQiPQNcwyWq5SqGeQ2RUZtwNpvK7DzKt160a3Oy
97W7rPIzCFsfYyCZbs4tPlU6h2UEGCy/cpIxfNC9d7GyywgQsgz41HqKdyjjmDFm5TX36YZoicNR
tFtNeggGKHnXesa072J9OHS8NjA3wuOsJXZsaNeBz2XlrJ+PFybRWaZKDYoW9OS5lpsfksLwbh54
FuiLQl0S0gFklljHwHy1lUXqDsnrGc05wgW6cCXfQWitg8pU2qoN+Onxya3QL6WQAvm3PrAOPRCY
jzB2PSeP+5aGCFFggppbt4Uu9Iv9XWgAwCQat/AGnYyFJ+QlpayeQA24pzlN1Nzxn6/QaAEf3GGe
bx1KIt9udCNpaBQzf9BQnwKkDRK+MR8zbolX/UJK8V2feovAo/9VN9G+gRbkBt3hBlGlmYjM6Wl7
gaLUi3QTL4qykXZwVGNKI+2H3dudrq2W1AJF3KVI6dxsDup8XMexYDx2lJai/JHRD5d6cqGQ8p9T
w4HLl9BluczPlgcqkFTMK+GeSm4+oUtLra1mK+Y/bnTcCv/ta1Q1JKG7zIMH2wqGl5pR7jX9Wo3y
aZem88A8PBqFnTWImR1WWPhArNMyGofqafvoBqDc5od56Ma2F7+/jqU5Q7FEk9DZnx6b0ljAgvBY
yfZdhZ1AvaTkDgHWXOWSp5BEnpRqZ5aEZxgjSxWk4pR62lawPOdx5JNwj5BBq/D8mmYztLmER0bT
aaDge6VxrN1tw1pINJVMz9ARhDKPhbZTwiip2QP5sgSciPFJnR/r7sh6hxURKA2KeMvR5F0c0Mt3
Xvx+9JRqZ8l9mRTvqeCGaOG6E3KjEgbTIQUdkwOkfzqhWNNfh65Wv6tGCfS6SE7gnX/HuPXD/W6l
v9IbLRw8uCBUAWsvcd8WxDqiyy0s9saKew/QyKdq5UgZDUuHy0lz0St+cR6y57wzCDzJ3Fk46FeS
XkFIFAByHI+74Ik3nIr830Uii4DO3zpjcgC9RmFKsHwIWK1vcXM45wlKgnmXFMx9av7KsDacymYg
Q1ueK4aG1SMIeEXnCHBMPDew0HLYuQO+mO7dcqOfN+I6ae9q1yPskncV8RIuNRXhNgbaV+V9Tz7r
todSX0i1vbMSiSbGn38594VhUWFoeP0DNMWnT2AO9XwdaVmWrzTGzYB+Alpi+aaMIJBTq30leL8b
XNC5THa1MZXUH9Wji5U2M+Cvq6akO/tRtoaSL9XGhROe8HBhb7zWitBnANAs+TifVaSmnXT4VxDl
QGqJuzw4X1Rl7vpRZkUTOnwfj3VkjsilW4POSbDZDMfvY/kWXjsefbgyM5TjUYViRNGMMyqDw+45
/gnvIoy/fRKuyG2+fdZz0+FhYm3HuXnWcHaxTO3d7fgbVje9hAALTYYcGxcFasLybaRiEXk3KRQc
uSyZVBE0DH7UMje+XRB1pjKSh2/32Gg+jqF1ARMJUA66YKnQCgkKyubaYaDw/QnBH5Ml+PV3c6bK
MJeubxcq21+y66TnfCdMq4VNno5OCGJUMMhUJHGPVkOlBnAno1sZwyYtsq+tXEHm4VaZ/qR/rviT
XZkG3eK7w1F46/0oMPelFQ4oHm9zCzf02L1uZ8y1aONAddzLSXzPsxuklZYClPXbapyPIoZ9VLwn
TScGteMhujrwB9Be4htA33bkndh4DeH7zxlyfoGfGaDOGscGDdT9C3UXojXr3QCILEPmVQOpJ9Oz
4DiQ+55RAN7x+Z5UT4i5MRgy/TeHiJo98lw5s/MtQsLfwoKvValcE1UXkq+mgj+iZZB1rvTOfNso
FYSXli/BH6ZA/2jzk8bwUAnY60MrJv0l+RPpS+qVsjrdLAhnQtNYEAbfJrI0YMzuoXElgFRQgErJ
lFzBJF6dKLVmazSGVeglogmCbjNsbJIT3q/YO461BUu0WBZwOdjEWY5+9Fi798iu3Tw851aL+l8M
StWUfF1lSI4vcYt7mUBBRo0N3hHhnJWmxfhC8B2B5TL+UWYDeKEtGUEA23kWUyBvwxkLdclI87Cm
GVZEQFDnYOxepQS8Ehc2T99gEby5jstTP/o/5PS3ElYVk4Gkz+YsNWKlkb0K0TEru8RIAXBoaD8F
GWaWAC3QdHRMxef6wXcXPMLyTkPwj2FmZJoF9Jg//bRv7RIAExTQSwskAPImKYCZu4w5HmGXQtv3
v639KXw6wRtZsvqGMkiZtq14YzaRliDHR/AJbL5MLKGlYAh6r8eY+OqmO8wG/bO8avV6COujfRJ2
EMkl2ubOVWl1Fux1A8o1TOiv0UVqg2ZN63QSlXjOm/r/QZD5qOAg4T4ByW/hUr3aKcF25UdqEh7k
EVHh9k3dCNiWmy+B+hAFwrhJGNCDy925A85KHvsbucjbiQ6bsD9yuJhM7nauir0XWi0wFHWRqiq+
pT008W27k5BRdo29mn2Q1v9MPOD8DGNdS0YSb/RDYWJYXOcWItqCQR4z3nqPBePw99K1ytET4tCZ
KoLihKrWPa1kLfgLnCMSXvQ7VtUOv9Gjlf0qOrz02t/Q+PhU7cJIStaDltvesv4l00b7hY0Xkcjf
GnEAxrPm3+10liG+ihwj2L+Q8szsiXSiNUphbhCWp6lfn9xW9QVT8G0p0cdRB+S7vuByq0Qlb+en
b6GLE3PeA8jmW/Sborr4D+0hYBZf+BdyEVAbWGxvHVZnTcoEym8UoLXBFPvLcK7piRBT8aqveYcS
o0A2eHNQzTKRooFt6iJ+Qm+6zJLHtXRp+HhfbzsGCJIbXFBf8AqbaJCoARDXZ9xLcD9YHVRGCcaK
I+Rt5GuUO9+UDVFd4WHVDVkDaAXDnoJ2masTGtl95sWzHYKEsk8P+0tc5MpVY5h19oWTq++2JwuI
/HOKtKN7ewx5oPuyvGLeJtj6r+KzSooE2pDMtxV54hIqOo4nUmnUdnvfznorN+CDt+1ZdLoA4cUR
gGT2oPEwePK6Kvl7uI5LTomE8yKtKzWzs1iwp/YVNtuIiEBfh9pthDlScpeb/VjrY+PZKipRlCBg
XWnZr3+xMo8Wotn+ANuFEYkBJKm0NkYvfokD1rNPd/xDVdViPJIOR0jbGsDrdnBpfcTIHMj+Tb+p
S3ZcfK5y3Zjt9Ja7dWUjcddCwkAtpSjlKzanaLDGLIQV1Pnfj+L8bqcUNFfK5EUSgIl0kteBGKQU
u0jxe9XuI+La0J4nOuZr2Stp4MLumVeI/IyhX8X6jA8CJOGbp93dzrFK2IvCqFecu77BtstvSk4M
Z1ucB5Rnj4Kzz1eDhTRTZ+RonObbHXarCSNEb+9Np1EoJv3Pl8SzqSfDKZ8ZXSuDHt0u6Aqt1GQ8
Ok1vV87Mxtlwr8rNeT+B4dC86U7itAjLbEC9r6yM2R+icpZ9STiaEVsnOe6zLoDhV56Bzkhp++ds
lbtnkvlqYIP+W3aINFskSwBzZaX6qOABHue56thdSe0rsAmF1Sg10Fd1InkioEu8gwAIGRn/DW/S
lLYM0BayZj+v457Sjg+L/NQvk25zaRkXIJb2XlobzK64fKH76aVH+CzOs2HTYBTwd1+bbZ4NaSNz
Zx8zKZG124JPPvqVDKOcEA4jGevflRM5Z+srMMVcrOpfD4W8hnL7kyt+HU+LgpK9XPNbtpJUeMXj
lgbS5je12Cuhk9P18qWf1iktGYewRyJcvyNGRW4F61yrHFzLWFj7/bHAKe/GzDWtpVdUMFuYnRCY
JiLR2/tg8/RueLuUtABKVTR6RrUMQI0M8qPQqEqUv7KY4Ki6bwMF5Ep6vkFqCIOHW4za1QuuKEbN
A80LTl4vuYbOCy3kAsv7o99cNWL6WiG54Hw3+H8cc22DV2IraA+Yl9EUquD/cCPBFdVT6+2V0YWF
ZJse8symOxglO46xc1GpAgU6Z88cRmRg2d9FYqHs85tHgs79ljVtoUaOx6jM0vw7vRO7y8g4bWCP
JXe3UDIQAQfkcFzBeK0xSfb4VvzPm2GwKAkyPjt+SSgBstc/TY/cLF+aQzQbn5F+OwiFn+i6+m3M
/gC6xNQZQl3S8+JzQapfdmSPBp6yC/RZk0CRAgTFnFvA3ZWVozAkBRr4h7q3mQIDQ/k9Wj7EK9Af
/ScILF3xNFloqTkAMmdLP2ev2dtGjXKMUAhfLAHbf6CkxJyxM+bXwHBAsQnYXKpVPv1xYn6pUycw
xwniNP7koS+wM7n5fHBK09Yh/Iopiu7Dxhh/NFoQgE79Lyv3WhN1u74sWZBrTWlOkGdg8NajQCyZ
vSc4GZ27yP5P0jju+OGVJ338fmrG3pqddwcN3t8cJ2OegZtq2ZDt2ph7QQ/kig1BioUfwqnoGsII
QnceEz1Oy1gW1ZSfgBVOTdubrTiaE1s3hwjRLtH5ZmWWU8i0IUD/GZIcuQnkrs2x2yRXMlpKm1nT
Xd0nALQickFJO8kWdGCIwGvXR27wW5uYYeO2PwY1FOBViOhtkMSiVIfdPqkMYYlEez7MhNYf14hw
u1U2C2/fACxeGdokcEk/5n0Bdibyl7Zvlbafuf1uePvlr2g5YfGOSTN3ZurcCprLWZ7riyRxkSMw
A9X8nTQm39Fp6rzf7CEi8wdHrPdT4NptHatHitya7G2qZr7IZE4fegJ7CfoinlnoXW95K6RVcQ7D
/rktzEXK7y5L2qkwDsTFbsZXY2MeZU+EmbtejIXjO47mv0IKTGeJ8zyOqIGaZLEOKSDt+h/e6xkS
nFiNqFKxYiGxRDgW+tYLt6uRwipenAw00RP2Wga/C2zupbN5H7JRVDYuK3OG/43VJyIApAhPVIyn
1VYOVrSwRuf2FEMZeCDUxKkiAWUIpVFCpS1QvPxjyXqIWmHrJ04Zdyuv06DVJG9zI8bcKrslZ7Bp
/B2RBcPd5dv2c+AQY9bpfa6M3zIBhxEvN10SSSR4Nq5jnHlp5S1OGcYV/f9KHHbqjTcS0R26EmPj
+OawVu+TP2Y5A5y0deLPbXsSYu//5MNBhrHqB73IP1WZQSsl1Zolv+MMs82P2yFdye6I5G6wtlow
oKfI7F2NE58owDlZSmeiDEtZ5L6jzXoEV9ybPLO2afwh+wBd8Atvz8eabsac2bAx+8+jfm65d1xT
r9hQtiVrtRnYhxIgKtlSmhswpxhamY8EIG7w41kvxr96S7+7md3vE9ZhKPxmzeiIqu8+WTi5a3v5
7memdRrJ8GL3Z9VXWbJftefpoeB7hQYrDmmWvW1uQZ0H63YWpUxYNheOwysCTH74FmpLYoZFGVHd
DdAF3K8GhPduiTq2zKVN9rbDf74JJQa6IwsOEKstgejh6za34hf8RWA8/GlLZ+8uzVj6DVY5qVeJ
Va4LucGotUeHRwqFBK+lb74MzvzsfmPMmis4C+wm6rkP5NX4tbCjwyVJP2wbGIxsl5dDlzD0aWRy
CSUfXcazzwu4aBkXDy4ea/y+UX6RdUBPqcQfGO/mumsZWK8oWErjuKZZezigWXQtXt1t01icdrTa
8kkTTzkAza4cEsETYn8BaXkbtpekdh9AnNnLzHOxBa4CbHoXLoLC9L/9hpUEsWJe+lgxQYzexlFa
drsO7CRUMm4MAV4andV2rO8njzbRqAcJTvc8lqjpdrhX7NkJoxBwMZ74+Rp2rmm9tDH6nNgeCeNb
4fyLvjGUk2GjQAFZN+0/hN8/HXQPaS+zNHaYEVSeF+uWyhB7MuE7OOJnycvMAit54sP/daavPpaQ
574A9bqBXF8s9Bk0VPQd1EPCQ+IZJbQp041KK9Whz9EgnIwrcv9oPd0+T1J2KxZWYZwXc7DIX5R6
K0EXFkfxizBKUpZ+MwBjZsMZa0RV9XDLlSYTwPi49lw6KQ39G7ZUIQy8TEjFNScli+ntaBBhnDk5
PXO4fMpx9sk00jZDCn9bqFA7vgaRFAuyJn5ZAXmPjIBJ9DeOiG6x9il3U/T+hAD/kt0vwWQ/Qp4a
mOJUpOFoKkoyKliyTMlJfGe5xiVDOVqnLQUV+Mn4WZNjn/J3Yv7ZCQiW2PnoPyqQpowzc4LPINAf
eZTf9vJzaFSyKD2L/DmmOnZV40wefRQ7SA7dtd4VOAThPGQvMACGujyqh9KAlZ0yICpFYEJaLXgH
+YpXxo8UZyG/xnfTW54yNsdltAahAjODRPiJaUNhE2f1dYUC4BagZd8pTxc/b4O4RpN6HyR9aLp2
T/J6M8MCmKr2T8rI+DdONVrnu+pk5sL6rJKQ6bkrvw5mIaOP3maZAMRt318Bey2cD2pqJ/Op8jIW
Zsqp1Y2hBEegkgH2s0GWIHzhrIR/aUthXxsSjDO5NVhcA80Rp3fnKCkGV3JO516tKCj+NN/n6REJ
lseYPqC3hCnzM5mG56TETBTN1YCiFI89+TlRshMQIeZ61KRQ0tTi8yZdVDlRFzl1osEYcLW67pCT
h9CZFYv4F1J7XUi+ssmATKGE5oBQs9knzZ0dyr/YycLYosouwWbUzfMht5ILCrtl17sCPKfBlXiP
OpxgKJP0KENeUXxMJIc+jM07fcrqP+ohJYaJLjc/44uCFxdgXOMBhGwbZ9UEq09lGy+TBRKrwsKC
SUggjQ50GlLtILNC6dxPoyusEIod02DAnM5YzZxSBuWgPTfEmci5kSV5xUu7mqq9tFFXeasJudiv
H3dYN2l2Smeo35cjq0xOCFy8QWe+T1Yuj4iNVe+NGEdEWHsvfQkyRGf7FALT7gQTsj7XMHjdCh6Q
x71i8Fbs66oMSwBu5JFZXKU+Q5BH5xuUF0Omlcoq9ak3RXKLthAF/HTxoaJpfh70V8ubtn7rOrT5
umQk816z/Oui7uvcb8GSqYmGVu0qrbN7IrsVJLmWwCSITyXCNrMYfqZBpfaA/v05aKPrUWsAerBv
EAU43ZF4MUFaoB5yh5zKWioaqXNacitP5Lspt4TRFW5GfwSvKewc4EPpCFfJxVhPzH5/Ux7oa2aG
nLPEGRoBZ0zqXq24KLNh0Qd8NyqcjSlpv3e1/k+w8RvCKA5F2DoHHRr5XMoWM59kb8R52rQh6AdF
c28WVT1r1C7hqzm1cK3qts9URbVbIfjo7KdpjuXlYV74bGnNxpwMpGQJ+Ny+BlNM9ez6MVFTfPsf
PrOMAk1GsxxWqZaIT7yNHOvCWs0PD5Md3o7XsrPkwSMAJRzmgT5Gwj1OsWpIKWyuxwr+0VWCLqdi
O8LQGHwEqMzPVFN3Pnkw0X6Ew4PyYMiJBiK4zvKNW7+STkncA/ZZePSfG6SpaW+zug+qm7xBgQu7
xMDmndm2jZHYH8b0luwuRvQgg1Gz8H+hLDSAkN+MHHYP62MfO1DdPJSqnYd1FEt2x0Xt/mFM+VJX
zzhX+WKadRiiUmPtRgCrKCL+zDhbMPBSBeJhP9kBw8hT6ir94in4QIrAmIo49j8wi45WwLIYJyYi
djz7KlprC0Y/yqO4XR7J5Y99q/gVCZlOHbiJ7WhheEAI2+4wJ8T06+5LFbUxaqfqOXZ1gaQhlV+G
MzSoi4CuvQFFVzdKZIW24RF2RWfbdilw/rXYxE6nTWBbA3aQtLBvK2nBZyq8yOsev2hpdfOpgDf6
Q3AUBbuN2+n31AYMlxBEtSgCRnODt63weFonoXUzctxDE+AcEXLXiRoMR5ktMdpLjv5b1gS7RwWM
xRa6XmAfVp0QDQO9koUH7rwPZSel5pI5sJyWnvo3CLHUCfuYQ9ahdBuGDHV6NPI2wOOm8coAcBdJ
qPG/dw/bgkOhS8y2A4LGUdJm/b4i1FwfJR5Zk433/1yjvIbU9M3F+hmwHBTFJao3SwqqgMf7JbbD
/MUVOMcFU8RXmbvUvxNvKhCP7kXnuADzRnMirsHufFMd96YCPgKYmCw1dufIrnmZS/N+w6bNruKo
9Uk6kT61qIhoWGb5kg9x5a9cfgg1I3K/PDNjx4pcL9Hb2APK1qmXeKMTU/dJG/RxtHR0+ynfr80E
2kZwm6nyXVhjfyUHLaAYpqV7grCPRCSgH42Lesx4dR4vJBgFJrQOLhImKyUtYGSajysoVGImT6cr
/r2yFcShr8ZYbiI6MGrVDtJJ3CewH8uK6RZRy6Hn8azIwSWswi0QVlRAfPnZMiZRlT/5Y6RmCB9a
RITL9fNjoc7KKMOVkzC3jMQJGVpU+1vmOgsdaZtqRHwdvz3XBNTYPoKLJuZj4F/PZaiosOT76OQV
5/bQsbqmJpKGVViFyLL7zlNZSiiomRVKxPQsEoR2CSURKJdKwOqgpM0KiUO1AmHDdAhfQPiSJL+o
NpFkwJWYngD55I3M3s8voI+2a9bnkToUyNpzZQQ7QlOFvNXaOavpxn90UYtVOUDlDZ8i16C4WAS+
ofh5VKUoR1ipjXLCx3A+i4N1g5DJqEZiMg551iOsH3bdhvopNJ9uC43gMHZpCnIJYE0dGwu7pctF
nZ85B298ySxWlABwzH9vjHQS4Heg+pPVOYIwo+5T5m9n9iTWb9v9mQf7JsOlWLdZTRGWQSWL6Qnp
hudk+jyEEExWNj+3SCNvW5yvrEbFy6o2GslRL0ruT5jQY3STJ851/K1966Y6Di4sTjeQS8krMB46
QZzK7j7N9tUkHXlD5rwNd9cqFuIir+nqX8fpO29cIURGM1Xhi+dJwwFdERHzzxGV7OU/oa8J6ge8
2KppZoDwNHeCdLqBJevWGeTy6NugS6e+H77TcDazWJO0DpH4RrUxxTnUZclkqRljAqJN0kKWXPnB
p9X6WoNhmSQoDA3FAB+aJFOfQiMZljvIAUsWmikNoOg3JgcRqeh+1smq+9cisd+hT1PVMRel3Dw2
XBQ6Lhyi7ztW2hSkKljH1loZxmjLfBGLQHzD+3UPRhm0cYlrjPfX7TjMTAiAacH0+qVkXkpprrGs
3TzivhJf8XgaMA834QB7/lkyA5f9ohqSa8y3zf2sptDLmyiitdG4Nv8s0Yy7zIjBM+CJCk81nXXS
qKKAFxhYkuHm6afD7vjlRu61vJ5uUxm70ormdtntkfSB321q72voPekiCrVkfiw0MEn0MfDRy9Km
A7xBtNwkQX8QbztnNEmjj1Lb33GrGKVD6uPJ5Flf7Kc15k2qRh0HANJFWsV2Ax7dUOZp7rVtWdQF
BlAgRKOnLhHanZY6MpG/HJ3N/BOnz33BZ6zxN6IpOuK9QNcpPUbitlnX+Ix8ajHzPw0Kz6imo5va
UHplvPCqYBbnU/C+Hln3NL/Pj05qO1w4uDK5xiBMbzcagN4+PlSchjrIc0LjnMqc7Nly60cvxqAP
cnTevUUI8nOn6p2U8VBj8WKb0c+UHQuhC5XfCKx8hneIJHvsmDTc2BugwSPqJBS7S4t16dth9xGJ
IdQISGBjs6bs+jwM4qJHCRh45Dov+RiCftnpaltQ9dWEr22huDyQ/pm7UGNtFNPAapOrqdl3e3pI
aSaU8KeuJbG9RFX+5qGxe2ASp2VlP8K8vkFH27T9mjw3n0lUn4sZNirJkp1NTschAEMDwh8K4xlq
737gsWSoyNjXiIrMhc/zJ7gD61SlDbHI/QWgaAl/aux0qFF21C2Vnfatd03Hu1FJ/6VxbzQkj/yP
L3+OW9pfWtoRejWTWKSgSuGBGvmA94Sa6zjIuqVcfP5K1ZhLc+72N2dW17wOvBToKjk+Sz/q/MW7
8zYFP8Ly/Q8S/0bZ1jIPpzvnBobw2oOlO8nGuYjA7LvM2qM0uOoxcvvVDSVzaDlgXrfFHoR7PhsB
FaIH237cp0aubi5zAikPful9pWZCB19c2XvuntS8C90e33EnnrI9XLDmwlJ8y0Xu+ifHzNQaN3N9
qqb7DL5IXcWc1mdE+oVJHDX7EA/IllNrz1pIunRMPomTrwuXk73ut1Y9242IUr/ygIPm+szKnxh8
FZym8e3UufPU9UpwQxljO251FkFqLDSQ/X+fUXZBmP/ea4AO06x4wPD0ZU80mfjkexPh/dyrlWCR
idYR/45nQ93PPapv7UpgCHkO5kbJzICwyMR84DANaGDkfnrgWL2jXnCm97sJTVTYR7LaKHjsxFu2
ys61k74M07YLOzg+nrY9zAzay4brpiNECm5k9SqXX/gKut3KJzSEKaHc+IlPwa2qWbkjktRkbbEw
nEohnm+nUzyw5Css11C0Nj86n9/gKjgj7uFP+Tx/gYnd9EWLbxj37CnVWfbQ+Nx/xOZqlkAlIysV
6+r+AJuY7NZUoi5zfzdXZJueIg7ayMB86ikeWaIb3SL3RBkTsmyEf9MFTmljuL4UZtF5+5VxyZeg
een6mtKovYmzGNHvt4rWn5ed9DDRkYofEZWzqfwE5UKzejbBhsrZCxAZhIXxBUtnkoPdy2S4YHAm
33HemrEP+ZjSmj+pReUmyi2gxhMszIVhYdsyPofIsX2psCaaT4z3UdB8THMPXzHlMKtZZlCe5RDy
38lh0emRaFYgtz2PsANKZEm7PgDPyGS2x0B1XWx2Jq9JYSfAhVAq31pTLp7hEKh5h4ZUZdMycmXR
6vI1yANogamC61gcWlTaiG5E59RTtOiEibht6q5ycvUfKD6uO19ZP2O8DqxI2AiOznHqBlN0/ITA
s453K0t/9jV3uXbnGLd3pArXitiZXz1pmZlLxfPUHPU4BBgNmSMLsSdTJZL35Pm8picbbkb5C+g7
OFesOJWE6O6ijSqSAcoik7toMqXE5DPY+V8X+1joa9CH6YZHkHGkhVgngrAZtyysH71+8jnN+FLp
PvwVWlDeCVcr7DFUXbvVMylcBWtnu7VWDoE8QLYR1PEB3C1vCmRnmfT6a3VkAslZJLsUGnQA/a4W
gBpwA9fvw+zT0rhxvircb1yigedQioXnP94gC8iBKvOQWfsCFvqa2B6tk5jXGkP9qZaY3ujQfw8m
U+5pkrwhfruPmGvRRDfPT/mp5EMojnl08aDI0NEeam6dlnsr7rmo1to17oHB6j3lS3YPkrH5Z0/g
FSgjAyFK25N6rIE0609OPhn6CIyahNAN7pD/1hwDuGsfiHpu1E7diCoi7cNqpD6gN5QhsUH1vS/s
TMcK2khDT5pczylEWvTh8VKmUx3y8hligpGNJlWN4aLEvKgHpVp3ApZD35GNwLEZqpLDIuRwJh/2
RDN4uVOTCmZjb/zYPc6NOOrlxvF+/bhBHDVGqXuGR+Px+r2XYipW/xmeZPuROLqJLXeNOTP52gz5
QIjcCtFjNwrzdWvz0vMr+2klV7fE1b5euusDmEyMsIfzFhiqhRVCIjQkHZwonBgk0N7R9uCgOIea
dL87cMzPO/osG8E+Teqz8wEnf4yYSu/0ooYe2kKORpiJtX3fRSbNl1L6+Cx0p/lQ7fSvs8ddpLtY
Cp4B+vF0bNMQuN+kUS7dU1sIQQEGltJO1tdjgmM1skxpIIRkWjaF+gZuP9+tJ8LZVK3tw3Q0QB++
zsUKrCpIoVxPkJUuRq0JjyW+KEUJUG2bnnJv/9vXJp0PHyJB4+COZjL6+QJuBHWmwq5n0y4Gd2SM
eGE0xbQ8CZr8/ChkjBzH86cN1fZpzLx+6tDmzv64Fzr+gP33Cj7suBNE38yflukMmi7VcPTMP5SC
NNGnHl7IHVp7k6kRAo7NDC+teO9esSJELZpwTeSHgAEDoyW72rlVacQmjQN7z4Y1piOViEZoTvmb
1MNQmTaUsAdxzEbJZdOwoukPPn+xX54jDFEk1EKBSCao2VVpYBqPC8w00qsNZ+KS1kXlkE5TqYmC
cHyiPD0HWaUUTWd0J606Z2UyiGeKNE+lxKkUksdrpT+2FHX2cMbotrDsmD6VsJNF45d2k5UPrC4Q
gVnRyAOUJ7snTzjtJ+pZa0dkA+FmFVWfJKAc7Q+damrFwbJ34MN9LQlpIQyssW5EupX3t25vpkDU
JXuLgUKbSziVAeAu8TiVw+qKScDHRRDtO7aNkdYl6aLkbideV0Wly5LFBDq8r91OGOG5Ya/gVpBF
0xNKU6IE8+BCEd0bYbtYRff9MujBscbpJkKiLSowXOEKmcQ35mXybrtLDWQRmp6of9BoikzS0E6O
tMqjPSBSlNvmL5a8kMeAc8/zuRfNi66lBFqpnvYiJxc6wafnCNDIVBaY2VqcF7LsMBii83flTgR2
Pf04NwrmDIQe0GhNfQwPjlWDt/5gsp8LyG3OoR4pAmO84AM7/8wqp3rswP0hVYI9SOcv/B6D2+n8
DMqZjlXQSNWq1cNDyKEyfJHemuh+h0//0T4GuES1GxwyXQ53o/icG1/ZTWGPoHkHw4WKY6sm2OHt
iA25JMA25Kn4Urv61a38ORmcz9T/I8Qm3MbLV1VgIDzAusvqN9o0gWmK3MDQqtfWgXEBDaj7OuRI
bX7uIovAHd4SA8y7BjqIUQTyPLy421IUyNElylQPORjLbtKmWK5hMFYL/5kcTOCj5AD9ljoAVSZ3
18ypRRwmU+XxCmdhfFJAJcwFrkWkS+6DRxnuqSsAqQ4QWcVpzix07QaNs8OR4u2geW3egt9BbuB1
n0V/4rSAMjG4Np6Anct+oCeozEl500KetNIcGv+UUuNytfYKlyVmjaVmuHXinbBOh3Ce/tbQgx2I
mdNop10SDMtlrwS50KjAEE0K6qGVgSyt90werzAoi7LADYdN2zATaHyxyFT3EaKcxQrj/EfaMxEm
rlVHlos+5n2hk7fksOE7q2ilS/246cYDtw0SH1N7hSFfr0xrz6Fg+cwSmrBeFSK3CwTzlOJ8/Dvd
vyuEPj2yjHp5FL463m4xHm+YGYwbNSAZl14NiU903NDNDoZidjui2fZFmnP3uxsXukqFHGtqrlHV
K4gHa4ohqI+cLgsccKKJNXm2HlV2p1TVZhmmG3g4ddefTxKviiAJPqwc2nTy7QsQ/hJNgbjp5ZaO
rEUtL+5otmL0rx5U1D+ou8z4VICY7uF131cdkKpGvgPkwZuPVgu1AQ5SZDfRxDb+pUBATaVhHHw1
uF/g4oF+WSVy9t+X01l2vmHuX/UlQkegu28dM0P74tU8eM74qWZALwBXBkZSEmqd4wO08bRldbUQ
l85i850MUdZ54oxFgL4j2J/W62FpOS5VWwcgyaEqFdb1QKmJ3PfZxVYRdQAIq4WHf42l3MfwgWWM
aDjbUqUNv026UZ4VaBgZ922DOx1XjOdbjxpBRdkYl1oAlHYabR+dNLI1bPN5r2Y75gkc75qcmxVD
2vjazs4eDo64Y7JKKyYIbJG79CgL2tBLrRjeEp198k91FJf+klwaKcCn8u0xwAiSQ/eRx9GUaize
OQa/Ca/gmYQ8kC7+FVw5AN+IgBB+NoiQdXUFyETQLHmU2lCOvrLSuSSQtpdN2xWcQqVJQ8fzjk9Z
VCnsOM1ysxbaWFr/j89fD9x0bIFnbnsrFR1y8YIIfqd9ONNUUj+ncD9XvZvfEFRVrnfO5pLkffNV
6Mxl3H+WU6+kbmJXly28vVPm7qMCvB010sXqixxum122QbEFkA6FrfmGFR3I9zansqbZeI/u/f1g
lkNgwml3LI21M3ZUmFqp5D+3/oBUcMOKEnblOyXGClL1GMJprTqHAZnsGtp0Tmp+RKoG5k8NqTs7
AHL/ikRvv/d8zJLGs27BHDD09+Dyjooliv6gxETFqjUh4xvOpuO3oDiQuWab50JxJ/MMSaSiDR6i
4BMcLTg877FJSA1EgFHROsxQKs//lU4hdhYf5VXNiMu1ycQ5kJEG4Unl3gMVAx0SAJCiMTyspGL3
YGsLs3OAqycplqQxgiBQ4NxSMHoW2eUag4sHjhB2podwDuPjn1y5cxSWbZLAKLWzX0+thMKzvGr4
OY9FNn+L03aVpe7lNrZEmPOarZQPls3+46Pr6DZYxhYVoTBJ53X26SEKkRyWJQ2XwH9oyyd8Iw13
Z7s02PHUjd2MW6piI+BE/LQl+Zao5g4yRgmnLjxlvGNqRV61WEcYRyQR4/GMONjYm7J1Iguj/mgu
AE8D6FI0a760Z5lwyPH+BPZfftR0Y/uP5siPDRxC1pIQaFqdHaLxO0jrXmqhKytavSKF2dpOC5fJ
ZAA5UxCmd20kMekXiyWQYs+Ua6cAuoyVb/wwBcyoAQo7XupwTENbZ6GkyjeXW563OgJGs+HkQgo6
LfEMUgVqHRmvhrTtbaYRpLMn7su5MKAIZzn6v+lZonYFOMmGZM9QkqpS1tbZa7TlQx8hT469XNxg
aTMo6TPFuahcQejLRQpGDemH6CpNYQnnv1ND3c1VxqBJA8ycXAhwcPN0s0NLpq5bkDGzirDw8AXh
1apEgtOu8x0aOgxs4g5W8wtA5YaeAzNg2hjB912lfWvX3+muJzSJua9EibiF1vDlhrt3zo1FNOGR
3Y9OI8bGYFMHHCfXdgBYb7M40Ar2QFyDYMbcC1QpNHtRJCI7vQ0AWQqjXDJHMIxpQWtkjYtCxDip
XRF7a5iQ68eqZjtZ9ANOLmpcBAidR44/lUVavYblv70IvGWgKy+ql80a8IhGkdv++4vEuoSQqTeP
EuQPTBHfcONmHbSZVNUV2YEEpulqL8DMlru8F7GHXByJmDtBWnJJT4fNUc1B02fcRhkulgvSRD8Z
+Hcgde0L8kd5DiCF3rMt8ngju2GVemBelOhiorOS9R9YlCTmyAbXu1zpxwqjGDm2QWwbkh7Wvo7n
PzSU2YFuXGxNEVzWSPYT3PTYhydXCevbaDEXWO993W8a5ZMMEDpb3CSkAW5aAwx9A0kZMbHrYdVD
sUJx074C666uYh/eRqLPZv3ebadjrWQqt013LjI78WGoRsD2xspfCfwp5MGEAD+U3AcBCF8jftwW
fRyjKeBEpBOjTttBNOuYoeCQF9QsIBUaiy4ffHS0VRsAdI6W8wqpTYmPElbqUQcN8OvKTs3pi/I5
DlX9/rJC7QKwtkuXd9Psh2/FtA3Fd8eNTMtq29YyIOsIMyr8TiDusn2s/ZQJw99wSaST/VdbQRyk
EJ5rMrmyS7TsX476Qjm4NBPmyVNTt0E9mxCPcQi5Ty8uSS6StijYfisMgKSMBPs3EoTpZmmSgEm/
qktDXjInS+qnHNKyulFl0pSrADvn9zI8kzkyk0cQvllS7mILKwVWtwH5hAbhc63zKvq+9knmFXNv
41OiZmGBmG6aqFrLBeiFwyolssNLb484jmzRHR2u4wbI8wiiBhQsyt+PJLVymKL14L7cR80xUGl1
we5F0D6an7Iyk2LkD+fVxd2E8p6ybQ9efO2m/m2kUVT5bGIklFbj+FYj3fFEwTEtUL/GbbHR7+Iq
h8JJhoP4qH778GgujbgMvwKf6vRJcapdq8m2YHEVPTrEsvDp84Q1nTZjzc101q4vMT0gsBDmtell
IjmSQ5+Oc3nS61IL1ZC2FgqUaEm7UBWajWx6gU/iobVc5uhJ8KrA2AxkT/iC+bmeeiMsw8SRwTvc
iu93tex+e4AoWGSp95lVyLSh69nXugVxz7pI4GlvRdOBntxluDZbfrRvY2hUszCnsFmozW803zIf
a0ZzdHklrMt95sdvBpnox1kINZ96N4wevC7EHzR0KkY9QGSoeBOgCrv39BuxUCQ4iSAc85rnxygc
u/XRwcg6qiZRgqL+es7uHyHpoPAejUHaL+YNQy6+InrBuEGaBT7sW9+vrNO4Rj9YWLfOtRqLgc/N
IzRnqxZZMN+alr2Tc6zwrTXUN8DO+Fdi1GmT59xj2UKSIXZkwfZkgRTm9a5YAMJP4RgyHUkAJAKX
SkTkdkRNOhSLIZKtGKcDwd3IBYrhInTC1U2WI7BuruarONa6voGiVfuTGHORB8maDoYywRh+Id3W
+c7COBgfAZrkbiKkFqNa2Z6AAMJ6TNfSLb+ccnWOw/7QPQIbr4/CcDDFn/m/tdDT3TkFo0xbn6Kc
KcKBa4dvWnpUbi+tftdJKvcRieYI8K0AiT/42S6I4AEWbvcIaKMMDHXd79WSNOQ2rBLpuOsMJfmO
0r4PpktctxbtU3QOK4oyd4cSJVIQI5GN2mhwmvC+LPxChQE06w1R3lhBskn19YCYYdE0HArEPMgX
mfIT1b/Tqc/GxTcqLZCdpKSG5w+QqW+oIFCcbnopKPFk9WvHGcnOvvFhQyF3UAFp1hsxa0q9kF0y
YPn1E5vz3YJSYybIOvO11VOVa77uooZdutB0kkTIvuLWtZYZgFbfDNmgpC0gxG4JOztqtiCloApg
TQLARVLbKC5jns66DA0llIAyz1RskYJrrP0mWVQ/KJYOdc+iSVG1WocDApAXyL+BYMCNTOF3wKZo
0/Ya3TYS7VMUXKBoAnOCAIjIuzbLuxz5/+ZMK7byF7vdQyt+Lp96+BQQ/7KAQdhK+0yQBdvRiZzN
QTxZmhY8jC+/GwamrUgUu9XKWX0x69v5tirrDu5NZ1Rg5rREn/24s8gsgAiYaWleT2fcKeV6/irz
FK78NTdZ5gmSNMqWgqnT8/h7AAjgOWUkAJpKVaNxb7gH43GnLpQIqiY5BFGEZ4RrtyqRvaBzKEDZ
PreYscruorVTdO3gVNrTkIx9bNlM+1Y+6J7p2YhpP2sXEH87h9l6z6QRt3S2fqXyKuTLjQl8GdXt
oYVNQ+69DIh+MAlbu2yt2zVDIdk1F7DOYZOnO/KAzJnH6PVBtKXbyR6dmJZLr2UPQ7jm6rQnKsBB
8AHPy/5FxVu+Xo2KGQ4FL9CyW/98Og9KWEUGJ7M4gA19is0sSdY+X4W0KJ9wm9tCvxSzAUiYf9uz
O7C5EPwnvlApMuyaKbmIXu2bxdxoD3+UKcnt34oliRbAyCRC31htFDR6VQwokkErLfxP25xaMKQH
CMqMMUlp+tcVwjp/LTTYni5C9BrsdU7llNBPDi2yJjskDpQKF4OjcHozZ5r79apHnCvrrcfrBaAD
kgojiZ9moSLSuYZ7xrgw4Yn7uqKNC2lfthWDNVBMPBQxUurjkvf8pE0w/B86R71dg2+yg7yYcxSV
a01/ezeDhQLxWScgA8Ujt96IQzNWE0fhadpM5lTWyf1YU33ET6dal0Si6JE3u4G0KJhstj6o8hVd
xZuh0/qxBXNshMauD8UbRwaQxQxQnQxpN3gFfFB781cUolBPmFPCX1P4f8uU/+i9mCFvGyTLMNKg
/BuQCzqhWMjH9JVsYAmBnl5EP4oUAzG6espr+l1p//XLgZWQQPpy7HPtVm2RGoy8xJoqQQF8ftDb
7fyWN6MHRvt7OIGgWQ3nlkUuvAJcWLX+0F694TttQ87q+6fvupsdxYseuNokimiq0xtgkGdDJR5X
pYouz/lYPjtOONx9tb2uPnfaio21BG+jNmxk1FLO2qBH8+2NDrGAk3k4dcEtsJIanjAgQRHHM5X8
k6DKfDG+HMYf/GexKnTWTaPE5OHCRtUDn0b+pzHjb/qaFDl7+zlGZ7Cwr+joVDIDndP0qheEJ9Zc
HDj0hnSuIz3+Q0weFygEt25obTzbBSGBvQOU3cr+Zk7DWYyOAiCOQp8CePQCwv+gJmV9tFCwIeTk
KZ/m1+ufjCYMT5dTKOgV+1Wfhfnkvp+6fSGVG3uGKudgEcKaWh/ECLZF04T7ZcbZK0JNRCrib7za
Gu82YJFbdIFrs5IipPj5aMH9GQ6zAlEq/pK2IEQTZpiO4U9DeWbA6SeOGEqukLsMXPdcwbmvWUtv
2t1/eFWeV2GOc68oy7m/RD0VvtQtY6SIVyEgAu47x1TkjFJHZ9I3O499qXYeN+dt9Z9CwsQ8RHp1
r1j0bbxIZh6Bf9kpzkRR83wfmtfvkEoNylCDzQgQ93ZUNhNvoQpjgNNw7a6rieZeEgnvr2Mt7PqK
FIET+nrC+GrylOAZP5er29d8+B2gRu3rUfGy/S7qgT+4krK9I3Evel/YlClkAYszOGxu9Fx7WVRB
sMFbbDyKC0yheizSiPBe/v32aZEmC2IQuw3Q+Z0NnVL2SKRIEA97oK9TyLBmhkA6CCyv3l+Lpldx
L7sZasrXGYHBCEcjPzaNJggsDcTlb6AiCmKp0rRRXfnSyBN+TfZuBEI+yTxkpgDLnKERqhHUrpln
Rr2GSUq5OOYwZBjx7y5gvpX1xPoKeFRdo4gwTJIN/kEieXL7i84IJf6edJsGuJfGhkUdU94PU63l
uIcST8j4J7HT/36ioeu8YU0qkjspmRrUvb1D9jEzoEywyovC3F067yGGZzz1WG2tLbEiS/xm0Ra+
43kdVLa3csAjyWJXZlJAfUJkCE/g1vLZh96yZ6+WhBfUk7EVNAinDpjeEoK2BsRicwmOU2GBk5Xz
/o4R79lMAboC0vjeDls4M5U1zoeF9pMBB3pokS28IIaXy2D39nZkMeCvVccfn923Gxb5PqjOfU3Y
r+76587nDF4aMibTZAYKLZw+h1r4AnlWc1L6qk9ZGg1FPW0jWW3YwQmveZIQ27tr2WPdu58GTfoD
kVTKfwy4ENP/oucKmagw2B8DhbFvv0mwtlj/4eb/g97MJXL5t/qPNZB1OAEPE6NlrANPx//cKh3l
v3rKt7jpwxoSo8tgY2pE/a87AQYcxo8eMWwxCuftvy8hprQzIaCdHa8PzIMM7E7smEj7iLV8aNRM
nxFxmiHyoCweAtN46ROrFnHOy/P3oKztA1R2+lwxmYLXzC3CHqvuVmy+qnz4aOLR+Gs8+0QeanuT
cARtwp9XxPIeRdC5VShHaExuX6nIJixnB8HaXrZvprk7mcYHW5APmMoAIeV3Ais8ySr4q8Sewbp2
KeLIvg1wTivoR6wQW68CveLNXKhD9W53Eavucx+19udMp2FNE3vZ4+J50HCvO6S9hkcC2rOm0MUa
xELgv3uxG688ldG/YAY7Pk3YGZF/odGHrIneOqP29kwtbsQYxUA4zSUGv5KhiT3vaRDcT9MloAZk
SVpDnoPgZ+s0Q1cacon4ZIZLedeX7YAZJmjr0kjIloC6VRb1gjBdP6nULwA6wG+tZpdnMTUZYBiJ
QgUgUhdEX8eri+o2AoAmMNBi6CzCENd29gqaaD8lvCMv4hL05+h1cC80cM2Sljfp+6FQ9Rds/0JK
Hd7MJqG6PsPW99bBGOPra05NEuq13NaBYOX2cC/3FVrZozNcqJhhRBsTFILV86pvYwa2tUT8C+sv
oVquGQDOST9rBFdjJBKe06SmZ481GAZp9+QRavSBoB9V7AoL8bYkJPMEY5yc7tbZHCurVLvJm4+g
f90MQTn4KOiwspeiqx61MjLILCUuNmhrKDnA64/8vcbUwXegdWv9xqZ/+3BPs/TXCQQRhSJkHfO2
3i3qVUsmfliS0qgv83xxxCmDZbu9VqLqpaVxKycOGCMqI2wEGi68yvkEVl8vpoJmyszmB0vF0s7r
gXe+QDCcE1nY9RDvxOu8C9u9q1fEfHTuDjx7LhEY+UjAEcUIAPkol4IPjQoZ1p3mcpm/+wQu1Toe
jklh+c458cp7Ve8mXGWHr3x9zGUTgjyrJY3U9utLG8QlOOQMrI9RrCPQN1nJ6Id5bvtpW2Hrh5La
Bkg+mzQ5k7FrkgD4dzj9fVbgQOjHRxLZKx2v7yEkrRfY9u/Y4dm+C1Ya+r1aHW4ZlsbxxTSObrnZ
NGyvW6QnA2CmCNlkZGSBBRN6l6t2T1DMTQP1erllU1W34Eyv4cs8Os9UBxE2cWD7JhSdIGZ6hPUL
Qe78Ca3jqHV4rH1SGNZK5NcNVsCWl8JAUbd3p1JYDm7e/0ZIQN9LL7Pyo1C2WLuclPaFs+gUykky
YaoVcmq07fcsn+NZmzYtyEAoIixmGcoURxiKMO5dGLGo0Q67xAPpCN3h9HqUcwodQE11p68gvENk
K9MuKDb61D+mNl/tYJJUU9bKZnw3j3v0TbRKO6fGjP7rAbEW0kIOAc1MZqIogKJ2T+NQGKmWkJNH
+MYxprvAhQ+9Z9jFH+C5RxEPFlEVF9CbWLS+Vzt0b73Ugd/1xMQYJT5IijAeyK3IobkG0cLHtrv6
3Fgdu7iUk4PSQlnVdqKRgYqNxCeidfbkhMf6CEByYUXbIsCc9uXBt2o3R4IEfJ2oWi4o7vqDInGF
f42HlAf5zZzuaispKzxPMQ05GvCdoZSMaxiNkS3AmOX7mMJHEnMBrRp3VCiL4jewRFZnvbT4ijt5
HMC6zKYApJyLq5H7Xv+ngU/oMLIOxqILI87X/eNbqDAUBpyYWo31HT0ejlyUKu8JS6wPpMXLhvD4
avxjUuXvxY6CUJBL8kG4q5Mif3S7iAhV7F8r8IrjiCf2Bu4pXOx+oPut4bIe9q0KsVQHEqHS12eq
WHFwu7cmydEV+3r8mIE/Q3IYI273Yt5VOO0RlNodHeOGtCLFoQdaGO9H3HpWp2fIodaMNT4b/FVt
adoVaQaBDdMmCvcTjxyp44vdObbSO2E/aXD2O9C/cGy6gRTVzQsCz9rsEWmFeeWwKan3hGpqBija
1VCMIhGsYcVHtmPvoO90IuDzdl3+eUNFld8q0ecAGLMLEacBF/Cdiplxq9PSTrk7uuGpGheCzTpv
jsAiY6KVkWSq4U8AQ6Zwcb6WJcS80P3di8UNW+7KdXT8KqUVYMystiAOAPgzNmZO1Ot+bWND75Nn
30qnvu2bLLzXmd5WAZ0wp4VtSAphb+F26eBB+rkLn8oUv+dkbVRuIfQNJmCzQDE7S2r2wnif57S1
gmZcsYrcpy1jZ0dlmHQJYqXWCxic1DdPnNH7vdGmOlaahrb8e6T1yGxm9qzidwyF6cB9g8s4aMM9
jBn+kn4JZAtXO6ytVAYM/ItPuOhR+f5Y5FQMJeEKAHUfR9Rx3B+HacdQk39P4mYQ3xIcojRYehma
NOtLL6MJpSF+SEtd/4kYLaW0t2+9FeOFNPYlf7N/9zkLNUQNaLLkDfaYBwSXkLWoC7kGHwtVKS+G
JLZYpsDL4VPtcKfNuUlTAlVoUhFcuyWhofTHr4CuhJSFaY9/E5Q9XO0o31dwB9T9+kXdX2pmhGfD
EXYv8ZS+RbghmIU8GE3c60f2XixZpHsa+AZ2jFY8ukF3ut3Lfk9DuL6Gt2UOVf6IA7XV70Z9HuJt
Zz+aAkd9FQppjI34Xh9tS9GOOuEnqJPsK7dX+1RA9E/9fJ1+dZNYoi9SB+xGhSwyyMPLCSo35hq+
DX6IOtpBGDbleT0EIiFDxnW9I+AI80OvuouBxr7I7O5xLI3FMK3MGSTKmz8V4CPHmu4xctnZ0gK9
P+6IDMgoU2omVhGKcDC83sRff9uo9bOU9R69dtvsxO+t3nBLXV+43jcJnHh+RuHytLCDcebyvsTn
jf73G0gvBcIUiX2bWkifSnpJWqKRZuy/MPEvfRwpmCcoun8n/3agSsPVznxmE9kLh8UFJTIT+jT/
pI80cZYMZoiIOs/5UkbzY2vAOD8eEC9zQxCsPCjQRzWF6u/DeB7Wd8j5n04XcadML/tk03DS4mbu
T8fsakv1wATuD1AR04vTg6601d6D6yg3JFjoiamW4JH1BGY2UGk/fvoA02X8f5niyctdXC4l1Vga
G/9xcgkTiQxLGRNruPwsQ/sqSexMZNxUNa/ryHZW6QOTSs35LvoXoRhlMH6k8g2skD06WmqziZVn
DLPI8CwPz3VvocBTLhWRb7ydo+gYT4NQn7K59rZGRw6sqMnjoFk2BQ6lK20mn5xw3ODPwFoVc3FY
FxwLXZBX64kLyOfXhE2qel7EX7ZVJq5MLHj0Bxw7jCt16a4qw/mAjMXceGVOjkpaBWM+EW5kg4Ub
TObhxFkZ2z1G0v4lTmQ/1SDe0uJ42CVolihWklX+hmD2a1YpjQpaNh4LY2BJNT69RDDuTSA2Jfsb
4JvKcxPWhd0rnwnIABj0tmb6Nb6IdrH1HSDMrp33xU0/m81ki3vwpDpjnLuYWzyNk5kb8cxZnszA
OZIj8AcIxKaP2/aFUg2jaR73+xWx3kiqljDHmBBKW1Bm8d+It5kl7duKqo996nC6kfeoWu2vQPHY
1NYcFquRZwITlr8dU4OA15OklPhsWCnOpOZ4EubovUaOWQiX7L+Tbly6UNWo3jpOv1ivk20pZura
6V7gVzKo1bmLxTXgMSK+vZV3B8T/4iQjbSIfWGZ+ugam06uSNIuk4ho0w2ZGhxzp1Cx3bSSsOwPK
WBVf/qsfY9kH6JNG6ZEAo6GYZxgzKR36sQbzfgGuyMfiv/9rEEH490IM02IQT++2FyLk38XSLdBS
iVBEB0I4STnm5Isr3IXwVqEkzBqyFjFjlzhe1Ymw1D7iEmqtN1w8rgZAdYeuksOd/qs2Ri69FtMO
70ZDp0I1jVeQWWCpimG6Yl/sKR1QfyUj4xFw2OrC3ZM+ak2A9BqO16pyTieiQdhliRHcYXBerps6
JdQm5QjQ8YGJURP6yEffsOKAVto6yMynp0mBWOM8zQjUaXJxswsz6XNfzfUP4Fpuv4u8zNvHauT3
UzeW++TDSQM9nhwLt4Enk9FXbi5hFqumrPA+5o6HlrCM9s4hDJmlbMET9BOA0ulx+zKNMLlDKg7x
c5LcD4QWou2LA/pC1d9fCbwC3X0a6nTFjEK+BsKfzNM1l4ZrkHMaUez4+MypQZo0jmblIHRun5a0
h3PTaIoIP94Zb4GMKPF9dqPngtGDekOFz9sNUH+CXtBd4brIfT94jwrLwnoXLbDHkL56d+d0IEwc
xVQaUqgpE5VfEfVCdUDSks4Cju6fwDxyLmlXrqg9xKf1weHboC4znm+iUPjPE/t6QrljE2Ne+6n3
/sbxd/OkVtGdiZeVBhmFrPI3UeKukrXwxgXTShWvGnBvK1dkMYD18k/+m4AkKeXEWcc7QhP4wEaG
tjioEkpRwnUpoHvRTGpWO8zaZH8p6oJC0Zj+vUBJvwJUlKir8qRBqcrzvylmI/WaVuQt+NXMZyPB
qojs0nCaWJgCETVsV77sqZ2kRBld3lkgsZ44ic8wNlqG9AViYhnL+Zg5OxA3w1xabEP6Mi9j1KYI
M8Ia29yhtiXzrYvXdHaXk1Ymv7Oz9vCkiEddN30TmmSn4IFemq2rinecdk2iZgFMF635ZEfVx/1G
FuycYQi6d9ewsWu7VKogTPiIkS2fELOcFY/JLbETqUuOuBtIZRFS8NQuG93JZJFH2OAPNEcJuoGm
UJ4E+Ds5D2rxBGpbTkrpWFuPMFdZDz72lhXzsPSPtcU2Dcj+G/rHokVfR18UUlfETiwXx4BedBdn
1396HPeqq7lGHvDeZopFr20KAhqRyeJ/sU6/DjQuMbwk94jUvj3LsKqba6LtjoQjXq+uyRiWcKdP
oBf2gG65pxieKk11jp45OoneJEMcR5CTR3eZJFnVDOtB9hLiKddy7NJfjdsJneMPgggTdLa16mhh
ZuLQucSwEW1yP5cqDtDFnGFKWAY8O/nEWYPcOhWUJBMPLlF6S+UYl5iGfDndCklUJcroufOd9ArQ
JBznVNSp/mBqs8ZS0SG2GMrivwB+GqTlvQXPB+1JBZyXIN+mh9emm33x/jZb3L2nAcaPu0fEnaQv
zlmEowwNGYg1UTkUjVcBnvygO4GIcpzVShAaGJlKcA8w6c86a5k3OB+dyE+6RPTrzDYx3aUxpnMh
9GZ+7mEyfR0vU7o/lW65pcvMKa7EFX5YmdvoXZDkcTZO5C1ckpsKaNpaqVBcSxzeEijnThhYiw7A
9b1zUYhmx24Kr5wlriOX5pbe+aRQIvKIvLUS4ygcS4i/LgZFPumQsjl3lIOom117/4jlFVzmMRfJ
G9YsGwgQD0tAujxQQsaEHe9qtw8gqrFCLJEIk6GTTuieigEoJ+7KY8oS0m2rZMhmlk4NjH3FtvDk
pMnLzLwQyyJkOSpdzoxoJxnHfbn2ZSGAIyFsKF3aeD0tB4NwjsUNAQMklM5dn8vioJXlOcLLH1pz
i3DJRQm2l309sMLsN32DWeGo6izAxqEVs+2nBlgVp2wrPW2Ir/3BzbEBvkwd41C23b9xEXAPPyAm
hge5OTy9KmQJ7EwsyKFtL4y/QpvHQ8wBo2dG9oBGSPceiQoLmzgFEYBa5IGtNzIF65k0nPtB9+2F
rZYvCQHMjkEl+sALRf8mrg3+2UleBbp5gdraKBvFH6JH8YaeMuTGsHqDQjfo7RtDQ7C0+TTdwrq4
Hg6lTeivs5DhzPZMJCpESPhmzkGQn8YjOQPcRqMiOaIa+kAOtHrkwLKFv2EIPbeAmqIVu50c/PCY
s2HpYf5K2s2ak/La7cqne7S0Uf1Q84coP2alzbOdcX6YM3oa0HYTxCJNgo7t8ntxH6GUM5vo9mQH
NYpv4fboFwcemh5DIJgf4XaTReKWpuVakq+IotBHFp4ZRhgfk33h/IYxXwk2Qn8a0JoZ8Dz9VGT/
U6BGERy4KI0X8fCADmJ5zHbuv07JzSggptIYNW+Si4prrd7fmfe11ZbOZKvc/Co4OyMDR3IhO/Fr
4PCoHNu1WLU5c+43NrxyRyo9g53Oe9kIamJl2VOhk5eN4mGjrk95pA8+AQ3nweahvG6OEGgiYTUK
mk7iDcOmSEATGm1OqRgNH54JZr9jsRMDLKtYxf3YYOle7jc1bNuKDwOR6DiIe91D+kxMTn4HLPSY
h0gfhD4puvXBbAkg1UwE8kllSq54XXS73MLa3Jf8LhM/NaD3Ctylfd0lwwHqcz3WtMXHrYw8iUlv
Qb/meQXQh80LgQf1IBhFNVrfIwNFtwULrIQiWohDxFM4pzP4dyDEYBbLQhCiXCcvaXqNlGw5kNa9
JWZ+VhtDVKCdp9gHqwiU9mHBoRBTLWmhC4FZPDmgIWjs/hmw4gXdB3y3+Mhf4PQAfDuCyxUeTtwA
Mw4SbnMwACyZYsf3GqeSoUn5FFotOneLP/sDhVM3iA26FvRVgbqvPZyE/cfWlA2VGI3MY/EqxUr9
etnoT7ydusNZVOtC3KSDuPHdT/+0oCpRU78IUcDbUgg7j2YnYRa2GTsjNbaSz3Od7FB0Y85YjuUH
zo1RN85MEjZ8yBpBCJr9AcugtYMUbY63/mgIEjOCHn6X4OTutzSf4z1auB3B8gfYheQHKYLA0wiU
y/vwu0IUfS90YQT7sO1HGCOSCltwTObOSENtnhe9wQ/+L5mhQd5/9jwuN1kLRYzrMJoDNoPn0fbw
j7xfY64UbKewWC/1Io12KcxsFx9TZapDyCQOoD1udzmiKA6rYehrJe/F+iHZoo3BdjxCT16XsPMo
h2DfOIWvRb665ZB+aJLDpG8MKWl4CopoAS4RD+ammbxiUSL1ejduR7boUDgoYolFP5JPTWWO7fMw
jlKzwTmdAH26xAPrQO2nlPKARM6My6wrH8WNzqgtKI6tmF1sGydMb2eJGHK+/x4ujScpsrslA110
4jtz5eYfaY92z+wuBKkVHwsE3VC+brQlJu3UyV0rHsseYo4QK0jezKSRe0vdHTG+bU6Q7Zh1uYxD
YguA8cAeiZ7YwBdfyWAcHCihTuXOUAnTUSRIuJrYyeQcINOHR5sSMKjR3s2TaDBdsJoENe04wXtC
y5Tfo6tncp3PpmhKAlzHgJZKBhrDYDTyFIigBLFfecy/tC58LozR3iNFLcYNGGWdLwrMX1U99M7F
j5g89+BK7uYL8qRxf8WTkVHAqJlx432T2vVu0mLs36g/76QR1COgzphLkH0t9j/qNcmMsrscHWro
vFaa4v7dFcA5p7QG2dA48mFZ+xzvbE33bz7s0ClGgG3HVLufLlA4SIPLekkol/V7dEjmIshTwpYh
XmA9vd5Eg903TwLC1yHpNVHX23Ii0Dn8qBtIstnZDlcDdjOLQpZTEySSe9RfLIWgIjDMI7aDP9bD
pp41R6SqjEMEx+ZqHhhX6GDa2q1JrTahVHnWbjzkkEsVIgjw/N30pUrDt4DbhCUyO5MPj9qLWcq9
BCkd/1vCZyP0alddhyGU46Co0+SYLkxBQTknGtvYGAx5ZY60zLeDnvZItcpATiLCU7li5UDa3znr
hEmqE9C+YUPsqmq6p5EV9Nzf44NOAlQxwiRtfN7ZcI/V+8HKlUythll0+3Syj4jNoUWO4Atv2x9j
yggOsKuI3AoCrDAATRZN3BaWtDg8mVU68K56A3V/zCDneFciGeSJUKPrgBrWXYNCDoPhz1B60lJW
WdvHbk+IvKrhyMuaG9ZTYUbDn0gba7KR+NwfKPJYkdUli2qrcyFEbpP5cvD3WrW/uQvrUUVnyhLl
Dk1ty67KYQv7LB2Z6xBkg3ce4Icq+LtAJghHcwYNhQcViOt8qn2pP5EU9EaSJ5my2Ae5I31tsXK0
jW7Yw6Cd+2FxckJl3dTyRpoNFoNGm7VFd4T/PtZmJvDdtD9RSnQjea+p1Elbxs6X1knyE0Wbxnvr
zmpFHNPxGBvVS7zlgLD8+FejrmWUqNgs0p3okCDvMNXgDDlCn7UzWi2L5YyYd9yF5FmuG+p7rksk
ZBNATqaZOMMGwoBHTtYGMCuOfCP0PkNFUwpN7sMdA1setnTps9LS7942fpMwQfbgz/OzFGGCOyLE
BNiTS8zkGUjX1kUHP9PT84CkoaHvIvSR7MNADyxqJeFAlWZ1W0h2JD8b7sfzBeKpEfYijuUvl1Nt
Vyh4CDG2LtJ7sWX/OGY/V4GpYCU4675kWCqIup31VOW71s1HFMIevs9HY+9CexcY0cyXEdZ2kZ64
UomABS87TJ2KISu9MEr+i0cb3OvAMIi14YNFwwbetOP/SquEy7Gwq7mdqIsvrL4oyy4+BPkCrh4Q
rUvoMmhNZ2UB7lE6VEHd461w1Cu8ewOEI5+u2KZLiSnebdDIJHexqI+/5NA3n6zYzQhCS8XQhha4
jJ4RQySMLpgTcsu/BborPZe49B01ZT+7wBnAVeENgRssZIB6C/X1yK7xtyhnZZIYwmo8yKNrvjlG
1lGV/Qljwpo+OdG2J5A1TZs/avGfx5qr/iKMlkDRro63aZqFx7KuZNKYZsGQADBCwV5qR5uYF4Hc
oqQg/8XjNtDe5aoZ819zp6mEsFJ5HN9lomFrKjXdhPCEBYmU/Jxs3HhcaJGukTFuJoDWj1mpCZBd
3OWR+zOqX9nJR2xhWWDXzrpB3ysIXBJzc3PNsdJ139QPIl0NQi4Js/FTjEFs3MQ8fXgo6+UgotVQ
l0OJuAw7Vm2stKSvYHzwFNwnU+qaRWx5JQ3+b4EpQX07FMS+uM/YQvycWAx/N8/+R/tNh7dxewZM
emGVMsE0BN3Nd+oTCDxSTFWBnFIC1UxI4DA94ZyHY4TtdZndfXOi5d0GWEYMGrKgtkMzqDkqAfNi
bFkZUTO+oHoZ3OYL+qqCahayLF1FlNDe3/tm5VMiR9/JAIIekjwGX08neNEUZ/1MjHB2NTw7MURQ
uyKygUBp4pLr0T/C4RvKKDiCw9nXtNLN9jKJeD4VTbLPbWlYW5DftzWA3uhM+kiYQ3fEdhqRoZHX
W7o8PvIHcBBpb+8MRQUiclq64bArzGAbv8WZ7/Duf+8FK3rtO8pbAklWN6frturHekdn6xQ0gBkd
eQIt6Ztj/0JA0tfFglZPBPGYCExmaleL6JVKmkkQAQvNpAG+MIaWqBKX3/ZqHYN4HEBCB6HPCb7O
uyEZ45I2SzdyDGk8tg/k+R/DN7p3AK8Kkn9NL9bFHkC6XJ5M0KRsxa38NIWepFOnB8OrR9HAT/2m
Ob+Xg98CMnNcKD3rm+2hCWPSYvqDH8Ia8QU4kKc5YPa5g3BImrzA/TM5Yi2kPFUKmPnoG38AfRfh
Cva+EZ8q0KvX/UcE9kRB51VOpuM9LcK4vV79ZpdMlcrdbLu4qPXCkMlM0WfAUiDJPkHNJEthxJjG
nXFX+/DPytNXyPPEQEG4p6xVx1OkcpUOlc+kbXlt4yEPhbsYgvBXqc4kVzEpjp6n0J43q5MX++46
4etibHe6PhZQAe+/Lj3sPl32gxMm7mIBTT8/v81Nh0owqvX1nrIqOVF/Upf8pHTzTRXHsN+nc7Yf
pfprEFDVmtjldUrUl7r6aYKpjcxLnj7X9WY03wKbZf7fWwTQgHIyohEv8NYvEal5e6KQV9scgjcQ
EuglwpSdsvwpViJiun22BzWUCj8jG/1xOZcJ+uum5DOBX6HslmfGyAMDfz2nh8cu1TIQt01R/8Uk
+D9QRCFQvgtTGq8SmBlLVXb2kJYboC+3CuOU/+3v3z9Xi4YqLXedVsRpKFTFswIPf15RMVBW6bV0
DO46LOrTXK2k6NcbY1ZD0YOdE7+D0JEyjYZqRSzAvbmIXHjZwtCLZt5SnVkGCbA3NC8J0XIXzN4P
VyYRaMxzarx4yzYG3/Ypkxhik0LbWZm6O7q20PJoJPaceWKrvx6aHysEvY81FRJ1H2L56KI09Vtu
ROXiDFG3YmklIsxeXQigyhigppKyHzK4Z/7m4J3nTgYN4ImH4ufmSNlANaWc+R3TFBa1x5/JIYBk
F2U3kj+7vu9PDe6soTYoJmeqV6qzQ8EX+R3APYEzb8JyFeh3mA3vCkP9Q0GE57PDcv0t3tR4PKPn
70SHvZFCViQ1fTogBKz18FJEEdKFsMfUM3saD/Txpi3dIbQwHO+DX53XP74jrb6tH9FtexyEF6gh
H+RFDZAjANeeVpB1FAOZ6uUUseO6zovP/EcJu41IdcqChRiekQObzwVXtPD+iIF/pNR4ECKlwbVM
E+jmJtDSTtHgOMVbMzF3t+QwNDu9Yoel2zVxJQj3JkwI5N/v5ljvOLCBZ+T01fqC8O6UKra6yrMZ
hbbtXE+T3BF80642jzI+CfAIw7YjUMiwfHqOTMZTS3RGEMqB9vGEonxwOrrnNBz3GPEPCLIkm62Q
7pd4CAqFOzRs5SXdkHy83b2h5a4qgXUZh8kNFhR5mhhpLhp/4K97zaHSIS62qRgFZP5GPGfd/Ju+
u8EGpuOv1yYc2JnHAdhBqs5ob8W1Sksajbcebr6pMmAagoH4T+JMzpE7KpqKikiD6SYl5nIcrZSm
zaWH4Gskgfcf75IAp+8QSZUPFcVJcdQmXXZr4P9v0DY+/2I7/Yguq7XSBr602XuhHtg1KkCsku1d
9SlqWSnnf+1tq9U8DZV8cMC/q/gmltJmrms1q0eZANDbHOYgnaRZlxurzkVpRczflygtu2jifAJ+
QQyqXABu41xUBzHcMHylkJxTl+ImD2hid6EIOLy5OtgZRuz8M7b7XDOcZH8qCvn2TiXsiZy6XNli
hT8HzVh82nG/s7Zo7S1+2SXf6BDYUv+S/h7LaNN0xyHHBDqKaxAsfGSz7JdEZyUzHGxZRVr8ecmf
+VHG9rY9103H+AIpi7hkzQhVV/Z5cr8+6UHAtFxUJXbA/wX/6YZUdkaCysqSBktu/CjuAq44okGS
Ygx7Cxd0ix4wsLqk/Ee0rkExFZYvPmUTrVdvHzRBUcmjiENV9VxGETGDwHlqSkEjZU8mlxjQA+Bt
0M92pAZYC8T3wOxNFz4/UVae7PyrN17j/adROPZ8w3YMVomflcTja0Ld/S1g2RO32dtvFVqXaDUd
hPRJwMAdIPWAvhWJ8/NNOph/vdwSuIYjCV1FbF0R8WZGNxsX+wjR4mElTIXxP4hkuNB4/45xjzAj
KgW1N6xjXZHn0bUrV051f5hlRORVaVcCkiWq8dsqTf+kz0nJlVs8WEetuxrZgx+NrDZtUBM+7FOo
JqDcaP0jG9CSrN+6IbbXwpv3NPLNu/v+E9DndU08zLf64QfrYlenZPSPz/XnLsgmAcowP6WZIX54
dfrrthX+HN703RcLJL1CtdhIbO869HD1PK0n7J4edpAqE/flv9lRNq6w6rqJzRD6Ns3jDVdLfaW9
fPAIsa8YcNpsoV06Wl+ZUae7u/GOYodZm930PYwzZ3z2Os7nfMGySaxQh0NGgzf+YuuqM6dUzmn7
7FfJJ3CssBhUBvDPND9Aknc4l00da3ek6bEco6kIOi2lll7OfE3cDgtpFQI6LSAVEkeel7JgTlEl
qB5iQk1uNT77RIwlONNJdOtsz7Yxow9eNKxB8idJ5DqbeJsBuE3xL1xPWCEpCARBcX95/450J16B
In5ijscZiyNZ5NXXrMYqrGrGNFKzM4E33tj1G2CKSGp6Ion+cRe0khzJMCXT+URMtStm6MZU/Z/8
Verx98J01dmtPzbOtzrYg2ZklvI7X7jh0mwxwVYjDVN/AJmPGScEtafCr+9jxnrLAunJZQMbRXNJ
0duzR9Y8kme0PZ/EIrNcvq/YM2lvkdKOTUp4TyV4J+0WgxclHGHH/kSIpcP1CvRYEmMyZOQDWmWk
m8MJFX/wL2PBts+7dsFl/THUu6IuNnA5d51qfw5XDlE+Is5ChzBedUa1OtDyex9zLHWvvO8HMkD8
pEteh8NgeXtqLGa+axUtZNDH5BBzCZRtf8UB15ouwdRmYYFEOxfsOkCyQOnXN4qWgKySs3Wx6Omb
QIQcWgeJD3Z74Xd+Qu5TQa/DskIgZjAzKKAvZaqmnF8Aa+X9ouM+zxAQrO+dburIafBBpwhZZ9RA
Quk0HGvIVrfoBdmYAGTYrpM7zkO6xn5lVw1dhMftMQb3/dFpek1N/RaTbtDhSkf28/lW6JABXcFZ
df4CjApwxIKztKCUY4mmYK99Igs4rDAP9iZRWPsSV1a4HH7dnRhU4AkQNZgKbqoOQKk3K1jTPY8Q
W6/QYUmueaXSz0xfUxOOPrzT/J4en4v5gSEiVNcWMW/ie79Ob5VvOcpmHClgotegBkhpRwEhpKwc
Bv+R0asVZbuFVv1LZkGmmj7K6YgJeq9qnnaOnE7s5xpUu+4wBKbirAauB+Wx8JNMZYw43N6mSTxs
2c9SGuBHYOQ6uknEKjsPtcvo32KXysrSzwfhOOI05yrQI2VqG1JP5sHmvaomDljcz25jPZgaHxoR
eHSh6rtPdWIbrmxbos+X0I+gphIEqM+5iCHQXzIKdnWR3OPt4mBh7I+KpJyo/Q3s4/kBPfgEwZ42
N4Y61V98Ws2XcTc7CWcXh0sG1FdhLr1D1xedQ+GwAIshuEz89qlvRNkAm5uy4F136yIMdZqjl0wi
NFk/7lf6nI3XvHgp4rmWSyeCWpsJzSSUhDtQuktDRNR9ufirS3g4xHpwlhm8KvXN1SpIYw33eu28
9brRXtT0ADyiYiGs75LX5ZT9lj401ZnLFQyBiX07E/kIOtKEDbdXGkazoiPOohJ0UwsjQHGwugd7
zYYgD6DVEQpSHYmEHnf5luwR3AeE9WesB9NvP9HmNNUHdy317ebKLbQSHgJbaxZ4a+BtyB4skaiq
Shgn/zb4MgEizBIGvnDyH1NiJ+Wjhmw1f0d/eUoKDqm52zXGgi0Bjcbk1+RqOaV233mcLshWGBFS
wg4hU0aidR/EbU36MNlfCTbdHPW+baVgPLv/7+wzcfVVSUdS2r74qHmoQ6Xoe9CoZpD6OqDseSO1
62G+ZUWkNQsugBPhqtff2Le4ATjZpleknBbj+cePT8LO+QRsErrqAff8npZSdmWfdJKFv6X9HHpW
oWe77ejXyiF43FWucnJ8IU3/LvTh+vdqma0ff5N1IUeWjnA6M2EDiG8dgcUdH4URddeP4DXNXjR3
Lu5s+mZJrFdmWebA6tAy21zx1JOQpSHhWML6yf39QZm6kV6E9fqC+7DDP1TBdOpf+Abc39VzyN9s
7c8BrAs0F8423FvSKRgEdNmSv693/1ngccGBIe0WIU203DFrfUoqTQnccN3DT412aP5JzgtP0hNv
HIIO/hoI7nm5COv0bAnVTB0AkgZeO3pSH0k2ZhrgcfKZFmQdqjg/eOa9yxKD1EmMfxc/gFBhOfzl
/gRhm2Hehi8SWh3iwadHmjkqTHM0EH4ZzoUpEQGuH6J9r8TSAIOfM6b74JeLfMbMa611hg6oMHoC
T16r2KLUqj/76rtjK/2oeHnit44QM9vOv+0lLkf6mPSBsBq0lSW3nusgAi6mRiZtkHIV1l26wkuP
70b1Z6jeVyJb2Hc0aPiSh7PwmKYyoPbC3GxkTILpo2iOkNwucn3cicSa6u12iU6nKI11lUDZ0Vy4
N/aHVZKnJRHDi3wCiYovymVWGkqEUwqJrXQKix1QDORnOfRLs78jQUq/bykU1c5GGlJhUQ9PouBf
S+XkXgMArOYMSQDEMx9oPJ8kwWwa0sypIyzRvVsfn0z9tjdmuEEmwzyFtOBZ98CuT5nZhh5Gmm33
7Bs1585quYQ4TXWu+og57WLh2bzML0bOWy/tzMu0Kk+XtTcPQhRQnmChBGfCv2uBXDV2l5qp/6Av
awwxi3MO9Y/uMuCDguXYMlfYYzXtjo3vh5nFyxeNj+RS9iRw/O/7OqYkaowAs+o+enQtbuIoUOf4
Y2D09Z+vH0Miy2+z3zrrh5fC9fcU04Hck/VT2ATxT7FURQlRO6ed1tj/zrhE4+z1EGKigl5buDSN
9Q6q2i1CqqQsdYCuhGdYwSx5i7MDKGoZXoyIgewEpIbtRyCJDxwkg9PrcjZJfRTG6enp4rYG4DHO
YpaZcuKnOP2GHKk1AeZ1IoA0NbtVBZjo1GN32RsriUxQypJre9ErZrZjAr6fx9eLGDlVfWyT28ol
asQ3GJ5K1P1OK6p0XEPtAvWMbQQb4UdcNMLNn+KXH7utK1u65CSfgPTNevB41VENlBeWULQEEwH4
pClYTX0KHRJEKZhFsPV1XymqMfOmJMMjXORdAIkxHzMEDQkuvAMPaVKDYHSUU02sHwKOC3+MJiyT
rnty0ElhpE89dOXvf9gaWlMA+TQrEhJf+yRW4SYOM2nR4eOn/o9fS5m4DZFZFq+PyXoHOHTQlB8M
pMmIPrb/XTJ7tBIw2fXnClVtc5W3IIZjd7BW0yrtnSWaEX0njQ4+ppASxuDe/gGihlLBfRMiQ4v1
JE2nERh5uixDq3RmmJtwCy2j8vhYXq+AGWVHHhyYrm1WV5mAkZx57sITpoJuzCOqoBl5Cq9IoN2+
5chw20l81Iba8f+w3JBIbcHa4veYwNVdRUAEDjHD5Lfq2y8ApLIATy/wuYFC+WedE31UpJ54SqsG
hFckv+nOd+x0WCbPMsv/pny13Q5kILBS9I2jLdj72Pl7amjVei8bTzOe30+oEEGvKB9mflcZMo24
NJAwZlMeZm/zGEtOQ6kQelfME5uLZiCrH/OjgeGRqtxyl0H7FeotP4CK5wbillv3nI/6L2Wy6yfI
dv/PtvR+MvAJa+lizo/ExD0TlN+rDBicZ2LYbAqIK/z6ndkdaRp7qU8W5iZAsX8VndTbpyqzAqeA
UWWnN+bxjZwUwZU5QC90xnoj+Y60et70jQuIKYWEVG/jCLVvXeyeVZhtZlnTXoVDoi/kN4z8Re3Z
XJrq6eyOSAJZUS46864bvWRWcFue1fMC3916A3KI+bggBWV9ICM1+t8lhocRbwvdZn5otczU02IP
yRwODSbZAKemQwNg1pH7Y6XxZHcixEbJE5CQTkrlg1qjjoU89Z+YLS7XqcGMK7SQ5WPJNVaVMQkm
hyJSf3UIesdAD/YwJ63ecsRFGMEz5jmcGw3rhBArjBcsT08JNW/hNKyr9WPpr/p4v6T1t3zT3SBC
xmvSkPlguthawTetagyyswjc3aoGwRlLi5ITuDlRfWho6FBwidvIWVktm0Kp+JzgSEB+wEPebQ0E
xy2Hb8O0f0EBycDLTJ/z49dLIv/hS7e1v/AW8x8/ukOpTncn39IyogjckvAghx7Dmc8Qz9lDuLQu
+vx70oaKOA9Sh5d1JhiTV9SzqKeje5H6/rSDlpjA5eqx9JE1Vwm32I+5MwUBHZUiCtz+uPtPU5kJ
BbSNa6H+tf6s2wvF9my4/VXMPjWYgxkiXAwWkat+CUuSygRRK8fqwL11Jh7mYNkAzJPPutHhEmHg
WvL2j/dvXyQgOk1oabJK65Mlt93gofqwYN3oGlAlz9dAc++fJqkIPM5VyRKxqumVk8MqHtfR5Phj
LXtA9syf4D1+s6ylLlKJ4z0JfFHsxjiXYb0GN96EFTQj0TN+hQl+yniY1v3MFPSUIXcXPnmWwGE8
CWclQx1EciR2vAOiW1GPTqh70FqiI8Fd/tVKpffFVRDQJcmKBkmXGCe8VFM9PxnEa+5SzELwNsu3
fckgY63iSxm33w59+G9hxhzIcgboDJvgczm53ML6s0W8DEvTDOlZaGnbTrdlMcjQcM6IvZuHu9dJ
ro6KZIXXtOOwOpFd+V/VQOe98O308ZnnrCPssY+RApH7yyP04DKq/yXM8Hl+T4DsDseKvwlhDS6X
r5Ycq+NhznXt/nbouaKPjitrhmoWwznnHd8ovSoLDdnu4o1xM9zcQ+srzgt+QfkkYH/ipN3Q78tI
AIR8BLRSWSUG4k9M9KUttSUmPAtLkW4cGCXtbTTFlSq7EvRNBjsKNVryLXA9LuekT1gL8zKO7M0L
NTD9/NW30DVSAPTnwWrDQpZklZ4XdukT2+a338T4Q+bNIysE3AZCIXT7DcX4dqCKdS+GJAgax8gb
rJuhOBqE8f/5zZ9TABOVBMZl3wbnrZEHgcLEU5DcvOL2Ed4Wb9cJPAuT2IUI08Ui+ipnuDOcmHgm
24QAXt/AaEDsLY5PlvLTf2Yc0EbRZxPrT3Hjvhbb5Zmv63ujmvC0TyV/TZZfBkVBr+5D3ArfTuT2
YQE9mxbqZUAqoX1lLJb4oJmJlH8wlB+XqtQwBg44QJHiYQ7sPGXFzrvZoFv4E0Hk8AANtaoMcg+J
TcLQi7Ep906asFROB7UHix6xdNLcfdCyaqg0+u1rXJ0F8B/QpavC06EhwdebpqNpSIuQxB2jON1+
Rh1UM4RpwS3qyLWrnBygQUVDEq9fZ0+V8cCOUBanCFnlFyMxSoTugMUuUFna47MyI2FdiOZq290t
HP1qKW31Myzrjt0mySXBHp7AgeaNjrUOOz9hYrDFgHguzkPMHGsAExnChqivJ658iTXwDbSQrH++
vcEVb5n/7VCl4QULJHpU2u3Q1X23pupdT8YGP/5jYJfWsE6XgccqPN6wdHhdhTzj1tQPB9bHGm6N
Oigf3/AT1oJ2BOcyZ+ilpBRwJas0+j+LrP2ZK8vXdA/3XeRWrn/Q0oT5nlH8UMOsygS6k61riIhC
plvX/nQ8p5YnSuD9LIFDb9yrBs6++Ein0jZAUN0lP4iWZVtIvZILPVNnpxUTFly8i4nB6uavtTxj
XkANiRsFeMhA0rMgALFmlrhKUc6rdFyAZ+6noWTywVUuKJTm8abcpsDxjxUS2kBvmv+v2hPxw1RO
qU65c5lrOrZY18cYT+EySeIXo8nKBrVS4qzDuubA1cqnlfeeSw0IJTlx/EJek2BSlOk3a6MIcNYD
3CCy1LVXA6ebOtZuiglaysXbZrS2pyqnT6pxlr0TsKU8BPHuu54tEAdFcJk2zZeWOWk27glaIqoS
mqjmFhsoa9mFIHTbPdS8m0PN2PIQ7ff3N7zrK8ClvdwHM4PXiTA7fTI5UjUiLIUcmE6QCw2kzxTF
lzFx8Cknufjx4zTwsirTdbeMuo4w5rGd/mY1C6OyR3fowYb0SY1N4WYuYcXP45uNdUd0sQWvE6D0
1FmhnXDgxEsy+qZIsFEHIvOQR02qw6Se0NHu4U8wLbx4Fpa4r3OZSvcbfDWlUC/ibsQOrp7yYr7Q
rh/Fyiil3craImYnro3nFMqsZ1frlz4MDRxnML/pZ27d5i8CiaNdUA+WfLmX9qquBvBEmAuEnFCX
gU4L+UY0w+lcNZ5OkZH2MM5EZH+YC+iW4L38OQPA2LHukfIN1y/9HK2CchXC4OlSKDiYY7ZctAiE
GIQRfNJ9Y55f0BD/APcku3du8KhVzVRtKBlEkDeZbg9hBx/mdf/BYJm12mrVcZlWSNHaHKYchC1y
/fokb0wAGUApSHIBzDS2DHBVhfaJlm3M4a3S5L9adJNu/Fz2qHlh/Bx3fHGQxUe3Kwc4OrBSHXOh
4/zSxE/86HySw915HHTFjbc1TEtJAW1NWYsivOV62B1qBLs+rGtZmYpdoEODE/QIpqBf4keYrF3j
2hYbwVIatIqxDTGwOx4BHOoiMN8z1eY5EX99tu/scA4w33dP2L7VOWgYc+Hb0ZBdM+XDKcZOzGBH
mrHptNjOE/PRj8rPii6C+LagMHUIVGui6rPomdD05p+99qxLmDyDZoKHzOApFS4qfyeRAJz2lK6Y
q6geswE5nGOkmkI0hqbe4rTOk11FWJj06+bjKYnR1RWveiZWVTjexr7xil2kuRi92XzkPWJ0lFWk
3BYLxAFxmImhvxWDam8HVt4YR5OLUCIl2Srkgl1R397JNdtElkqlPBD6cQ8WgPDiS0/PGxr01ro1
XNey0/vfMVqMSn0jeY4rHO6tiTy9nPvUIiNRrAZWTA5h3hQM1zTi/gQeVdkZI5wpuuwOtNAeQ2Gw
3mJ4Bd6KgbkuWyAKNlLjMtf+qV0LRTK4KAL8P640qWgfeO0WKRgx2qMFzG6s4Fb2H6GE+50YuY48
Lyv+Dnyamll9pXotz7yNlEDo+ejroQ3MK3xSZVAz0JOY2QN9Erg9TMQsBXYFpY2alRn5sqqet/XR
5gkgG8EHlUmazPBA72N9Yn3d1bra3iKrKjAgYpFnn7MJLp5HziFavsPWsV4Ep6sM+iI/HUzFU5gh
SvitPBo48mwVq4A4DrufD8VgZt5i4dXu+x8cAm3S1eVnRu0n01UkjIXti7TEYVZQdVMqULFLT8qy
52YZgD3ywWbxEpQzKxodZN0wnOcYmAPySXAi/TO67Z88M2LpO7AFtCXYto0vJP5R1W1k9q5gI4fx
JPNjf+hRlcFMdSp06R0gBGccXFYXTfwNigtFWEK6r23SsCgjAJAEppChEJbu7M8WnA0k3J/XRLcT
1kj6ut7wrjYHwEtyfPQj9EVLOL3L4rs0anGSYnj64nmb/YnASOoxSJxgPV+z995H6FmUNItU7/Xu
loof3+xKvh/XsJdYpn5gj6FrLjEt198JKRzvUJRIMAOChVimZVaVZKtFCm2uw3GzZweQ38Ior8kq
TeVIohcqTtP/apbdhUTbXf/n+8SxKgiUDlqMH1tIHIrfMrDkQ7rGyTWZdbH3qGvZwEcolBGZtzwm
9LEYF94Q9xqDM3kqBx8EJMa4XgFMlqfn4lAYIdALNY/Ulj8ft2qdv63QMHECl9AeLj6xi2M5KOpM
Qvqs/T7OhpFnTK13SwI8vcktZofMl+JP/d0Ch9mfBxPOJSNEVA8gd2PZZnMoS1l9dh6xZ7UXurVf
L0fiRiCs2p1rc8kpn/lBhGSHeMcLzGptUG+uKtRRGbpwf1xKpIZ5mmaaXbZlDxtXtt+ScaE5WVUF
tJq5NkxaNQ0uEjMDhpA2hO9yQadGFJbsPLZJtaw+frQQQAuezPFn/F133ArmrvQ0kdCXG0jktKlO
ox0Fa3DXbvakNfF8KXxr5KKhSRYnaYx0l2UxUleQfWZw9yEGB7vymqTRdoiR6glLQ+BNAmQkZWC+
NxU7kOCAMkVDhqmiEzIDGromcIYHNlu3uL3UbvTTmeEfhj0YOBhp0RAk/NQ0LZJQMFXRvzjuPPmI
2ZEDB5wiWhMQ8W146rn4cSB2Yop+zrTy/DpnpQOs2gPqIFuilkWp0VEHbinSGoBg5TDIWonJd0Dn
6LwaHLE0KNOXqQ4c8xEM+Pm4c1i7cEHGLjRBxaOcc8o5GyLEl5RgMrEHmGOxHfJxzDv9FjQDtvMS
1NMh6J2pDY/1Mn50Txe3mg2MBJ2eqzgJ16XV00hhc0r4b4iozQA4GW8Ms+KkgI007+Q+jM4fzsZ8
qDlYja5TG2FZMg1CD5zePyz6izLoYO2XKWhNiXMZef0HSsMKrBFzshoJy4rlbHRkdR5pKZWgthC1
Zw2Gh19Og3A8oV98Ps+xZDRgwROEetmY549FYj7GPdJTIhT4pC1ZF0dEucFv28Y5r1Kx7bs+Et8f
8k7TzSRnAoqMEhexoBVK8DfwhO5pmPnEiOzFIBy235ErOdNz4069HKWE1TKIZEFEd/z2PlrIqRXo
ERrg26j3SfA6vesVZHJDEKqrW3e8PWqqnc66bc2sBLSrJcwz//OtxcF7ZkCeHDk3ilalJVOdWQLJ
zowlSnEU4chSG4I/DTIIDUJVt7hbDug7ZP10SVn7fTyoNu/FfMWmlfc/gVZo+YWYlDCI2pFjglOS
zR9kyYaAd9PtU43r19+LD6XbM5PLHNPAcq8LGF6nwe+JnxEEWTDChCpYw5d8Uiw76wxBshebFpB/
3p9KT1fBW36GGjDpwXp45R4aHqySVGUIbuxMIBRYEOgxrwhTrh3oKmjAJ8rcRGM0OFW4nNpn3DS/
kYIQ9IeNFJsqpNzLBmGXylfqD34hnqrbWoChADpel9c1Vb8c8oKFia/vMplWKGgFOmmM9qec3gLA
l8E4mI1fRz6IJ3jgFMZ/O/dbzf5Cgek2X9sLWfVGeUs6O7efLiAU4obVFGUvQaoodafVWg/hWNtF
9SrrgeqVsUaiHpYC44aTAm1ifnQ0pPj8gM8qGlEgI9z6am/Gc5wMIBFVGHvfNUNIC63E3ehq8grX
DQw1PJ1n83VwC02KcJbIp0Hz2MntRD59dwdGentuAys7uq4jP43Hgg45mvgMhJg0dKfjEsJ4OzO6
QEhWeWx91DTlb9Zg2xkD21FpbAd6OV8lDxawA1ytEvLP+bL9NVOcni/htIHUAnCftzkzggKEm3o7
S2VzelaH5RQX+IzGIzWv/d32o7590eFm7d7dW99qQnzan0M5mseWlRdpeZyxSmBtlNi3XIDavWZF
i/whowH5oiQQtPDJx105rl43dzb0t+ephDSqHTcbbt2axvxoXVxYcJDl7shCNbTLoIRAz2wg8FQZ
a/KgJYGayKveYd0u6W6UVdBVLJbdPWDmRLJNApciBF0WYfbcW8TDSM9Hasc7LNu0xq6B90061wdM
YVB88HYA2dY9i4kAli9Lgaotwn6HEIgmzy5VPgvuuUTIdCxmLssYPr+o+2+MGetO26u2AgTm0bwO
g+U4PIXO9UY/T84O75+sDLg84EhGLt7MZpzY8OBegflr4y0moTv7Xk2A4/X3R0bf3GUtavGQ8I+D
14ivjI4TxPQYZ0IFIUMer1Kt9AuV253qaVWjHSPZiju/Af01ERRXGHh2su1DB9dx6kRj7Prj/mpd
lVkwRIikZQRgVxQqlBy3F0hxmsQd0D+tFtRzTC9iAg/wXYYAIUpI9hax5GhQmVi+xBddkHU772Kb
CY05pJu4dYCvYgWMezWOqOcR4B33MYJdeD1B0/3CiIuTrCJbiwLpZ3lL9yZGlnVUEqUULMSD+2To
cco+QXAc97jMziR3UvtvCscOaW8dC2E6g7+OgP+AFnny0TMfzyg9PorjtQ+yTAeRckMlzrw8n9oC
IAJe+W3IppLDolL1oS7zoDqwFSmrJuSzxjTdS3yZuVJ8rF0QxXzrZesWSZTPqS7yV75uV/7vMN1T
qNXbj8c181kSlq8+lNwK6QN9PHXObzK4I/6kIC5S9LShuT+vkWvLyCKnu95X175yRNY5l3zgbE9i
FzKvdktp91r16VpXIbwIoPyIHn3H4oEra8Qqz5yoFH5iwqDcJiIw6iIKuvvNYwN/1yUifTvTIUrq
lufFrGcTzydeJyRCdlksJHFOzwwqhOUs7yMqIFjJpdnzosAw0uiLV3AmawWuTsaFSKsMl9bG47p4
I2gayUbCmCHjIw0YzRVQo+mCKAKOptmWOXu1VUmV7nOMWf43y7PMpt75NGI/X4nrTSnPmfG2BJM1
AeMqeQKGAIO8+3UnKNs3PQdtd7Cj3dZ/kJzlRMvyNjQfaaR8Ci75gY7vyfbYo3JV5q6R7ioZLGqW
d0dxdh931UD7670NZZ1UVDG3xhmrjX9tP+J2m5o6EqhPdo0C63UH+142l4oq+WZ9eBttAO01B/Cx
rPV37lXG2D19UcfmJ3er625oDN9hOxwNtJKxq4/UTxSRN4hsC696ex24f5vfvs+oCZxQ5Yp/QRoF
tksLmlj+8xRp+0Fq/TEO8bgxIkDNfLVPF6m71M/AeK5JFSmWbha+X98LlTFjcQvsxrz3qKOisp6R
2flWFv4zCGfyZGL8Bl98dbHBfslqbDx5VV/dDs0+adWbzeIitm8tf1NfmzSZZCWai7/YbAcMy6vM
OxaEKDkDYn3f2/BX+Njil+1WUfzTW6z3cosAh2s1lDkNZtH16UMr1ISLpoyFTPSBgAIKQcViZs2v
D2pab34RnKIn1Nw09+p7O+TYaggyBjU6EiRxnWsoGrCgwLvnkKU/Cdu4jjhEpLYEUP0z3/zWPcxz
x2a97A6tyyG45arAxhBv3/jlNmlJsjGOLeFbf4yua/eMKOZB/QYzq9ebtjdbpbm+kVXrD/+5YUjV
6KaIeTHBpl70G6uSFQuAxfzETbblDrUudomZkZtpg1IvslEaepBGyPfueZAzjrENO5aw4UkVreSG
B+Tc9MPm23WrN8TsBfeUb5lqDkdJmBpvb8of2+5OACO73Igz2Yqp3m+m5srsg0gDKtqv0rwMp4TW
O5Wiwz0pP7sKWDYatRIOhl3UmTo542fkscwNAKhKK25JAaniCE0Lb69YNpr2BgxHs7K2N7CTn2Th
okF5a0EHvWr/lKvhjY4+ZhqjkCjLro1Ybp0NXgFL83quxcmYJacRXfgQaDGpvJKIr+lPXAQvHYez
c9aAmbaFfucP7nav/sG+lspmXJU59D6QWS7bv0c/yQUlJsx6YGtD9G2Ev+/r12UESyKX2g9AQ0s/
YePNjs9bNUFvK3vxsPd9UR/5qop0kFo/3f+/dtzFC3lHsOnhVBUyS5iecDjfQe3fZgU4iVQjKFGl
LTPX4Zdq0Ue9MqtcTMAfpNRFGNDakq6lefXB2e8GBAvuu/dwwmLAvx4jwWAbVEqzE+XhtW0h6Y1L
v8XLApSi90DEm6optzUchIJ2DLFtuNdGM9vPd2ZIJcPh1vM2LTbP8YK4OIIr2N6bPJ4hNU1XBD/o
IKR2iHN2LSn/nHGPiZ0Vf32XKdAw80Tr+7iH71XmTGuVSAiwyd8schWSfFuE/bTu9l4WIbn0rI/o
TaCQRMoWnxD3A/ZZIouSuYSXJjTMyWZoEGD5gaF9LdRk4VXUQrwwz/nhTyQYf4xBIiYI9zisJNKV
OBVxoge5VvFGUK6B7dAikQjH7hjvHD2Xojso2TXD3L4xZyrFSS6eYPKz1av9nf4Rokzm122rp6P5
Yuqiiz2n9s3ytZxHYFJB3grriVsFTg27mtXDIVaVReqySqE9xYTAdureVmjpSghzjYyxvdrupTlb
61hY944Zyje9IMs6Csqd0hDzEAnEd/JMBXKG/cZbhOCvDo84XaCF4e3DL7zeZSgVBQDmXnfm3H92
KEXr32ONA0ziEmFLmwrwla5D7zLf4rrVs4q327R/C0wpu+mZ0hdGRn7UMoD1qlq4smj+vU/Lprle
WynGGct2VyghoF9suKASXl0RZvKD7Dpax4Ec7IZesKEnfLp6VM9H0Dzf6ffRZk5dCjLL7BkS01O6
OTCdENlXjKiTSgQur/DYzvDBmIPSgRD+Z5euxmQhOfINEjOmLTOQZ4xbhUyF0M5NwBVKNmE4m3X3
Rx1+RrOF+4jHTBh6Imy7sh2IjmfdaXT8Y1xtUmAyr5jvebcCq8OHJ2AQHBJPT1wqw59hXyn9D2qr
pIWUwJ4/0KLZByIL64zYPgp/rst5oxW/RCCGpHBrR2MBdwkqIUg41ls6zpk7owwBtVCvpe2zTR2R
ApxDTvlfck713E8kdzxXhreeWJig/08kw/ZUm/Q5Ueo1zihUMDWJcGoEzWktOXOGMDdrpiFi/y5b
OKLeXeuc2wUQXd8QituTiQ5Zca3UCofrS9kz/bwnXFo0JiIQvtXJWPX4ha+QsR/8gsMM7Dm7PX0r
5XV+1kap/jLZr/cXs6GBOGWR7YVWsswEmRikt3i2y9OsjQShuUR3ZQzHnUakHY+3g+4X6wmrNyBh
6ErTIhRZpXJHWfVPmQEsuTHjld3qVHJfOJUnUljf9XRIBaWw2wgDqVwuNhpuwEvzORylO+rPTRuq
J35t0FB6ACjhpQm4lTzubzV1+/r62NF7Ac07MKx4x9+MM+gBe0ImpbQMMFkQ825tgOEgH1/g6Vny
s8KshpmSByy/1qIcyDk+sCub48lyfxAr8od3TblV14AdMmSgDU6FHe4Krv1mUD5RXUx759p7iFeR
Vjh9pkiTxlwN4dEQR6r/Tb9p4LoPcexAKfWo2eUSwSo8PLtV/9q66fxF0Ve3iks4H5xfMf0FFSw3
HHaQkJmBCyD6MDTBekKrbZSnI3MLVv/MXCWmqpr/87XAAMfG1CQnrE3OcyW9FLA0W/i9JCPLsCXx
7BF7fB2Ln3drX6ojJOXNPmtBQ9oNdBuE/uAX5evIYZIQ3kdQs+Y8lee/hZ6WkPvkUd7OW7jsKVOU
VjTN2NnATNAOwxn/FLyGEsk6tFRbqC+KfovnGvk8bPXX5NDDlfvyKX/Nfie3FpUhLPkTwLApRYRS
xhEWuOFOwFL6Lp+uAvR3ZxaCEunyKlkNC3mTh5B1EHNY1q4WaIcZNw1E4d3GDJBU3NLlQhxnJUl4
0nOeUgmIz/HMkWFebUiw1qCd/9dmD40kWIyk8cPclNOiXwLwYKgUjLrtZlWX+3eVgV7vyngK0Gzu
aXXk4smn5WObcIS4Fjk6tnhBuzYOU7G3+Uo7jrrzEivarhjAddOw8u4uTT59VYebPwKBJZLudKlZ
9FmkNXtO1ZiLLecY48lTPfg9qzfTWF3T15dZpEKdvHUalHQHJZj0ZPu61Pb/khNxyDu4y21kI7s8
sVTk0qWRMM4AVbBijwHyqV6v1QSEs2RvgedK1oPZnx0eGcliCGPJ3tyCj0fpQAjMJ0QLoYcjb8vX
L6OtPkzRp0LaTFxtaJDm5igh7Fx5B3SnXYGFkuh5DRv6eOKZrWuv6eWlKwZVlpyFXhX0CnmzmPeP
XyyCLHcOth0KBqyYfGdG37tK6N3w1YszPxof44lDjEdQNhmTK+7zCY2Qkvyx20861Tx0r2ckNsRi
Vui0S/staLYfGcFg1O0vJ68mEKa3ide4pFDbdQYVfCu6hNHX1h2nc7X+eSnTwwE0oHm5KGEkrWbO
C86jFzjHZz+X2C2adlqEmHLI+aH7OLapTgWX26iWGPiKwlks6YGU5s3FsHUkPnq7x1qiktB9kN60
h0yb4A8ksdax6SmVPKFbPRMMHgMv4vW5IUvLufW2hlrX99YwLMtUAaNYPE+MeyFIZbFb1dDqlPzP
DlsUyTFU0gzoa8W7jGYybbFEyH7h14HSDFZw/HzUD8uirLL3RMSCqrR0za27l1UG/sZocMG8O6hl
/JkngluWSfLhrbUAwqMxsyWiJ2vPcSj+trOPQmyxOX//oGcBpae9JVv7F893Zt3PewRb8jnKChGu
Xfl8h1Xfolh76i1MjUwGRhiPXfKHQJ3Lo/Rypd7+h5VwoSK4l77RcTLZBetO6TZuU6tTj30ebLe6
fb2XO0QefO5y8FfDwbg/3dpK1GItgDcT7+hdhliumX0+LLf3JmxvifsfRksNBx6Usx0kzyc0Kr9z
Szkzws5NP5CbS+ieeRniW2xJBVbHZr6YLDQHt4EyODEHVwstRhT1W1/JlZMONYr+13awJKTFI3c+
xiy+lkEXM0N2xxGRe2WLO5Q/uVq5l0Nx0fi6qWUXP3fcW9hOP0B0NVx5LexsabaqmBOiIUkREu89
ttFTUeOvw8cyBJB7lml0uOQiMSJw6S+B7WF3NSjqtlXs5rniUYGSaoZ7FKgB9FZdDNlYNyohli7u
SovEDGzoPqVnfrk0UyqVd7vmIkciQXTjq5DIciR+2JRvSzYfnjdJimlLt+GxEWDaam17TvwIz9TE
QyDVhbUuOEPBxa2H8oF1CwNCytOz7c/Ydctg7YxNITUcst68HMmlnOICtNedfOcvotbzodMtEonH
/irR/QQ0KKdQkDxb48uAKe3aV6yc8jT09cFKA33ms4W3eRhc1RbdfwuQu+o1u3oBOf9UyfBsF1qV
n+OTky4WvOXFyxQpq4c1mIv9x2Hnp785xRzmYFo28Zftm2FTqkdTdVL7rgZuK1ddq229gyJ/SpCS
j6sksQTMnPzX36NXvW3hTH7NfcFr57P5sYVsDL8YEsekwBuMe7Ya3nA+wMseDiU4eY0P22Zyu+5C
ucjxWcqHak4Ghm1Njy319I5PAV9zRiBAvEEJsNT+4ajsRD/n+tSikAbt+a8nr6xtZ4fRPkx1WRRu
61oirTAl1LcddATdc7W/48pL7DWyQhCyR8cQs0Dvm+mimZn05HaruuGLT+nLjbQj1FA0YIZwyLkW
6//QHbxbGpUuBd3OozxoZBmeRKqW3cvu7OXNwEAVUoV8QczHqO9m8EqfveFkGwbJyBd68DFzvHjE
2cyPd9EOTiUxMDTGJ2rzSIw4N4bky47Z9lHEdsmf4yQ9sqb62Eb9oFcB54Ei89dVrYAHhtGJE203
P+OpBeNV/7AcL7Tu3G+AcMbY13Jq+SwRAJYOhiD9Vn/5juYnFRAej3KrVfdn2yhR3t8nQEUkXfz/
obsE/Tj8JcPKeHKWLZNZqP69X8bF92Bwpl30+qJpsCO08Ue7uWs7becAYrur/CRLmXROXqFv/mNl
zFRPzqv3rQHbBGlNgM7OmjZ4WqLt27XgL1GlCC5PIVW4ScL0mL7HuLVAjHAN9Vl+/PnIJNxEIVug
UuH2/fTUfgH8Tn2kpmGyiwHIhrgaPg9XC45V3GEonHMhcFM4g5Fzd3yxHt/e2nDAwV62IEMT//V+
v4VLpV0jkLV2w859OyKXMIoR6MmBZW0sD0xxsg/TTyCpnvKhBs5onjKcjsQIMHB22bXM/XsXtlR2
5+aWtC6tzBwDoCLAiL17jlZ+NCYnZWRvry7ZbIlrLyVh8cLKZI+GodxEzTONHCUL9JvcJlJOvZAv
Xqtww0e3pMprSceiL1BVZUGFSXiczW7JowBlZu3/6kqxC/H0yDCyjv8XOa6YbN6Xrl4xI/zBtxsz
Y+HTJmpHF5fu30Of/CANEbDumOc3jDkdAiJVFTZAfZxjFLxn15jztTvw79Ai2Nil/do2fjSYYKIh
Xl3izZpkJn+RjMCNq3LlxkHESmqA61ieqffdIp9y1oKlNnIprqTG5eHFhlqZv3Fo7gdL8sbZdcCi
kwPrBzFt5BqObqz2S6hEtltaZO8q4Fdp0t0DDFR5vz4bxKyysVSeCfVGiNHc3F382ddeNBzzpcDe
/KDfVP3fc12yVOM7i9kFLGL25MqLxBaToyzXyqhEya2HESI1qWoc88Fu7ADioTNXMW6nEWuYyp3N
5c0tHgZlyL8WkizFnb8Wt6uQZsnQRrgTM5Sp9ZKX5u2V9HkBjjoOxJmdK4+uwoq3mlNIaLTdSLPA
84EI5T/+FE+nCr3YAs/Qo4Y+Wq19XB5oQ2tpoVO5siW/AU1WMiLoTz3j+erZSMwmNZn3vs3RlBon
OGwXD6rSp/r/50Dlih4Sa4hiBBF7Xzh+4bU+33TIItSHJD8/1V0LIb6W41GAYQjfVrsoyLy9pERR
EuEduOKOhLHdZSi4IYKqkE+J+ELRLccq5U+NabBAUHNrwsbmOjPlxxz2p+hR1EvYeOqgvgs/0TIy
0KwDXRW1a2SkWzl73jGZxOMSDSoVTtSlqZnA1YPiQexcq/CEBmX8UwUy5KWH+O18niCymqP0AMIp
dKD2bsDm0Q1GlEbkxHNyh4D9H2TDjvIbYLFDxr6eFuvhrZDjVeFDxMLNpKLxPnJkfRfUvyrj3riv
X0oXs8mARWv5+fX0uuXdVITogCwvvE//7RYcggqPGFoN00wMkAaVbhCa2Ag6XlpS5ByJPJ/vqBcz
lZceNbIzNk7rEf7P0LCQ6/xqHYrRnrQrkwmjjhwaC/uzMiDrfUMadkmZ5ySsNuNr58eDHbsd/X+r
GLXm9IItZiYVREXNQckwJXLOEohVcSFdGn2DUuiAG3BeQnTTFTD4QGLAU9+nu6Kyc/gGhWvIuLBr
JiVfCbsb5AbEN2W7YgA1EblfwUCfzGR6rGwKbP/cYi0DBJngCfEbaYO83gN2M3PkRAKyzGijDJoZ
hA+4KjEbdqsxlji3W0x9nyanrJ4p9U0+4bF4s4G2FKK0ly58JX14neJ/GCGIYMFe3G/tG5ecueZu
xQIzVgP3GDqWToizuDZrfD6vnohLtWjsP9u6KjzoL+nIm6wuyyWLS72veXpsuh7OodabiC8ywjKG
YMRyHRq1VvOSpYL61YB4aXPqu4I5GPlkH9tIn2HMbg3LzAipyOrPuu4GDOQc/5r2DyLn6bKcfyJO
AAOy3atnWEWJhnFetwWtxiakW9h0Fad0hZZVGbqBlxm55ROar7DmDtBvtz2aQzhB2xAzzIb2UUhY
LW5SE9eIWFCSCD0Byuf/KXUjNZrAltVjooaWwYeSA3uI9AZKqh4b7l+fWEu59mcM7TM4iUv8KSWX
EGpGIHy8vJRqY6aGU/w5zcSwQOqvzRj8lI19MZqhDwJYjvtyFc5uI1PiLGiQGAgvh+kJUy+8arIu
ah4Kq4uejP2twkZ3kyiy04GmfwaAq5r5w67FSTRBE8c11T8AcKGOHUrSfRSxiztLcnYPit6tnyRL
ZZy1ICx5U1yJTOM0O9oL9ZdaF3m0qVO9EWY9kiR9WeZZ2btCrdOhB8xlwrEhH/XFfOJykLC4BByn
KCiQliIZ/qsAQWMBMR/DWbGHAHBiRW1dhU7u/k1fapQQmKw9RgtUxcpiZAOeJbQJSyMhtzhBSLOM
6BW6PPcB0hzKpHxE87qb50td2eQUXR7c3fPtZ/xs1O+IccRdJ9DHU4ccWMCxqIbb9kW7vIbV7Mvy
zBPTYwqKOh8F7NZmuR6TDOiNMG9OTeUwHVtSU083L30j4XOnlR6La6ToXqMjva6RusV61e4obMkQ
sMIfovfF8KONFNMXkryhJygDB3Q30U/2PIffhMVlT0kzVYExi6cT3ebUd8Z9A9RLc73kT5wFxw8R
uHSuXFm1+gMYZ7PRpX3aIZWo6Q52exF1bgItcca9ho/YNgI1LWhm7ua9dgf8Sl3AFwOBvNo82SmL
Jp51dW0j1BdvTRjKjprG6Se6mOJIOM0DFdz1gpGy80L3en61LeI+Bos66L+onGG/EXSHxOb0YfRA
ebmoDo+EmqOMEBcMs0aV+wJ1mjAwo2aUmd3W0jYRhZ5O9CkyA+EJdmwQPCcKUDyzEoUPIY4GW68C
gbTNT3wPBhelcf3WDKRk2d1YaS2vyXPYJzYxiivRuA2aewMboCtv6JDm7GthIIA7SvHKAjlmRobH
VMzJyTPnNWAdl1op4R5dCUcSZzWYqIVRGxp0G7YkvVgXMxgAq61If/aAmgePA2po/pgW7wgLijuL
9KS+BHnVwNFauvlRDzlS/LxE2SC9myaDUSYGspkYPtrYSTD7oGZDKMzbIsqCZiAnZ5Ae+ACUO3V7
R9OKIGQrR+RzMWUm4qy0LR/ZZ1ocK2IqsjfSWB+i9EJn2fO/ACAaLkNjdPl/gWByptKkTGQaAI0T
+Iusm1D1nQn4Xzo1hF5+XDGKpb7At9sd4arflrDvtEnR6mt37JYP3b2xy8spaV9BAIAKRL7Opy61
QLziWx90mP8aWsWLhArCCej5fGsAWRCM8NPZIRttcnLJdjlSuWHeKVT04dLgw5RLh4XQ1ONeIekf
uJ4Lcss0y6nlIEBsIVc8vn45JV5jMnLe5oBAT643xixkSniTBddQYRB0U0gFo15bQOgWoCV7GhbZ
ov2Wy1DXbvQQYCA4QtnwEKkuqvr2Nj7wto2IFHFT6WSbcHFzrxblDQXLGLLmBbJvjgRkMHzoG8vt
R4H6ljcwbmR6e7LY4PUnC6X6IPBErSoEDNj8gfjrZ+aBZKStCXPNA5HXoHvtEM0/H/hWyjIPpXd5
21u+MJW99P7hBI6K6o5mQo3AGES0Kw2ABX6GlK44IQNn4Vi0lO4SaX9aOO5Pbrwfyqc42LIW9vJ7
2kb8h1JKT0hkuTwSlttXSNrZS1Jpb7MFsXZ6X4UXInR1H6iRWgGvU9v9t6xNdc72c7m38mc7OUWV
sW1Rbl/Ll/e2QyYLO+YivzcfgVI+wLSFjEKZoNOcGDoJ5koiSC74C1WqMxehVlV4Iw/Hp9iNf/Et
CaQD3NNbwlb7+LO7KF46L+z45jcTa4lfi5IfVgJaxfqMuP6e+F0aXZskNEGuYQIsaKCADlOnoIpQ
XNv3+41aGBSnJnK+7zotmKy42j03CsNOTC/TjvSTx8R5weOOGtbcWfDIRw0kYtduemwIY9t73YMU
pgtIax4H1eB3pj7e2/i1c64+7pSjh4bIuuBff1ix/K86Of4+PJ8dudEmxHVEzsVBptCQoFT6zcAh
HjQ3zAvLoUgpDeyKM/cZ5A64keQJ4ImrTaStcVWyGLygSbHseKrewk565ot1mXiRN37apXoS73b5
13zf1pfPjBvOZ1fPC0LCNFUu90WBR5Fmq3Aj/2NqLnI8j+7cuPONWlSAuS7lE4A5Wl6pEDrflaXN
0m//AqPdv3GcHhwNZIQBHa8Z4J8NqvZ/+PJg68cw2BGL9+6nsIH0rkEQ85wrmSLsGHjEUYRGzx1u
DkF0THCl3SCCsXJtahQkS827U7a2O0dN2ayjuZ6NpU8xe1E3B0i7T0qhzva4ErUiqfHZLnlAuHOT
oNlCVG/DWZ68dqPbjc6Bru/7H1JJGBBjRq60edEljzUFIruUMRgxw6WcN2IYG6zLgND+NqyPIZX/
tRILEAzpqujZAewvHfMH+0XPMaSdYkHfR1Q03Dg05HpsSLvQgyX0VHPqd5dlGOiDskxDXM4C071i
l7U5VAVS5pNAptElhE3FSog+41rxmqvW+JEYRTyKfBNNOgGhpNib36RN9c/kl5BPzdD0OUKEWoAR
+8LNFcHwVxO6nrcTU9OvAdoL5gnRkd7xfFW1tChHqMAvrZ+gaM2cytFehlq9XPHedzFG8depm//j
Xdo8UiZLSuC3Jy4elXqLQOs8VX6DaAGgAqaNMAP3j+1qZ6dnln4TeWTXu7bZ8WBG0UiaIgI6qqR1
1I0aBBhTwCEY3tP6xD5TTYnbsiW1GRwRKFSq1lpHQTKRL59+ktcDbHSttFqnjMr3s/gvm0Y+sKEg
nOFCVaOO/WHONqPT3BJPZ9wSWpIbuD4olDg+pCthf3u4LT1W5jlPyF/6yLPBYg327HkX5959Rp65
lmtrshV7h55RjWVP/gYyFN1zKpo2OTTDLSD07UPhGBY5XOvDhwc/Jghp9dTGotUI5CBOXP+4z1MS
tm+JL1g55GsDBKVixqGh7BKp1AolLK8tOjxIzXxyYF8fFwMo0fIW9L0WaNsDTKKgkxRnfroMkH0h
MKe2v+ImV5Ok9JZCI5cbWDIormhdphSMfThOSnCHeJbW6MF+PCGc++zQtgzuArA3Y26wa5V+TIIy
+oW27SPPGiYhdFmQzJ/KFn+RvID+vAi/DDAHjxH7dlA6NPyl1IUlrNR3ev/HVsRMb6yVgqz837td
WpJV0fWnrA18oZPti83xDN2c/XoNXHzZZxmo4Q4nrJK+idBfVO0m1VxBkRuWAWY1v8T/u4iIH+Sr
byOllVrL7hyrZegtLpjfbyGCsetd6/nSkI7BrHfjpI9HMDf1AcFV6H8wUbjozJnJycqLX6hZuzts
XOIpMYxxSOyq7wS3/f6JrRE2h8m3cG/okcjqMOB53Xxqe4/HaN0k9wYrjah10b+vLFK1vHDb52/Q
PMHRRfmDkSi07Tv5uqhI2z4svccycP8zxo3bvKx2AmobK+Qywlqhup2obhP+8xaHYtTOD2cq4Zvo
1V/TwzGPyxnkUQr0n9AZ5E0UOz1EyWstz2hPB9qsQOSqyJa6ub2xchnohtrhk3uTFo3m57CQqjQC
3/zrgk3W9E/KrMdtfG5HU76Hyk1H4oqA5rfevSFudTHAwdQaTaXrXYThtuG2mQyzZrKnf23sjf8a
WXIwCPY7XgGKpEtJAbcIcvbSaTtLuD4YkljonQ9IP+Ii5e1PoOURfnMUcp3LYgWMZPFO/1djw/Yk
ehdtQIMAX4Bu/3xzJwrXqMCBlzwiH8Ad9OVjvYMR3V7ZkO3kxYSYqQ9a8VudX/pvL7STRPVQUdDV
6OwK/F2KsMHmiuBfUY9ccAkjiZBmQXqcjJPbwV8H+EnnELx72LOpgntJqxfGBBHwL7R19UPqDa3k
0B1YUf4WslFZO229eu6bj1tmBKkcgxivkWBDFk1e14+ClWAllmDvB/BPLLr3W46wnm0u1vtL+FIU
0ZImL9nGi/V59Ei1bM8nJ8M+jyAndZXzv7mZ9fnnuraP/CY0thgs5nnNuGKCa2YLjXMlk8/TF9M7
ma5W1vfJqepRtwzwG21XcdS5SGr8mu9cEpByW7iKJHQWfxIJIYescMe6dDVf+/BCKBRCDDewnEgu
9XPWR8nTmtCyGoPBGMYl09Qng26tHYKv9+F+1YjTJvEZxPKnGYFNenCMxcRLdYAfT5pkGyWsRmlV
2c5z6sbw5P5KS64P+RsNlvLORb9w17PjTZ09/YIlRl+NHjz8EWw2kGFyJ+6HK7xdK4kRab2bppIE
jUmX0QnootWpO73uiM6nRTHrWnGfUuvDdavBcckSTznJgDNLF4CPXW+led6pZucjxja3nVhrUOHI
1BE2+ZJN5Q6l8+Q0Sb2nrnrbDq6H0j9LWo6E+wEAVf1z2SF4u7WwVUrzhgm+TE9ta+MJueVzsQtw
uDSyAv626Y+c/R5cJYiXxwEEsa3uWGApePamheYxCt2oBC3sKkmhl3IdzDw4pWnsk7O5FM2HLJDI
lIni36XhNyTc3QOv/y25srHf75bkRXBmfdPs09UjFhJDfc30A5a67XFNwySaQrIPqjwY8F98mpHB
ryJvD/ZA174TcCeDcsUwF51uB3bKkYNe3TF6JsMGkmrlq5oV0yDwMOwD7s1VfkiLpukyfJ76B00V
T9S/0WAui0+F3geY/HWnM+eF2uWDsQ8SzxcoHa/n8ADc5dXoMLlVJavK6mHsVqDck/QYvgILXJk8
WAOlCJKKe9J0m2w+LtsuJdz7DeslVnIYag+SfU4/NYE/GOtAeei4qfYmxeUSnW/ywrXvk7Vszqbs
QiJ9N2b8V6iSOHmXZnLP0hzr4HzMwpPP30BnPvj/IcLKeCoHeo3AJQIqxOiimT90ASP2K4+yCnqE
8NojN198Ptk+GLaIs7hmBgnbRDuUOzAMPFsxHMigZzGetsnyRzYZNkSeYu8CF2QCdyddBHFb/SVz
oNyhcwlOIox8dJ4FrScHI6b9PYLkT7f7L/Hu+wAaHaPyvCHRCyhjM8uGzhdzNHaxFf8yNdxSgWUY
WBC1Us+X8w5SZ605WVilBi65FCA9eZG5SjwlaasuFWTsORqt+bAa1Vw8314yTEsPDyEByzVXC3zq
FTNV5yXDxrLNj+0ZvYvG+iWszgtNDMP/E7vzdkJJakrLVKr2k08jM7th0AtgonKWR/mYiFy0IzZ6
KepT7eTaPIvrPxYGKUP5J1IO0M1adfwJriRt8o0VxGiaygDvFzpNizXAeIsQVUwZV84jRwnWPVLm
vg1VTeWpsqBD+KOOVlA1xq4C2vmNMtw+xvS9/nYOe5qEPpfMdZ+BMzGEKKyvxUwdr9E5r0t4KT34
aaq0TNK3aNwGd9MEcKrl2tLXy1NJPuvLd0qN1Z9ik/tfQyEh38lvJogxN6BwpbB2tZ4f5AzRmlaf
3Y+tygaIZ6edruxXzKeSga446MBhsEMkK2H9s8x+CGuNhxHDWjpYHXCxVxH3MkWn8sayISm5GLzU
eCoYhJ7p0/cc7ZgpswsMSTi1+md/AXcEwVsUt8V2KKuR+3c7gOZZmwkiFFgeoCyYJ9MwitNulSd+
DtCJrZFCIVNZTb2on7zDiakUtE3BqkWVdbqsegloEEF9Unx/mJtHRWb65Nb+4lLUZp2wtT+sdHAb
1ItFgm8MiEn5TXL/3PXCdinLHyPE7UVbHrDm7c5UcT6dOiQOdq/urFowixwHV2MDVi1AK409tGKL
8P3IKTjQC166AY2WoupQoxrDGsgFeSN5mVGE/m8mHZmzIdV10+DotDr2mzDpf4kJXiL8gNd1+PuS
Y/OEhgiqnzXg+GhUp2hKWyZwcGRndlWT93Xq5zTBPC7sumjV545mT+aSJFmusGZOiq7swKogsfEt
vgwfq+u/d+lV6qcalwbI1zPjYTMW44dxNqXCYiulX6PoQZ5QpzBgpQ2Gslb0zj/dFfIaoRK55F0j
ozxtPyiP8AGEplkI4/DDeC7LKvXhuABG2N+sj3++9LicDzrYH3Mu68Ar7ler/Jhe3Y1Cho4wcr/8
VXRsUEUrWFEr3lkwLsBSGFqXUWkVz4tyDSvIMKh+gxhuHbqJ/rcaZeuDFD52gj9BkpF9Xoqcm+e2
1cfgq9bj2vVFfDWsLj4xZS/MeMGBY8cudVFPcow19NLC086U7tIxRqjlqajO/Y+ASTfjd7pUYeYx
4IIyYH+vUag6Uif4rVa1Fc1NRd0bXBuAfxZZo+sXQYPdOS/6rvmgQsbQgXA3ZljBOKCwVQvf9rzj
CSD4++n4SiD1A4IOgEWlIOAVmIomDPaznFzMrE51gPwvD3J8zgsrjiiSad5CAi4F1snK8eohL7F2
F9SaQtDnakutvLXZU7GIjhIgqXc8bSU6d+SsGKyPDlKCxalxHiK8C7OYFuQB4jXSzDIrW+KizGdZ
ia7ruqkVj+472ejcZ0uAf9V9AlOTO4aPaKKT3oMnsC2ysRuFtlt21tStMtfTjCeSyQx1c3NpEWBT
4g2BvSI6IpUM9lhsJyoHK0FIeW8zRgUewENdlPa6YoFdHZxskALgAwBE1tx61Rcq2j6QchKDU1Ga
oBM2QQv69QzSddbHZmNF3Kug/kPSjCTK+r880bjSKav0CzVzNAVq5JDInVAX+vFZH9KEV0B+d143
g1tqAftMgXHTXllhAQnggJSG4JD/pKhc96EcGL+zEl30GzgfH3Cc4vlIcxGeikqqumtGfNaiG2z6
NNavbqQfPkCGv2r6NSYXVs+kYDVMeyZD6J9JZVT+IetmDxWduh2N7sMTz2x57tjzbMcNlyMd74+N
16++8+7NOpZZ5RRQUN3yzPXXc9gp9vYfUcdQ2gVm+jLAtZFYyVMwN8SJ7oLv6DhqTScdYIiVfctZ
oPo5SVc85rfd98HdDwMWf8FKDKZd3dB+uaob2CbpJ1eEzsAWxa/qSLWbb16/Sh4/762k9olRkfCK
S2Au/9Q3bPAXidLXuVWmhaD6LWFcliR2ExpqgXBeSl9bKj0PwyNBuVZF+DMCiuUf3AYTxjETPIoa
n0qRjC3JmMKAzLRcbvwBbC5eVzjJdkDjdGzIOPf3JvZ1dAzlzu9Zh4WuC2QSDusly3tM1WaPBst1
9GLSw3MVQGAVXvd/6uVGGR7LuOdoEuiiPLWxysjZOckyq5eDWmv6+xvcHNrFjxO8ALBD7ds/Elwy
sahPpBiNrV1c3AYwIAi8atfKAxmeYJyaRz8Y04S533NjM8IyxaiPGeJZAdhr0cHDngB99C0coyUd
jhWwSllA4DHW5NSFUBUZgod/IR90yoVhpiUyDYLhuup42N3noY+wmhdHbLgAucygm+kPI/hB3v8y
nwyWg99Yd14GqPYO30+0XjArRKFpJrMiRIPbUkOm0z4JLsJqSYx1lV1wu8d62bU43ozn67/+q9wX
e7uqEUvlS3cU4N/rp6Lx2quFFwr/v2Xm0Z7TaySJV7ZBw/3y+HCxwzhmV7tZz9DmH708bgxG4rc5
NgeGWCzSblgjd/VyajB4j/eSdq5kLurwAMgPoG6Q51tI73xLouy500oO1RGa9VV1kVswgq2+ZEsA
qleBoh/Pwshz6JyBtrZcAdhd7u3tWHDTN238fWGoEu2MPtpFmEsdUOVSMsSiXfmqISI0uWETolFX
ADL9odrR0JpDwdqJR5/gDsmPY35hV68bJQ9v9wOOZjbtB4JH/tmHqDIbqaSlRcr6nQRqwrvUyFBJ
BMmYhrij0QW5fchVrgjnc+jiswJmf/UagDfD8K9mK1HAkQ08W63XsKT9Dc55/ITgZIuEvIk0V4ob
tTrZ1rRBBGjhj+VjyZWZJiZt2cep/MA3JNp9mxrWOgepLBbqyeOO4xB1NdTE6MT12ywlUsnglnbd
gDqQH8XLIill4ZA+XCO7f5ZAIP//ZzZt+9J3ALZeI1VF3vwHfpwFIXlxOCTyEy62I/iW8Np5wTAZ
Op3hF8B/HlIFOODZ/5KqoOm3+vdil9jBCELjJOk4qEfanpMEIDtrUAXax3wXejJXcR8cE08AI/4P
UOFm0i9QGJzUhtxIqN2nvsJMWP/OHXzv9NM0V/0YXFX45dyiMdUSfQBwI5fleez718cYI4Z5awgT
XbBx9vQProBBSIF4bd+xHUDb3YL7c+DIPnKBSOMUJxZwBLD/oQ8NNa3eN6c3X0SQLtRRv+Nzbw0T
SxA17COfM/ytgE6k2xUVK0fUdXxEiK3kQ+s+vHiUZlx3qziDj/B18HA/m2kzYjHL6MOKxURwhkWD
KaF7UtZ4AQz5aLuDh42eSGonIj3B9TKn73cMf95Ni/8vLqBXAIr5X2ht2NAfT4OZ4wdYc0XIUGbb
uhWy/P3z6VzE0JjnQYJT69gLDz4gqNbyc8HAEiVH1OXxtWZHvdojWTKCR0LhXU/YyGbrGqYhVp/D
CllmRRGI3rdo4ZQ4PKfWsVjQQ4Oy+6kgknUt9jDJbMnIBWATjSMsgxUObdb2JWu4qRkX4gNC+xSm
fbuZy1L+k38wsJ7/HkpdNJaRhQGjR2xVXZlzO27TGgOIJbXEDsxE96f8SiYQxYOJO/o/A3l81CEL
Jj4Rsy6g/NNVFW+So1g4dOS20dE7mgNCvy3DpQSZIAM9rphdfWSxFa9LdcaIJ+3Dfnv+8Fs9kxz+
LLrDjTkrecSTSnIrubHiuEWE0wjBqtKIjm+tHHgy0oYg0H1RykKobCvPTH4c1/dVyumf57HctDi3
yDNg5oTlkYGUoGuWetAg7jksT6UVX9gXtBRgFTEGk1hDAIPBGqmWw+itfVJIHyLwd3ZLWPZE7+7F
fjFaDuMbQhKCj8/e7mCFI5I3PLU9ZVcR3k6Ma1bbUdvSoyxEQFsOLGk1rycIB3T5ZGa8bMrImz5I
TEUcrPIgMsQMcX9w4uqp1I48tKbAoYm04JTL5+6Qz33T6R1eTipfmz1Kqy8QJa/vlDmoQ0k78Bzo
iEIxTelMjLL/aQ1IPWz2HEZr4O78+7W3PJfooVi0T5x1nJw277p1V2+YHDL8LGEh+yWDwzFeYYmM
+4vX0Bpgp3iiIbBnbMzUrF6fkGhW0o/37jkR1L/2TsCUNMDF+LqWaAtpdRaPD2kmOYH+ZXpJf1+/
BJB3bAE1QoL0iX5M4RYL+SHBQ431k6WFT007OuHf04LszzrtQPVsO38BJzbEEHyVXb9KM8rhYEav
b8cFi/vSGm0n5d4NL9NUVX+URirFDXWCNsCo/libI9p0OQ97Yk3dGUmYyLVZ9+Y/LPa+VI9VdCdJ
clFo8sdpX0ZRAg2c2ZY7qgLFRhCPpqRQs413ls9OGVOo4/EgCAVz+A3vfK3yy5GfLCtWH9IE4AWG
Ak6UkmK5El8IkvodbMgjctq3uMnT23YEbfUyjmadgAMqMwgX/YoxA+tP6nRVkKDE8oiLpEBVK/y4
XLajfugTtXKsnK5uQAC7z0yhAvzLQ9KF9nmHvMa2SkP60jDr+6Q+GrGvQlAmyZzn30ifjTxns8M1
gCHwWQdyxHJeYbPbksWz9JdAlGYzPCz1XTa8DunErCJeGuliP72vqdX7/FVE+WSabN1K4wpER9JC
OaUYlmf/19mHJHeGbQyQ/oqfbsBVKheS/CCKuIAz6S+StcEKFAekgeg3f6RUgosp4YUdCL5aEHol
gr9ScC7rLPzw19t92qEnuM/0AFcQemHcU4pzrHU8wIG9MXcQO03fqK91MWeSz8o6iD4eCT4mM0yd
EQG1+2de4L6sMdWDRcWVifeHkKGBbMyeTN8q81FFNhX/ZDI3jjTOsGnluUbpi5sYio8RpFqezTdk
WzP2j1DLtqIBb5VAcJQVUJdYSydU4bE1eZGrwltSYpD/R3EH74pL+4C5xTqG7aCnkxIgNLgJ1Ucc
XcOA4YSJSZGGMhOzhAngsODV7u9v51rG8++jnMgt4xo1dkkuoF6f0a6b9KeTyDIDw9u41gq9cUpM
XQoe+16vM2tLWcMZ4DyTm4q/vaXKri8K1YtnV2qrw+4ozYHjWeKe84juKXX0UQj1E3AaM11gyJIE
xbSh3gM8y8XP3AG8pi0h3+RJJELuUENMg1NKQba8gqgZ6BvLxb1kvEAet32b7ufGm1OHXj7MYEDk
nMkNY/xFDpQElUUgvjP7RCNEd7YnPvhqAs1hkFbL6tskg6HKAIlDOvj2bC4MGwQtAmos00d1Q4YF
hlnZrLcDI7HTYegPYO42LNzLAhhgONbOTb/O/mO2Yo/3u3+IpgBSAp9CraMoAsxDX+/pcFEZ2KCc
GEZdFC7bDzQ4Hf7fXXi0fK9WjMa/GD9Oy4i9EpWvhw4r+XWi6imamEqzaUqRZA+qkCqe7uC/Vtd4
PV1NrECPBRoWMwbnOaIKpSRLW2g87xm8Kx+RlSdR+1QEbzs+HTTZIVWEDYJf3qlQyYX8/q4iuKoe
/uMk19B5vQACLbbUxdqKTHO3+7xGyFpWbQWpvr4dE66FU1Dkncwk7Cv8aWt4gY4ks76tADio94M2
xDyL87t5fJ9X3PO2UiKdfx4uMm3mpQKg7bt1nSPg5NVk6s7epVYQIj3mfRXqJbhg3cRsH8sniYzJ
mMC/gRHFSYDcMyVuXAzTAA3gIHwDb5CWKWFShU3qX6Hn1A4yKL/S2baJMz8FepG710QsHmwZcnAo
xSuiGAjIFdSB76KQVn+0H7HV8mApU8oRnPYtQMeM+ltqjNU7/aa/eEEdIbrWROlFvC3Pobbgnfcg
kNq9/wVJEuZmqguUPzWkyHOybojjJGI0KyEa9rTS1+Zp2XWGv9l5nVa6t3vbQuxWvhHQQzB78fAK
R2fJaZw5CzjHEbAJFZCBZRD5nOtDBRY3Y4WDuAtgrG7WAr5jxGMrUsacRBiZNljKgKsyU96cQ71G
Z4P1547ywRjbuL+7nqGUTcla32tMoWYu3OZp/5/vYfBeHVLpv0V3lRg8hQc/+PPnqHBJJlVwWkZP
rA6asjJcRK7PX5M4CCgGcgQLl8D9S/iNHp2//vIUsd/i/YhWX3nmStTObk7k4+vQPnqQ/tGr4WvB
54SuvTfvgq0iPYbBilC1dXfUuCzCENDBLMt/n7zoO3uWpoORhX9IpRTKv2ESBheYAgjS0ZmW3MhJ
zoXbmXsRGcWWyl+xD/QvQvjDdVFGAhzH/WQEHOzQHCn5DRgJVWVyX6lsNgJx8a/e/jNwrGFk/0BZ
EgdFqq0JlaIj9bvYhIs88jdUHQ4J3AvtjKdXVaIlf54OcsFqWCkHawjzkpByviuHMknFsof0RN6l
Iv9Z/wAmAhT3Ry/bNbICZwH81qlUHpn9abNe6dlQAPc/sgJ/a+Z3+HLU50QRgQuPsQCLpbBT03JQ
qA9AfHlPF3jiw1RWKuX3Z9cejLkwMZQg51PuVTInJ/s67upOMYcKKNjNMcOgczKETak3xphb1paK
AGezSZ8v+jePTUa8hcy//VCeg1lRcSwd0E19oT/0Ns0EE9f29iF7GvScgwLl7TNdP0VakLOvoTiK
TvRQWw/MW+NyxgEttshyOMeHdFGy5L8/eRC417xEY7vQYwmpRDFVpHVE6QrnCLEgu4EpM80cGK/C
htzkyGez3u4O7vnDcR8IzOmEjw5nYTO2156HZStj9gOlrDwZQikQMO3c4gV0sgQg3XlTdm0wPRUZ
cY7McYAvCjwGW1pgzDJ+Gwmncpkf0L61NG1OdkXL5kOCaXBY4BGZnOgZNGVe3sI6OdJZ3AL9sks8
+hJWNuMxwZbl2/Ph9NpDpenP2N3PhGsay7QPu2s1KOKYLwCk2JPsaM2FdQ3s8NnpEJX4r0V/IEgT
wqND/0+2vTvmC/0YoO7qwPuhZHtOv8M7aPMh/VGs/JsAufkk+orzl+yB3mvTrkDSiOchsp/ppVoD
pIYmCHyjayGJ8ZT1d0cKdEsuTruer/Me/kbpuzWWEg8QJjuXlsj+jXQkWcUZ9HT+YLi51sUvY5sU
4P30Ymcn0obEJWFoEejnK7FhYoHrFt8x89NEB1ejuZYPIQRZwpbl5HTxO/PnkBd55Xv8Thc97kpl
YG7VZpT/+5IEAiKmS0rM6S82UqnywkZ8+xjq904O+BMm7HHtds7h5eVdNt9pTwwQoKcryIlt/bOq
7akaY3bSGKSM8rZSF6G+Vekdmyv+rAQFDno9vv8TEcNNwFXmlztWxmRlsD1MctZpTxFH2VNHU055
+L47DFzCZ4Q9P2M0acfCnUkQXlNcaxU0+BzSUxZH83XXhpLB2sozSnNY/IP9VF0oBzYCu6ds5MA4
XsyhdhLc28SgheHHmOkDkkuKApOLu4pgE+DtrNS2jQCduOIA0tAmcdVuW7vvtTSkkH9ExFfolb6j
FGWU022Eo4zVir5rEjQb2MCBRl5DMXGxme8ouk7nCkrAWAqTG0LfM4YhhnmVCQ99wEOjUEhjlu+g
ZYNT2IR+ReK12yYZHPcRS9t6D2Q9tUr4QHv1+eob0MOcRM/nzTgy4e0SZvXWds7X9k+aSjbmxVX8
HzofG8qgKqTTKhbRf5YOH5SCcGCzD+NatbPPyWHoIElTolLnWoSDfXvTzHkBDSgxmmhcvk+a3+UD
k+0g6OfeIojVOFaRKYCSm6JxqfNnRfF4RHRZIpo5zT4I/yo0VLS2Fq906bLcPHhRNVf0RWsviWvO
vsS9P0scoz/CFGpLLTrH2w42o/J+hzZXHC7JSAiPAXD0NP2TAhPDhgzowCIusFWTJpZyi7NrB/Vb
3DWNZemt6pgbKzB4J16NC6oiqz2posy7HjUTMDeG6lZWQVosse0ChvFKYk34f9GB7tFnTPCiSgxk
vfKaTOVC12nh/BLRY4d42ICBqlsbwXAtBIHjcFaP4vMIblxPgHsxUc8mRUhrXxn2Js0ufykocZnH
iHmbWVT/zaorASLmtA65nXadl6OgcqYMpd/02ATwtL31TbjvJ5a+WoVbp8KT0tT4prUorex+U8pd
iHxup3hK1otMxiLw6b6yj9abiRATWrjgv/M+91GOuiqTpaTM/75NIrsn4sCKuBxfIJB4r2qmV9b+
RmlbTlKi7krqAk3nYh1q6Ov9H92HiB3poTsEVpZpbx/SIC/8SgEgAngue4CMpZJQGTTrs1ddz9GK
ur5tyYj/IqqjMJt35GmPY1bPnj8w83qv0C4YHaZpO+VS/39dYUpskMoUL+9zvrqQmT1PlkNNFBgh
9ZgcTWX9IcJ9hXKNP7vlok2op0k0kdKDZ4JMg6vJyic73d6FGLx3STN+aV0sXUKjjsHK74O9Ak0U
algBeLgEaKM29GLsG7bnmmqoskxvPHJFKuWIus0nT392sbuHvXv6gAMF0IEaY0W2Ny+vs7KSNLWG
6Sf0LcJpT0cwVGH6xXUmIk5i20JlRSvZ1pz/SDbIHTCXmyw6O0hlfzlSV+pmGMvgh58WGSUVcBNt
spbwSWfpZuGZFu+oxOZTUBDMa7PkRjEr1LZSSJgLqJgC9ctON8SgviUn69FAHBcDuf2pj1NW/OmH
jk7Hg30Fodfs0H/UK+7sdUAEuPk/3sfL81Y0KffxQSNfuuL3ojk0+FDNVFfezEQFhpJOJq2Uaks3
QlNIf0L1r9Vl6XQ74LSK9UtSzx9YCT6QI5+pLl7JJYFO8BwXwP22TuRHOln1cOCmT+aFrSB+sc87
kf6UEaKPDAK3BHKTE9KJlnJm0dbns0sCz8hdna5G1S+Esu2iBR1M6sfU0i1IFiOsckOlbpElP5nI
E5f4ztoTnQW02r4/lMIuIkF/oh78Q8xb2EFXiXADXZhKWKh70ue6leRUMofNkVFpCyN4Ri/VuF7G
4zeaHaSsB1omyAOJ49JT3UQemgINYau3uiFZHbakd3m9uXA08baaMlHLIj6s5N42cIqwMSMMd3Xw
jylcpCkam1zv313hgRc1GxyQlc2CcA4ieUKShtaPeamSH36nxVYGOduPhRpE7lf5ZT3Ujqla5wJa
QSrFo4WWDmoewLJoFBiE+xknOPZT25Lklp+QUt30ZhH3qsSyVZrZU0kbv7W2XcdhkAoTVdcbdPYe
igzUVmbj2fK4k3t1N4mg/M7o6ZFYHWUXHAK4RiiBHgXAWyOhqTUwPImbAJtNr8yd5Qyivty6iQxw
Bn2WCjjXcP5rrs1yIVCycAu95xtX55FiDGC7Mdbs61MD0ggIUzMXz1SAPQKw78KJUMwmIqqzM5xW
jZTywdH0ru/sgZajSSNKnb393TXWGUp62R2WUsOtctznthM1//eaM95uVwGU13NLyUZpWpQylL/u
ABKh7/jgciBTgPV5PYrzzFWTFFD6p4wJpn+NHgXTgOcerf5x5QzDjU0DFGt+t4jIkBEzHbW+o3B9
Y1LaXXDyKTFq0vorky1r2bSLE8yrHOZ7FN+ryoNvTjtyT/ihywtbYsh+xaAy66/Hv3g255yNzXgC
aQeIURpAK3gdHMxTeo8KKuI6O7VRskUApfS3gFt0WNcqWuIORt4ucFB9Qq7O/9k7iTJxi4CjpWlI
pRTc7/U4H3P8F66RNPoMTJ3uxmcoajlL5cPaMHf6UD4sQPyQ9Co+rtzjdXzijnn4TdhvK/haQBXm
GTlF5j7KWDqLCPWwp1xnrAfjzYOkRXhrUiVLtkX7t/Nh9zP0stiHvdOp+whsszV2Svj1fJcivCcJ
iJWl7mW9BtF6J+005R42tzJm0eKiN09BcQstBNJtmdJA0SsJvoMLkLwgOhZ9H0QoPiv6w09o5vUS
ixTqm0YOdbaCI5KUKQVpnINcftC7LaPm4nzqibBp00VEDOICmxlF+ALrJZySr2cx6yHS5tvbXKZc
/QvaujnPz0G7hEBD8iEdaNfRSv0P/SLLhvmash06oK/rDy5pFZsKYRgfzOh8SBvnFq44GLTRCvL/
sCrlXhjjCchceE8yCb+CeeYKh45xii/gJggt9XFZG3G/eEURxDmbmcvxmBbnVclXUs5VslhlqlQh
AjJln2M4bd1BXImdZsSaemyP9Y7gBsiM0MzCC+jqTUWoVIEfQZ/sxO2ufodjODAJ7O/UcYkm50Y1
rTzGe/f63DsAy13bX4on13G9Q6uvhTJeDWGrzms4u2CmRCkvKMrNUbTF4LTF48CwIv2uXZG04R4f
Ve88ORXzzQ2cxGdMkP2z+1GYucnDcDfEQy0S+3wp7TkzdqJylCilrJTB6ATkqrRJ6fi1O15zCEor
xO4nVEBL+1PJhs+YWLkiOPhwvaipwWuUr7wj5w0YbG0nZrNg1s5PWADJKeLqry93MbDp8dr+NJNR
jgI8sB6mqed3EnkVN+BYNq5Jsy/ZcYNWr15Uw1hGudxYmJgyJyveAEhW3lYh3UUmxztBipli7zVH
GRQ4gwXIF/JE2fdZrprhUdG2xJyLUki4iMZw+Yigc+fIWLr1K+AFRQ6h0olzZVgdwdpbBX4SPQVv
HApfNU9eHUgOhZhnVbmUPW5jgSYvtxWNeHlR4PLQNoY1GK1obVkQNhUkLkLRmH+1pPzUqJX5vrFc
xUi1qVrwV2wBUpgkiL7sAw3x/rtvjfOu5WqkgtcsQl6BGUXgraoJNo0V5YKeDG+mN3OfWOQ8brm8
xXs8O7P3bEigxq6OqgILn6G0UG3GBVgwsiB4wIKn4rd4qTPGqC4RJ+HNyRY20S7ktkja53wmRZfx
8TOeev4eDQA8OlFGNiiuoZLANvoQRgWT0yEhaV0EVR8uY8BvGHl9+K972uRZ68/Yqs1EvRp52qTh
I1ISUklWDWgsGYsqzG3Adr7QKp0fU9U3m2tAngQGowSWuVq35aGluNIINFuz/enBOAXXXDQR5IEW
YjhfGQWXrNZXap3/efjdyHB2jezGGp0C6yhnZdQ+8Bn1880qnFJTgwGmj5Lo7xNf/MBc2PZ+1GLs
E+4ZWP/XQ8hQgHI4EJ/xjay5JLxotDCS5A5Nebqkb+R1We0PWYBUDGe/W+tHZAxbee/HjtymbX1x
cI193cDmjbN+1kSWKccSL7FES9hSzINUy80SkJ859AHaNSL1mEOJW+REtjAP99guSKkQaZDoXeNx
DypS7nGNPju7WO5DzGBfsaxbaGGgHdKRfax8+5OLve9cyli8q4fUnwCFBnqfZ4/f8h2BcN5XEs75
TccGR5/7q+RhO1yAYIVz0qji2h6bU9t/hi0Xd6jDUF8mR/N0xz+j/b9uGX62+LKwF5G9nEpVQvMf
B9KTxn8vcYu0my4E2+6Q/AaPnPywDhuystyzLW+6B/O1RVDUkGndmTj6sgST5pm4DWZNQl4JtLG6
/gs9zuqqAt2X0fQMNAG7+MisfID5faKLeWberm9fphZeMuUg+cWd+0pNV+z3snB6IkXRRQdnHPMs
VGTQ37IvEL7/ViBf1bEG/JNsQn7s4dNazZwBrZV2qn+rGdAUbLcuRcxdG3z+fMVxFsax24Vm+MBH
fEmSPdCcnmd8vTb5/MBoW1V5Y4L1kY1KBKWmFaEXovYKl4opp9N6VXyxWUUXXzlXANYzLBKRmvyk
Yg8QZT5EBAlA0SqvwZvPWwh7bsO6S8UQgSVzq/NY/r5ZAbps+mU8zjVeoqztuPUXkIOCazyzT+Xd
zBCPgmnVUYBZJLM8LIW1VnkzsWeuJGkP7Br2dn6NrXCQSaw+Ku6/dA3pAUZ7PiqUq0DpbrZ7byxf
ZKk/EKNfYmL0EX1Ix173eqZekVHCDJoKI+4Ijj1wx8ruu81UgXsLiuleqIHQPNJj3+a6iKjRqWjU
bMyDDkzn+CnbjRKgDZVrfF7fw1xw54OsQ0uFmUYFw9DJDvRsVk1srD4l5dzKaYaxMdv3y2q9pyuO
2IeI8CFwsArhVbvEG5G43FItEMEolI8c9a34T69pD8sF0/DqJKNrpvA1Nz22xAO1qOj+jI+DVvHY
WnUmVEKYTLw5d4qQwfEmhfiEAT3i1YgOrDAOSpRfQAzmazHsh1bsf0E1R0WGJI1AUKtL7LRRE3mn
vY8braGUxAi4HpDn3VaJ8NQjzG/nRIezhqpERH8O0MmY8ZTVmCcPDRMCvGBEttLh/m+m63CKwI52
sQc/InD+MCqxcu4C817HjaeeqfhnV4QRMqvGbHM9P8coikHmxd81aBMPFklkg1zuUDO1zGso3Atx
hIeBPDNv4239KyyfZbVMtvyM/8OizeYu1/JBuIuIhAa7WGwkOG8tIO/3NxZBvcowOmbbhhnIqOtC
Cn6JaOAQ48mXZYm2SIQ+emneBRPyP2HENNclrc+cECwLgjQ09ekl9KwQVxKp8VZGKWOiY5mt8C2u
/J0XKtHaIc8hNljUISp5f0h260mfdW3zUQ29GgmFEi7E74ldLYXCFP/Jows+LXql/dLQ91gAPaGI
jLqmxpFYeBguPZf2CNjb9T8Dol3TrhM5LUTfzMQlvExzSX75T7+LnPMO2RgyiOcHzFgHFpI5POJB
BvMgLvQ9fFgbUIEvXVUnIQ+a2AD16o/QMKp1LawQ42HdXmRXXzUMVkQqiAR+jhnfJippLn9RCjri
Peg7yzY41/dWh8fj+Xv5RnACJOen425sPqLmIeQoDjElbgjJxJFL8vYlyqol1l8UIj4KFuENs0Nl
sEyPHlZFx7eTy5eae99dMCHjEapCSI7+VK9RJ00/BYFvzyB8zvbKjIrS2RDqdF7NcZ9DbpjdhcmT
5685/YnLHhsVLDzM+s/kiHviGvKhaGxL07VX0dm+om7bmSo4SJwjUQlnuwZpmxxpxEgPmC2AEBid
z78V9eGblLIsibZl2wWTljsiN1sJu2welWGYIDnvXTfteGa7sSjEboLAX6NAdaWPwbkBguZfs6L5
i5dmI8jcjBMpu8yGKkpYTrwbzVtlprAd3ovEokRYCs6QdaiczXj8JXXeICwX1cCYIUjsE2kkWARk
0RGUCIvHgu0Su69WFZNoIs5PQGcX+smt8+VVbsBZ3niwUxDg5197KBeUb8x3Ht+nJbXD3UKGqRnz
CBr4XUuqtPiPb5L3ZAYyWFfqZcPDnMlUQt5N6NHGdpbhgirqT6CM7LVz/cbZY8BT3Nk0nKphitTG
u4bEpIO5x5QcLPXG68dgTGyNL6msjDyD3ILfetqThHR3pMptNfFkSQSr7S3gS5XE2/tRETSaAPHO
kJyULFrHZhhb7j12JrjIRRYIMQ2nTbLMKPKtuoKnnqm1Qo3mlfJSictLZS9/RtYZDa8MmCKVDmEx
T8PmiNhMbTd5rrzVqnPsLx7O1RFmfkbtcmqiFm+hzwxknv9zU7OyQoMiRpdoqnknHLaCpWJZlKN+
lKvxA6CTmBXIf00lU3sr1JXrKND3L79s5JM24iUi/3m23i1pVXxW4NDKvRFTNBCDdDaZ7EmaAzaR
mjHQZl9JC5/rsOsXx5E5TUWzjXLppVXlrFN0gDxjyYkx1C/0HTShKCqvxTN8KIIpw90Xvx685npD
2yjl6552nP5UBSOwR2UOsjG9OhuOiZu2BtARN2rJqvRMi6MEghhDBjqOAMR+fKWoh4CYok3YL0/k
93WhM3wMIVUuEvEn4/W7SSY5WRhZHoc0Mp3cCMaHXPJ1Kxd1LWR/SpSdl2swgD28plXYrqSarfGP
to4hOS3iGqD1exBP6t6jwzbNh5SHG9i1NwS9CTcSkWHoar4j5e+ImY7liVhGNalSfjPNuhxHSBcK
9VKffeNYiXOnAq0kpMJb2xdqoACpbx250R5F04PdXgCrIjzbzvJj1FvS+a1Q3odHAVaD7xpf2M/v
/XZmFaWv564SkQc2BkQ93H0+BpYnfcSAq6IlbWD5NvcFnO3lyubKpEqzY2LbjEkzEiBrKRFBuNrm
MIhYycyz+2MDi05N5ub0ZM7j5tGGWU3ZQa/+hUFzYUPh0ovgiNogfD8HhgEEdXvKU8iYC0EjjFqC
eAE9p0rrB2oUmMVNktUhUPjrG/SMehytrqProIu+QqSFvZyKoQyTAB9iDK9v0IhHMffE+Xknnqcv
NeyLMUpSTpS3FHT29DY82jBFGxF2c/ROkKusdYQE+/k3WYv+lfc01OrAD9LOhBzoYJjVIoZ690v2
acZq9hsJww6qRFzgst/PyeyKwntmDcA+LCJs1U8laqf/kl9PHDkOQDtBX/MdSS7MjFyd46GxJPhn
h23fVL5zHMBMQbmBmi2xU5bA2AX0fad5V5Vn1VysBCXH6W6lThPIqvG8EBdyziHt8L/jr5eAhXk+
rSw8INAcxgDmTCcwv/ee25jN331m+LAZQu2PREnHiy58XS9tc+Z+ko/ngZiCHIXPfnlfOyYhDa0Z
u1TJH/IMmDAqaAUSpT4NsCBPWfp3VmtaI2UbpimmGQWTa/TxLWU3ckFSkIIL/MOOJZQk0n0K0u7V
MVWEzEMaVvetmsWTZI61BgkpC5K1oSCdADGsrjlf8MH3s0jFNpdyZXKDZMKcn/shkb/pHt4TJQi9
Y9UN6R2s2z8UTx437q6mWzs7GNts9aoNDT+1IYoX0ik3sn9YfKpxaCPsALodlDv1WKvf+DLo3wFU
xP0zWE1caX1c/IY67q2zjYQ7ftAkirfeJfpn/yESHlo2nzCnbbZ8oap4px/7OOhb7gzVAfTcojpn
2XuUjr1a07c+Od/+R+tS3RWLeMG5lNCnKTUWgte/7AGkQ/0MSsTWj8DnJG/OcqUUyMXY7IMbWMl0
mFLcjyCR4s99RCbBRgJKxRpz09z+NnU74Sb6QGHylrF2HDKpICkV88kLAi/3ZTj8Qrz3+hrx9XT/
RxqMshi9RaZT4A+E2a+nq8WljiJ7gsdhtq4sztR/w6S0vqt+bIjMDE0M6Eiyi322bQmlHtS3bPTp
wI+QGCCx3c39QJG9Fx7Otku6qCwHsH4xdFpBM9HHS4nP07jH76vuWGlew3UF4KzBTvxW76jlO7fz
MMQX/NDkOBppOLLM/4gmpluBGGO3tPoC1bVkoGrPl9OlefDyC4CnRjZKWbCuPG1IIljTuG/BLxtw
+AXBEtPZV3I6bmhT5Lp6vAvgPpGgR0d+h/E/BOI8TWSGjg0wRiMqAR5j4I1hN0Fyi/dDmlHRWC1l
Kw9YwA+pXDS+Qj7IqdHm9OJTaZ0Xn4hTqd8GZaq3k47S1aVcAgo/0fhl14TV4iuadFaRPcP2GZ53
5e5Hr6HZys3+HMBPhgzCobn3SWSqN2sT4c0FS3SrBD3W/WAXSw7WAue499V2oy+v//4tzxTSrYhl
LgCiikaf9UcRG9SIntEOvHwUsdPFCBcaDNg6nSQHQFJwJ9alf5oozlQ/s9Vc1AQKRArAzYb7uGzR
XlcQvhExJT+OWyoUsQHwsa1sTs+P5nVex+2r/uBVQ7vonOleo6/cb5dxSoKBAqNXQ2u6/X91kki5
nPPb4PAIObEmVHzN3p5NGic5hfNFLbUovA7TzBkhZ5cSX7jUxX5T5g0PRudlyUDwGH2KaxMJKInA
f20xkFmM03jLWtAeP2ZuASHUOjTn9aBatFEpmIMzsPomyGf6h32ZakVKRnA+EjeBMT444rsWxg+Y
NShDL1a2PnaHxV7ikGZyg7U+MlFdkhOV7b/zutdddv/4ZK0HyCgWot0ZwyIzL63Yk2eSyw97SwCc
HEoWq2DKcyFuDJg5HfabdTRIIuSrAsnmDMzJ9EY6BdCcGArjoVah3SheBHpbz7xnzqlj3TzQJibl
VPijrb7fzqApiaLrlwk2SUq0GZepbsdN9FqGAR4FjyXL0E6hUSSLCoHH3yBqdz9ZTVTCTVs8zleC
/IHDMzwbKdx85mY9+edEfjtf3gR1yxxQd0AHgB+vgFSVYKafo4XuPI5VQl7vTLyMvLHphaT110lD
cXWf7QL8FYVVGp/ovN2NKuneMyIB/QJq9sdTQFzbIqEG67nCmPf92CNwo1O6mR2ahhDuqegFo/x7
e9SgJ2kI65dPweMri7+8WwUvG/iwzWGgPIyGdiUtBXM5jOqxv09kwvCQg0vb0UBqrg/XWaYw4mFM
ADlqj8s+fC4vmi1rfO5RBHX/C7Zie84HpB1BAu859anVWMUM8+9IALhBLpaLwUFCRJ46n/FvtAlU
SlvxKm2cDtOnkEK3jCZjqaqg1YA4LjxzYXHV/WzNLzX3s+m6OeyI26VaDez7+AWx1C8K89bXuOf8
Vnyj2mK9NznF/bZEMH9tbI9JVKKYtsIpAx0W84rrn8NqJP6VTE+TGClVxYyS1B1Pryo9EwaEShu4
OnNYNl78mUS39Z1TDXyBL3uCS+7cpJXiRHxYXRIgLEkt2/1p5UCKNzgVkoJRq1rKY0Zvyt48rEZ6
hiT5412qbEO/xVYCzAYIb9+UqSi+1KlOwYHmZyaqI7ZdtW5h7Aj/4NKGKiert8Z0R42w98Qgiwh8
gvWZTdHzKV0xOKcO8yd853G2GBHmgqCI8mURJwdzy3W6BfmVIp3wH/PXDKkFR1uIDl+za0sq95Ze
9iC4nyedVmYsHxQeLCyIS0b3lp528HbIvNqx/aI1zbgxtI7PZ/vb9WCv2Vl+y4rLbFZJXtXIsDop
GV8H401W1EAe9yHYmODiulQyd0LKB4f+JdloGX5X9vhr6j2HwhlRQW5hy3pVw/8m82s+vgoilCQP
QWITAOQFgQEvbQTWs2u78jwwwPUko3JDQGW2ZivLLTSXO8lrccgvINRZRZ9rajbYOf8fmdqyoy2z
4sqBP3sw2FcE+458Iz9CNtJhaHEUc/jh6SzkjRi685LF4J386+sH9som4jGopjRMIIAhUbcJDe9D
/oVaPDl9E7gx6kjYYVrGxd7coIAlE0T1qh/uj6HiAuXTV/KwSmK/dQtEjOHLw92Z3IkDTebYCSEd
d6dR2phWOQyEXynJ2r5oibvEeZuoVmSaokO3WrErtr1FcmfIFZ+sKxH9GKijMJ1YeKK/hESJ9spY
5FAl8kiBwgkMl7REHHykky6Bf/zD7jfZ/UPVrkUyQjl4C6GqyCwfCCfsrLEM4caev57Q/KczjW+O
Vqvm3LqUzPM0lbToHcYaEiNtl0OZOwNZAlulScyPK25J1eqvN5cD6wNurRv+yw6q/PhdeYljLF79
oTeWGupPrP6z2iizXOBZdOO/dt4HnQNBomRYil4cizY+ruOeHMcQOvSavUW5v3GXXhnFlpG/MAuF
wENy1iYKSMFX6fg5SmEnFsuiOnsjni4/Giskhw/OMDW3rxKOHmC4Iz+lD0HZ5n4+5E9KBxbz9nKk
WpJGJn5MGMbrsk7ZhfWoS4SUk4mtCiOAHzYMmJ+Yf13bBelpbcEjFsDPTRgOa5DkjzoLKA9V1+Xn
ZEBpv9/zxO23vIGiRbzwNJbmot/AdphLsxB9pGUYE8SUHvKvQb45DKlFOmr6PJvRskFEj2cwwLwo
J/Fn1UgkRJ+1wSqT0vTPNyFDGmoW/D7mvBAX+baVxquIaYnmdUF52FqkduPVSQ7w6+EMLoGIAQUq
o3MNGgavLrZniAGfyJ1cvLgOdNMO7mO+Puhj798bcX65LkAKpF4WCavZzD8lgPfaBjn0kuTcZMbL
TaTeCYkt59DK8yUx7cUe2jI6h8fLh+sQQkDL9S6gccxffsUUhegiYJ0lAkTxgKTxleV96aE5FIEt
9GmfDUWMsWQvVmv9R/ovQMoqq9KTnpOV9eloX5Gcj/gZn25qi+vo/1L31JzjpvQsCYixeje4w17g
s+rQyClY2QtDPwn3g+aIbNOY9cnfKBRgqtsVeg1pIdA+o3OVBphYRTKmRdo5h5Eq0zJ7NkN0ed+9
uYdyqn+lmfVLOzCS8FwwgW3aGIsCmGrsAo/DTtBrLqeK9wJk4wEh/k2Xdql92kycddM/zmwBOM7X
r8EQ+IVrLoWutWqbJm+JfzVebqf2Qe+Obs38UBcHGm+Sr4k/63diTw53yvzcvFhXy13cbvpZqixm
YKeOSDJXpzwWbSF9jl7nHZwAtbKXhhxGpIItwmu6gbNP7gB+FzNsF+fNOI4ILV+i0501bak43dFP
MC3m9rPiRigpnen+JGSAmLiQwYf38+ASrrztPnXTQRS6KhGCMpRiefIJXfO59unxsQAPQ4H+Dl9K
//1x353hLlGmYd4zPR8pw/zPKlcRzM7JMsX5idFJvEcuTibN4Vj0m2iPcSr+EfYtnwKFteKdMmab
llKEg3QAIRLDLM2+nkNhHsWyTDBC0ZNvWz/saDWMm/1llqW7nupkmB5O9KAg0gHOINMwVJSsGIUE
Eb8jwj21KGdK27/sbYMX5vkcTlDgTiB++lcxiWpxebDwyNWLUGPOfPwG4IvbkDCnepyoW7IboZlS
yTznSFb0387o6BVX/MeuXqflnFqKUy0vwXhJfVq2p80QwYA8erooIOKb5UFQ01lGTODndz7gsI5C
JoDkdsxnK8lvUolS2NlAjqfdjb2HT8d5MNTJFk7umOPzlIXE+BZk/rCnN11BxYTSv+c87pBefddh
3TfVTcCByDhNSCQa7IpYj8MAxTLDKQQH5ZX84SL0FvTEUBbg2Caq0Wr75F+tRIl81FKE0Thj4L40
Lm14VusSVnRiAedOTiSWEO3dQrdAiyqB6HLstmLzarNLvMFCqok9W1HfLHbBxoav4dbCSpBA1f6H
MfLEdK3qs+h2lapb+Odk/t3xWmEFshVNs+OFBX1zS/WIYQjmLr0xxNS4S96ENSabh6GsFiFNylTc
3cWXGby9u4do3r2OM1ujk41mAZFvd1p+Te2g0DK6xUtHD2JnB5Z5cUShgL2HO+Ow82zST+tmc4Ba
CGzUvYwE6UBqA+mm8MZf0nHCSOsrgcxND34tdIkuR/ao6iAJ72fW3x6zjbncFIC2zjqmY18QAxd7
TJNyyN8c5m4Pc9BoidwtsS2lNlS5QqmxfoWYc+UUBJFRWoow6WeC1y9UpZu+YDVQNh6fo2/TSYQU
wx+c/eqFSe1/HFTvQno5Uahu+2JalAiOSoA5NLAwu8NypplD/teWsS5y43RTJ9W5aum/vhpQFfh2
UsdQbxasU66zAjRG7socPZEysagjqC4xjeKH2QwMt3FWSlz3bn4j1MN3BhWuvNoQKuNMdB8gR2fH
aEJcCBmMHF6mz4oUSDayHskFMoVRa2kHwYJ641S+vsbR2XQ0xAkfLkrbhN+NGNpluBxO9AnCO+KZ
q6TXkcoeQ608WhoJedwimX4fweopKpQeFN6BahyGJuhSsOEMdCvepsn9bgchmdXXh7bkv7jZHMe+
wYvROVgbYGXaKNBndaAqAleCS6eoKNftWNfQdMi0VXf3yxA/h5XLG58elgpISpRvJiUOJIgj4VD5
Oaq6khCYKD6ABRZlbsQ6x78rfl+FkXKVfB2eattZJY7RD4shclMZaEtdJvDNS8by+fHDAEhIf4uG
nR0oSHMOXCd8VOLn6NgLY9b5HD+WB6uAtQUeQYvRSHwh/Z6e0khK7mFmXLvRxmH9uJPLd3yo7vV6
/pVFcF9QubyJwWIOT2IcATMzDtT1mOfXPaTt75JHX11JdzGQzX8q0O6Y5IKT0YXDX5djjO84hVt9
4TnxfvrDcUrNch4+IdJR+fCuxNTl74YOZXrkjDD6WX3rTUN8rTYRBTR/5feAHATXZzNFeev9QQbq
AdI4e4IwTZNde0WyKJHxzR97Z0mjOnW4hYiiRP6evWijti8Vg8ds7i3Tk2gtZNQPD0qqXjSRwOfg
U/6R7BKTshxe/lyBOpZc+EON3zG8H19VomytSsg/VvQaB1UomR17Tr234iXSZfwULfljnQvd7qhh
prP22MyO95sJl27zh+7iByFHp4v1gh8Ofj8K9nyeTmk3p3LSzV+OxRysHrw6NeH9Y7A572WrIBpr
kkP223FqpiQcMOf/etYPB3lvNSXzdoqY65uuDcWdfW/KGS+gSNdwSFvjAtpwRU9ba5X/MGqnd4Wt
Q7OQZ4Z/L8BVFGt3yQb36dVbd3SRs9fX9g+D5LdpzszqT4jeBx1olYaTd1o1kp/UGdJlNW+srJTC
w4Pda8o0002cUMN/splKBKcFRGdHf75+vJW/Tu2L65/DMlGMPgkExcZuZpcs1lhhslVpmE10gvQG
h/yerEgE+YejY1dYw1oYBKI8CuVn36D9o4dzhnQXlzaQ4PEDaGLWgfSrIpjd2egfw/nmjac1XSrg
fUBwiKDqzzSR7x8Tg14ypsGZ0kU46RDQYdMSZJnQ0dloLQy4rQGw6Nm1f6YjVPWZkZLsopSD+Jou
mWFqX3crwfcjWOa2NtDJnVb56PRd+5e8v1Br/RzafkDK3q1O2laN+KexX3+A6QV6qTm5SDMTTNo5
nSh5xC3dTHDcDF6vSUNTnc/B8c0fxErSL3tWIl2jBaj1IqQv+b5nsycyj/iJe86LUuloFeaTk717
8dpNXMxYZ9RAeMooRzODLoRhI48MyNuTFN7BJ7wHAUGSHqWNg1+JiqauEatGEwToWOU5vP8F5ifq
SDDudFaSWjqYFk5VHjIxgYaA8S6Ifqa/z93tWeITqKY2t3ALCp3ZMv8/UudPSsgQhtALk0Fu1ERI
EF+Ytx1fDlqN89c7ZS6xxVhDnt/7pzE8vbJFvl+Vk0lzKzMCq6cHLMiCAd+Nwr1ky3ducfzlsfGz
B9EYZ4pISB6ZcFLiUwMKdRI5hViSSDs5wtmEbKWwCvX8ohRDBUtJzgbBgO78NcPQQWnGM3QfRc1W
miWyea8p07FZPptme0SgRPlNPKxBbzbpLRYbfa8Ns8ye3UQVXtwIzTlyhvyL/WpGltMJLkmrdog1
RgqYqRT92/Kl5kpyVFM5F8ZQhrHVBND+/fXmB/+SgcJx8iWuEtKGrMbICCjztrf8XqOk1P5NtWiN
e4vwfDouNDv3Y9UWxT1GtrsYqhFu2tJnmTl7oO4zsahN/0R7TUdcZKewTsLy97EbMWFw7nIKaU/4
msNo2cjQzWFbW6g/HTBMA5ZLjOOcCcskveYQoRJ5V7Z34AvO2+EI2XX0B/N4R/j+5YiM5oWlbeIN
Og+I5avbvdUP4Qx8WYv7g2+B0PCv1tEZUm1OhVPzfNj6MmpQLeLZnZenAlZ27SNiLDvy9NU8eOhH
5hEYNqVxNQeREEy2r8uziWGfaiY0t5VOcCKTcrhLBVffB0liRgs1bFKGOYQDQwDZkNzeX8QPijRj
wwEK8A/1rmOojH/cAa16aZZz1eLN7mZD6Op+kL+YkrAm0uqAtcQE/RPb97cKrOBuI3vs1kyIkRtj
3cjFB7k3VGQ6OFR2NlZfMJc2nxcU0CPpWI4LbIuneoiqBSI9ahjg51hk4bRLO08jAUnjyjjJjXgW
tDor6vSfvsoBycdpBvo+o2amRG0GWcHshpZxGkl26Kt0HgpQcpvzfUyocielHRQO2S7PpbUmyixL
HkBlboUQ2gvAgNVj1L8ARsyE5MOMLaWgMRrsglqxeeR7tM3vfYaZ8vZ/zCBW7jiVn5ha87ka+AFB
mtM8Axds4GuiMzIFzrhvfYmXLZnw+DUvoi4EXB8Dzbq2lLmUMGffPzV4+rF+0Vob092+y57l6RFg
OdQhrPRzBFlH9CkFxErV3Ji+qOSgxBTgewo7YF31jAx+o1CoXHiuWtPdOOq1zqRKIF57gxnwZd1a
DEWQdV/Mk4I8nlGmEmnKZd4YBW3ZIvR/YOXAwiXCFh2HEybL8+wk23DC3XYuWspcHo6JP5Zj/JeK
eEGmaatp/Dhl+62wHcdJWRsEdp1QkoezhD9ZpGPNyTDBq8aI3ONRa01aoY6GfXc6WG6Bef/oTRtH
/APabZdGt/oMv89L1dRMmf8buRNcVDr64Ko7SsZv9eCdOzKLSI/X5HL3CBPztNRokNZQzSJU93gE
ixBtlOUTBKOztB4hvLdctpKKMiY40Eal6tnRDSvKTLuVyX0nTR3gPjSFABYa6ktEdiwzpmt3/51z
SJYVGqNbARTMeBiXyORmU87f0p8kX0o+Abi8qw+VO2XHAtnjW1vo6FjnH0FMaZBBm1IPGomLU1y+
A16BTSE5+NR9z5i9rLZBYnDAzEy3w42U4isRg9Lg+7oLV1xtNkwxCokfTcwscAw6I3tfo0YIYj70
oTgpUTn/BFzPqT8jqz7wE/b87f2nkMmNTZxDcqYWut7P6SRyirajB+XQcb7qjuSnt52B8U4AU675
jU7NfEsUY164wI+80evu7upt6Z+c/5OfHkT1trvmYDpybp/q9h/Mqt9Ufl0rBN+eD9no0Nob6Oqe
BhgFLWmMnKgzPUu8lR9oQ3OXPd1YKo8KHifR1jwUwMw0ZYlnjoEvLNl8/7Mcx8yadOB9ZdiSulEX
X2PiNDG42rIhuNzVY8ThngQ/qVoHIDzOSGBEpXrWlq76pbZb/Sf6b6b12J/vKtHYZNKx30O4W4S2
b6+CQo7XM9g/pxJ+nPm7WW717RW7D+6Co8UCvMdgR6fSLS6wEhR/NTX98lTv3tiFzPSnhoSM+lYv
QDjq5t+ix6bdZRSXqgitZsbD3YrHwa49qtlN3dqiCfhAjSZxbauMAuS1TWX8s+kVL9JJKxW726JP
onLVFKP+R2keVdsBFpyTtMj+gj7QPMFsKMHX+yZZefWX0KJGxXffnsdVBqef9hvkR3QbPCtG0Rjk
0ZhpZ/gREwKEXO34PzXss2Yxk42SYVrZzOcIH3dhY0/QAt8Abr0wrS56/nTdCZulvtikeJVbJ6Ax
xp9Pz1SDhStnK3I7kmEVIhmCTENKuiyGqlkC8+YhfZk3IDxAGyMYIJCwMgML0joOLKIfsxQUrMcx
xmtt2gSYXSdi0UIoWhIuTgmWfi5WX7WU202b/lnG/RleslqbBI8eJJBLpcDQVp2mJZSDdjZO7B12
O0NaRkGM03PCVYkPe1wjzh+WEb/myA2ldWQlSJ+YxqERaM1LaRCqS/C2cRNUh9elNzllyLN9BwMd
g1llKFRY3rWXJSQXNGBW/hQwDd5+ZMjjxINASht4vPLHUrAoESiQemAZ1k8D8qtdi756I93GbKe3
170yhkY3IT0C+DXKyI9qK3KYBK4RHSJGLrdskyYBFZNWucqXT8gJ1eNgyYHqn3WLeIFYnO+HF9jI
Oc5V4fmRtOmkG2cAiDStYD1fXEvCJbwAO9AwMqhAAJvxd4i8YtPQYWSnzZLO8T3rswy6RWha+OTM
WDC2N8r5Lr+jaSVD5JOMCNHpixSDs0TZCT/81UtnZkSJoWGJzO+ojnl1YYOfHBPLBqSeCXQtwBi3
TNSXE67lKsMUgQ5VEeHPH1aCMTrBNP35DFlfglno2+IewekE9q90QX5dSCAFKgPnumExKkJk/6BQ
is0l6gGfeDg+BpQzYnQPRqXxgwy2O/GF3ichCO9bbpiTCR6JY1TWhBvdfTyXGvC6x4BJJauibmsP
YapnSK5tacUIArt9K7P87dtlVzTO/lX56cN7M2rK9knHKvncH7mdhQ8fGw/IlAMgTJpPYEeTDu6C
2PMoxx/aPIuvEZg0ILL7ZdcZtCMNHocn4zi9y30Iftw/Ir5oshy4ZQgWLujIvBZe9jRi8Y4eMLPg
4Wpd8oMWuuZrUlEpWafyuTu3s/uH/agPMLSnjh03togOg0Hh+7WNx93yXztUUN1BW0rGLTi9zfUM
/6TXVgf+QiNens75ubr985NIR+TBb4UbHmioiT9f/D3uq4ikKoknTnnKfRy5CpX2XUoUcLVQe29Z
V2CmmC913yvH/MZlb2hufD3gT4TcgRs+qmGlSV5ig2JoDMzGcv5gpOLzx4mXhqYO8df67j6gtcl1
Jno7X3veCSEBTqKjLeLjpw4FKZXmQHOEXQAx4hkNdL4yyvmcHfKQcyytjvksrCTHV0pfIB29z96g
hyjmU7bZVJ3NK+XPxad1U6LXIDluCc8HxLpwpzwK6pNOTepHOvfjfSGTTJOsP+jsx7ep7l0uY1rI
gpD3HNA1JQn3g+JMbTLaJbbi5Or37CR8T3PTCAGFODCAu8iRkNV9YO/KtxWbk2tGR+tTz5OkcHAC
7ZhAsdTCljGPBuGCntd+Wp/DMIsoftBumwOZ5c6OxnMkBYjIJVBgLr9CNaoOVk8nPjkmQX8W1lO8
vqwc/FI9qAAl8cViPyuf6z8TFw9REh5Wxce1CG2m5yzYbykLWCHxYTjc7pjGQgciWmgAQBlO1jta
0QLyepbelWEwOKlct6esdt4OFLo10eDBkP3I8iOLhcg0VwMRCb1wp4RIG8BMlwv7gNy29DyZcpM1
J1oEplA7DB4ZXhdBR3uiwFQfE8BL93POt/pul+Xgl+/jU2F/znskn6s0M9NaVXkli47L4KY5b3qJ
AjUv2keNjXwg2S2ObqueHD0xA5vGvu69HpiwjD9qpPDgwVs45Wg4Nnb6S4tj74jzwsDX/has/X+Y
SrHP4I6dUxqPJPHeKDCfDbbVI/NPtzvg2WrICCBJhoe1WD1S/gWiVNMuGeAcHFoPlPFRLA19bPyf
FmMPx64RIm4pofE9R38VHfVCDjcRwrhbpajaIDDOEmqETfCylYXI8lFofFIm5RrTvXER+hwcqbXj
C9AXeKJDiygL0O8YTy0CpG44TiGCKrpHNrqw9ZQVJtRfTZdkSvC48J28asL2ed/oMrrOLRJ/ggwO
o64q0CD2qkCdhp8G4YWt2ZpUDcwdGosGV/DAAnCi2OCf8yNdjUiM3Do+vUSGExw+SF1cfPW0W1YK
N43DOhKavbMYL19gvhpDB7FnOCajRfqZlYP14Di0X452HvEMWTf2/SbvjSFEeYGrpL7qXQJEXXaO
ko0cxiwXpVBXdKl/x4yRsUAJvCtTGJZQ0Y7l58r9y/6i0fi4VYhcU5HuO/5HPbyxfAUsUnqHzgLZ
xMCYmWercF91g4qIdijK+BHDZ47FbZedWjPIK2lGhDa4cHMGE5vxqT3WHatUVF73CU1MUBjFuZS1
frxgJna2g8vBUs7lS0shVO3PwUvtkAIBFS8bTW9fcipWDz/7lZm/3QiKoQf2EpYzFRPhjH1uyuiZ
dU7YrchAbJKImno4JnCcqIy2LK748kB6t1kH3PJc/dhVmKpFahbczvbNMwRqKd/oiY/dhbUzzAit
xLGfdeYdpgqu+BAPbQSmJWQMrt+37+q2JHAISaWI+dGxBHrSgUYJEGWWO3Mbcir3ghIaOb4qnmOK
7i32ad0r4b8Esdv71TWP3PGqoiZXVyMsTA08wjT08PhiaNCT2Cw/w4CzBtsVgSv24eJ6CP2c6Ggc
z7pvfRyi8nnn6DSEtNSCORp+es3zRq2YucqqXmwHLdhIswOX7wiw1dg5Wo51S5MCFr0mwMaymik/
5526wxBzdZ9ygFS2i18b1mTi7xedA+eovj3R0y0tTiF2ZZvzSusDh894RXQ+P3qLBTLFA5ICRsVK
Q3+XPjAcC0/KXljJ23k9acbi5ceLP5aemds3vEYQETnyUHldHRBV/4dmmxaqlauT2kO2Q/cEx0uy
fjJRg7hlI9nBgNYq5XrMbnufxftIUKk3JZ27kRkPKevPzY7uGomrXIHj15j5GzzXg3bQ7BIzhgEm
xV2RpJMBq6cnJXc6yU4izspzNCbHkyITFJtq25DRUbDES2aPz9L6HsliUChanlviYk+8Hoo06Pf2
ppiZCbA914D+kc1R4YtFOON553sMHebgwUKoTma5nfdpBtOHGHespwnG6MSw20S1eIFcJSCBscQe
95aamoZVNfMSgfFQtPg2Z+j9S0zWurQX2cpWUWbdQxGryANDUk3pEK8dBfUc9+infnW3ABDjMtKg
z4hDRq/y0021Gj73S/tIs1OQJoBeo6SOUq5iYzqR5ZkqAR6Hpaxm5xRQpIDUui99EmQoSEKxSrzt
HFNW0TdRXaekmj1IaCfa4tevihz0qFGgVFagFKUh+BP4vUbkb5mB6nOghx0lq7F3pBL7TxkiwOCc
+OFKBOxU3ijZpYIbAV5Yh3o5/j31BLJAwwIke6JfhoDCX4SXETG7Lsr/j/WRi39TiB9MbepLytu9
W6wJbPoHGpJy4Z8zmywECehNUIszSt4+o8AsoAai5KVhY+xJUBcGdp2AOZRuHFcoIcxYs5nAzOEZ
IwEf2DzndqiolqOPPQTJoRvVxK8GtJeJ5k6WIfbpk8CCmks8yZo+2f/AKPbZciCFR4b4yXGv0C7v
E9MfpkFlnARxmxdEggvkg4dtp0S5g6nG4+kMKZ5D4a9Or8MB6cDFXbfT1eif4WzE7r11B3wii0W4
SddjnHn1ySWpmykWpYulOSDhHDtxoyva0fBWz52/XFQbzoOkB7GcJFdFZvmhi2gQxNVfQs3Ro10h
Bhx+Z+w+4UbDJzzGgTmVqbfvaFSS9HVjZnxOckXrydcLAAbrCuA67IdzT9pJaG4W8HP+tlOkehD1
+BN59/DbyyN414kKp4H5jDVh3Agu+HU1NYx0mBpLiapakFSV9+Kk55UuXqoTo4yH6YA89wi/n3lT
NP9xkrAO3/1aooXScYCghcUTM6cRugWYUefXArx+itdDxhN8zf4NWXRsGdsOyiglSV1NmUWa31l6
x9lSmUIuXW0Sz1ZlYIvAxdoJDG7k6Hb9i9xTtOBNr3gdCWNvV9J0KKSJsVMFvHV5e2GEbUadp34G
TGpbJt8PuOO9jXbtGTWoeJ3LwSDlzgmZP7QdIL7FvRUrpPjxfzFnR2mjo2ZFV5UY7zBFiToS20HN
B/owOGAJsf4heSI1xln3cu6suEDRmcNO1OCRideg+VXwOLpS3CVhUHzHPyeP/S7XEKUJ17DOis1G
DsbwTjCzYj4p+XcfbHkSkcFzEcPJXyiBr04xYWnPUWMv3AdHYBiCtUHwJQb+/0kYwoyxq8s/yMht
3qOep3qc6GmcRvUI8/jngnyUBKvY9tFa582qF3FqdXZc/KC/Ej5pZ+WJk6GF7rzEKj4eq0ZhUQc0
O9TmzrvvX0LlUrLthSCtnWkQ1N9zZgjquqgZkNtDj6f5tO092IoCaCSf90RzV5KetBQCUWrtd6a4
UIgYJr+5d1m/lC1HHbYz7U+LqVoEDBiZLWHnTyjsMkIGnbOceH40ow2M3Sc5tmyQA6JzVpJ9Smzb
sUzB/OgwWaug1xIOyprTLJWCVMW2wqL4iVCirY14XKkcYFl2NmhuAbuRdUxDd9AvPDARQgtL2Snr
0dEL7A0co9p2lRTeS3eHruM0wiHgF5aTZT9uj4gHypLMqcgdOgEJpUlGCcb5nTMwct6AqEwAB7N2
03ZRCnin4e3Pbc0o3RSlSZWE20eCETfHPuJg7oMY2FsHQBDULuK8sp7Gp0ehufor5u63fNhTLnkb
eCvBBd6Hv7o+uvgvoCbV+RfFdf63CvkBvodkI9o+jNljzdcrC2DI7xV1cHUre77wLHZn8eOeXCo7
9DtyoVK1mMrq/KQgJp3x8mmS3Xz2BNHvIGXGZu8G8WKCt2/ULqE2KF9ltOf4fHhMzVqSJoCmWNit
zWh6kEeDHAkBhtIr1hY6P+HhszwFHDSayA7P+6x3GT/zqKoSyOIUXYrfKx54KxLznivC0ye95D8i
eAH541zlQolGFeKvZ1HYkBlPzfsbIdyeHkd+dxd9aRS1SuF92WYtP9iUzGDvpKE0ovNR3m3YhNr3
lyUnXyqiFvZi3isKbhfB62KIsTnidL3pWyTldW+nzEz/rqG1Jir5JVZ2+x55rdSE4CW9UnS9AFFb
JNaTkvlyaXtiET2/YkAmz3XiQS4b2/HKtMWDUgq9rxYSplLZIGWIxVHxB9uTuD89ex+oKEeQJYrv
YwrvBh2YEJtK3+A6wjlwh5TTF2FVlTxC1pBbxWTkk/dg38ov9fA7Svz/kxnqez0phvCyzlPkpPdB
ZkzvDbVQaQFvYYopTJv1bAfQ+BB5HsJuuapoScEcsuPHQ+rk3hvPoqS1Fl8M123hsL0hX/HRPG/l
YgGBSGIaGThJyv4igswJpq0Huc/XuzSdrgE/mVkkuIpdE1Exi4tgCoVeJcgsuLX/ksI93iUUtV+T
+VdzCBIXhHC7n6VdrucXhgQqM/xNieZJpXy6DBRJEh0tsNmRaIl7ElGy8SYetuoUVm5665LL+A+T
3x7/5WDixQoFfYPakN7ndMqiwnPLLe0MXFraBwTSSC/mN9e49ePIqj8B4H2qtx4ACas/kgigO3e/
QFLH5L6nx/7w9YhHLo0J6lf3byNnl2QML7pY3RvnXkO5rdXIfQM4pecVxDCmFqlDf3jLks4nyba1
w6qskl8ZB1v7X82bt76IL5pncObgSm97mXmgAQjs/O2ihhEunuoT5nN/YHOmT40fZbpCq+SOVEjj
49EFdZPI1aE/C0uAHxm22PE4T92Blt6p8BKcGvNq9du8pJKUGP6EaCGTc2hS4gcX54BSsS46QEwL
5DF5RLXG3rKW9k1/LnuIE8vGoPcTwkF40Bi90FduMbqi2iUR0EpporX2UkKQzp5vDhqOe629DHvw
KbVeCPHgKOZ2hN3GbvsN++SZwvOR8m/++68RqxwGzwD9IkO2MVM3gQQJY4HljjvaTO1DAVlJKm97
zFdErWDz9lHIieckNynu5Gr0s2PjsRnAStu7cv7EDCu6DPrpPV3LU3Np1YDhB1Mn3l/gWdXaZEw+
oDPlyhc9W5TgADDZUUMJvNv9nFPz0MfeHWRDnDYsY/pC3B004Bo9+qrGiAOrj8nBegdQUHnmeRRP
8Tux5rSk08frWvpcimky55T2Fl04Vt1Qz0eHxxmOXydgOOr1B6iBSjuvUC5CWaojHOALYXgPKsWR
9gx/jBrSHFqJrlGqGWIJWAteEQ7IMDih80Fk96A74blsQdnfgSTc1mMPHhNv05C7K+FS7nK9a8Fz
wGfidYxRhn+8Q/u4xyKIU/ihRBIBpOXLd9JN98DzZWkdGAM7fdLsHhqbIrnQWBGYob19ye02wFSO
ARCFKbDcxTz/96YAnPg0Ku2dFiGSHAgGuC5OxXxQ077jNZwUYRhgIgC5Q29dJsU8FDk9pmbQzBAE
TRJ993j2lC9LExENe/YC61qkN38oUwuymQJi1wylhwumBRrWl55YPj4vH7j1PLsNC/wfkMwvcuMz
cppehi3Zp3NAYo4RBiJ8dfnOasYLj5fgwcSCKcW7QMoyZHuVK3On0bIa186DyS6VI9ikscINx0h4
igI0dgikJX/biNNofq0DDeIY7wrboLl2R2xRIlcVZu24q4OZ6scy2G41GwZNedJWFYmCqiWBgqwk
GDV2OH5apUiLvCffBUw9uD9LDU7XNXMp7vMoJnqwplpraOIc7HwSkqDtCTtMukU28qa6wL7buvNs
mmSayKBSTudGx3/+oZscbaTxtE4tVkQIpK1TZzX4RQBSTrH2Jq4ygZkRY2YsJ+owXR7iUkRk43Nc
CTZCnf1Z32LcnNdTpgk0MsMwv1ak0RPRX5dxz8zBe17AQ5KJn/9eP1LY1hYoL1vhnF1Y6z9SZXEy
VeVSOfDlAIS/1ExMZzFv3RBHSeVlqLU2s344JRZP3PLHutNlMPZVJGSI0zZyXVREyuNSk0oLzEP8
QD20Ll14+8Jk93TC/ToM6Y0vS3rSf7Srouy1KLkBiSs6n/siwRBhFQQJ17WBAO1AO6iw5INAEEUw
0YZ7DsNuxxpKlniozagOcVWZSrU+E99nBgKoUH4fyMuc3FKLvZ+9zmn2iI4a651/yEAdJwIiK9S4
9f6bRXBn4+9MYI3z2ewq9qaq6VRtaf6e2UiR06asF/wuzGrn+QKxX4O0UAaUTWwJ3O6ZRNXnyViA
s13sH2EGmQ9fFk1JpsApfASnp8wWlxCW0w6B5WWA/B1M8B5iz4YwFd/MhSQYed65nmYex6qDXr3x
FKPVG+u0MUjslHaJYCka4fwLnW0yGI9+0IuYbuNWu0Mu62LtOt/KmMkuyu4Eqywk3vok8eo9EF1A
PYmePfiQhifC6+5ogTxVMr3yDV9vQTpd7rmpW2K5sYArd8c0992tR3fZoaYJyB24csLxclVE+uLe
/mAP6DhmeL0AyQM38KShJJzU9U/sEzWWkl+YfK+hzcknKCDzCL3xqWmBv6UfENCnqH0kxg6O+oiD
e6i350I0DZOq/Dbl4Xw6GRoa1dH2Igp7uCaCU8Pk/0Q72g4BbPGTNeFB5NnwaYY1KcfyqM5i+yit
vJDVm8XYdGDgfe+qyFjNb9/xDd/Cdurt1aydyYC5uvJ33Z4AziRYeTr+ql8tBSi3H3l2I7BKR9GS
a5ulFRoPhUrHnnVH8eUWCok8d/sY54LBtULXsMqujbarVTGoQHYdxsFV/jd+G3IhGZ+0/SDMl3pt
XkNzMtL5Fx97UVxWE9+kziS+Y/b3cm2Xunp9mm+I0XB81apUUHryOOlyUk01+SQQbbYylT0O51K9
2qoAWseUZX3CbPiPtLWdx+QwiT+9pY6aqUXFaJrCTYa+WoCr97TWB+CQm9z2LUAe/bRYMfRuRSp+
/qdk8+AQsjpRH6p4aHmp4+ODT6EaRy1g5xiXL5hx2ItTPcK+QtVdyO4eBEI2D4w2VUDcetSyJTw1
JFAL69FXUisdMS1kIflYithiwoHVS3mooxKKP2fhRu59RBCgpCxClCa3zAw+s/gB9Rrl4AwF8Am4
kiZP602qnL2Ut/6cxmF1kfZoQ5lxf+/O4Bc9w+Aen/tPfD9ZYzLpF0orUen2/WSLq+h8cYl3MmxT
cGxj+5kCkoojdt9ZwQTpAgXu040mIMTrXOmBOdrDx27LWsz7I1hGQOUpsQFnSRDDCJ+jYilf5IY2
MalvvYZUjSbTHixFcV/qEfoYx9FFW4qpYHVZ7/mgiBYODzAljzt3maEVN2vChJd7m1U+klGMAPSw
tGDBgxtfuvcR6oYmtzoHQifsg26bYsaa5sgPEX0ngVYuYmpgEOnaYx/8WdBHKdS7RvLf42yoEB2N
5GnGzPTFdHlQ7XCEPi0XPUwdSQPubsTs3KPdNWOvnlqikjPhbcqldkthnquIpDKfl3NXt1afaiuP
sbENdog8wxDqJFRUd5Smn7HzagjkKb2IuSsnoq0NISnFYYhDOAj+3JXcedIT4NnYkS4t5rLKo4di
0PROgLbItGcM4Z3NCYA/hrm8RUnCX1dci15ADY1+5r3qP/4evpOUE2PsUEqPPuYLLJP7lIIepa5v
2HOZstYNufC7APCOSDL7eT6Evu1uaYJGSgnTADzbneER7/w7mUzvFjJm1jYHotUgY8F0nKEN/09Y
vc2xqqngqgfW2tp+3u7nu30kjtPeWwjwwxMiQdcvf2VJbnzYHoOBMSnHU0p7qgmgbzudy4iNIpMY
eOSp4qakDRiCGht6XnEpYBcb9ICvOSkLW145QS13/mQJdsozI8KYZ7iHHWK8iJJfZFOVu0p06ESf
1uEpoNRc1eX7aDqOrFDIwTWtXE8L9v5dBJscIM+ZFA3QR3Rdsp+ESd+soEW3+hzuQFoYI/3D+MEb
moALIicnU3No5Sqx4LOcuHb3nXFaPCV4teLRfXfCelMeeIR/NxHBKHAp6d0U88AsLBxSVlFzFgIJ
S2f4UzNTb5xtPHg2hhvO4ttwuAJxz/y7gtNTtlwGXMeyetIPmIRhtzQHtQDlEb94hNzvaYNRQCU2
82c0gKszyNw6bWp6QBGkImlwTtGs6HgBIoigT3VQo4mB1Myta9zIGdtp3EXSe9ouzoLaOfL4AP27
ZQOOiZ9iyk40jzwxHuCgZJ1kyeRqHffz+GsJsz16ityF2jMFsPkVEFan8pzXuJrBpDcVwBtj31+C
hmuqk7d6+CLCh1R4W/b/Uvb8YL9mzoE1BBY/xExbVBIqWnko1oqg7FH6wft/gYhlflJzH/8MESw4
d7zn2zNUkOlVLOQS0MXj3Z3LqRpUNrEuCpPwDiRi/9oRyi/CEwdQvA/EnQM72rvD+bZOFCpFnkdQ
9ab/aotmWvAlw2hwvKMAVXMyvOu4AdU7/752Y4nplm60x9W+DwhqNuBbo8zTqVSKNySVh5DMTzXH
XZQJ9GZthH4pO7RewHMCAyPmB1aoQxt/kkWrd1VWZtWotqH9VpKI63Pcn7xIB1NZZcuHtuDfWaFM
PPPgYl/YIQaLVk7uejuRVf5VCL7873KPre1wXUjv9j8qvq6uMf5WYxF2bbafQJ7zkxXdtsMk/NY2
RlW9wfE4enoGZNgxiUky5ZCbr9a+1ecAGwb8vuBvDkvuOsp5g5ivoaWHOaRPdGNR1P2IG1CDexnn
l7Lbv1i29am8jnv6hCnLUaZlGINfTb9081NVM4+wDpOE3We0XCT2xcq5EkLk0kYFIz/YQ9ecX/X4
KySPKRzMU9/m4IH5XPlRhcsxxOyYRpaCTTtPRiW21OJwMSr7ly6HkgMQ8u+PoJm2STdWDiNRq6Lf
7rmQISwI4snCetYdbCD+2MLqtTWpEnsoYIY05cHgyUoP724PvG9owMgTms2vt9SKTh0PzSN2NK8y
evVsqMCeK/VahSRNQu952lNvmeKZFI3w+KLcz5SbRqQ2soo8hLCNOQ6kgVpTd6plXXVWVlrRNE9K
p9m1mXwvRbbqVijc7E23qrPeA4r9yqlkfoaVfG4JnSXB8dAchKj0eqQTmTyK4nWOequQzUHaDP0H
cgM2acjgzGTvDUrIP4C7XIkb8AGl49RghGskKoY9cv8dSjri2fplJ8jd1bALOhKpzEhJFwoAv6Fr
xtZ8pp+H4Z27WU5ONYjxiTBg8hjX8rhOHfWcRt6C4SqcN54oKmb+ZPwj/HqGLDl7xx5WVkcB5BzH
+lyeFm2hqzfggs9gcWX26ZHIwPc1eGLZc4OCkb9uKjs4njCR2vjiLprjriU20FLATrFSwBL6POtc
brbTWLwGXzIDqxcTi8Ki7haCLFX7Lm5h/2K5mLzxKuoVxDpL9M2v/v42ytxLIZ+vzhNmUNXm8Qli
ag6AkV3amxjoeE8+oGyFul1NaCczPBvtE+jf65ofGASbfuC+VlYD3VtVpX8asQTL7U1IVbccs0Uc
8wboGYmu/lQ7naSC0LAVK1W9CtSruvrYKgNzZC0R/L23dJCzqOeIS/92Uydy8uw/qwnSW5oX9zbZ
ljQ7QYgKlcQcsnx24MAg6etVUU3qUDUE7ez1UFCQ2DW8rPTYmkRjHTQKpwDY8ZyljRsB9QoydSZu
E2HNMStxTZcQJiKy3CwLKdTd8dbNLCZJcjMwVM0QhwsA5ITJefSx2iF87QF7Hoz+IE+2Yj9YNrjk
HC63KF3Rg2IRQ6QSIuruMrnPfE0YserjJ5POil5BU+YBnWNg9qtSy065C5J6ZGKQJRCLft9Q3Jd9
dV/xq4jqpzxkA8c/Nt+yaUNU0xQAi9ZxyAf1U7EgN0s2ilJw8yakjctvMSEdGJNT7a0fEgmKLLha
OIJqvBkLLobRyri4aJ6ZVpYQEWFXDdjK/hjTUc2rtouHINIylNLne1lhTNLZOaYzV8HNhhwK8W6j
aAm4L9QTyoVqCQ42irBfXADTb1GHGUjHhLlX5fwaehol6EcqiUSxVnC3E5cSKrrvfU3XM6ZcYeQ3
+xiY+pazSpqU/3rki7I7G4IxFIUbznQr3LYT4IsOH8dKpNpUbq4LRgmVGwvRP10PkQoGkjGRkLuV
5Im+LTxY0SETIee67puwJ0RmzPlwtNUQHE2WpYtnwTiuJurhvDPY54gsa+3SWdKaei0w6vUC/lw7
/cHx1gPZL7qu5n6O/r5gaTZoQfs6cLipWFxcCD4FEZawfbUaXFbU1rYZ2apKeSYHi+Zd8pXTbB1A
9/dESm9z6IV85IMqUo8Zvgee5XfoLU5X2SvTKmXgiWouPK0rxv8+Okh+ECs6QYKv9d5ooq1vOP23
IO5EtFi5oszUvyXZ/JSppItmAOovJPgCkfG/DU/V6uRmO3T+d9nObg17k/g+CayH0eHrrk8DxbgD
2o61e/rzN4QaySDYeOpCx/fmM6vf5EdMqKrwWpPb59BfI9Au5ndoFf+IOP9v9dLr5wz88mbQuo11
Zqy1UzsLiOof+1dYz+HFwr5F17MrXqQStZf061caIsbjHifwqhIQFNTN4EaLN0vqwW7bw6dIZ6dg
ItUzDzqCYaCiJqCgHBTUpVdhZCK00cPN1U3HIVGgdi2nofEKT6nRsJ/TA8HigzKIEPBixaFVAn3O
1CXVtyvmFOl+Rk8rvFblOcG3WSldmZOnnvGN80lgczHHyr3gfXDPirQomkDj1WCFX4A5A20Zv+Iw
Hptyud0c0iK7D6XzujzL1XwYQ2RqcxVEko29rbA/1ezVOWBS7KoVVQbMAyriknI0MRbHCcpaqiAv
GLf0/Xki/HKh1AcyIYTNt3y/TkBypvIrRkbsP2F38f0DzFB8HF+tPCmxAuOQAESdouffTuotMQn0
N3Y00TuIhWg0Gvkggaz30Z7d3s35F4ejooC29ZcUd52W1tty1GXYt+2Wh712ELG9fPPWhbf9XiiM
7fNfm+XjGBkdziNx/x+FWWJ9nHINsANkN4NF2qNsNEyLogWLRDekZNfXBZo5IBdyZvXy9E7jZckB
BNjePLm0BGOF2R9MmBKGJL9qCgcq2wnCkqbhv8QOIs0alxJJk0AqBlyYp3KFbaJYIUh5cr1k4qOJ
YUjfEwv3gOfgFqepCJVzKf80j/eCjyQuurqM6+K5e7CFBLPRvEeIfV2s2HGUAKia9pIL4BhF8aGX
AZiu4N1paKnY/IpQbiFXEFJON7NmwNj83NueJzOcz88v6zwwYQsKqQ3BMNtXc7AWQEn3rgHFgoq0
r0Sn7CnL95GWnwcIBTdAu0XWXkAaJtgedS9qUKB3yOhFknPObVpQLFKwAIJPNJvR0V66LSJd87dH
dpiOVrEZGCg39AwF3XGyYvptvoWFbeAjXj8s6i5yFWayLmrefYUvmGsZwWxnv2jnfgs2dbg1r6Uz
M4fTThkQU4dqbdk88W/zEh++T/RshGMhxPgsWb2Q3tgggRLmulrfzEBVIJry6cx/sY4CmX3FxBr3
PNeQazv+jdAIcas3YWJ/0SapWPThSHgNVK4sI0yTrBe1q5LFLjA0BC+Cmbt+j7uSki6gNvNryhF4
H7YyII5xHrv78bDMSzc+8KY49LSwHs6N/OWtYvLQxnNaGFRCnlYD3klC+HHImLBreryDZoKI3owl
FOH3/hcZHuE7rXLoWIdD0d15KMZ0IE21A3YtNjPO0GfwiElv12Xhq1/s2xOcgrFeBLVSwNc5Snos
w+sild2s+OHTrrkEnIvvzIdKas5ieYnigNGsBbINsFLGuc4dK/trjRrvsWKN7WIuia18lmuaPER0
SSufAOU+l2XqU1/iMxgBsl/u/GKazBoDbWTX3E1Gf2wGnfbZ56RWZWopo/fzjS/j8YS2Pmbz7vlF
tV7nfW++4FFbkj3pfZ+Ky5jBCeF4jw1dhn/SBzeOcEjafrfC3SBGRrW24BK71WjX/qpgKsyGQ/6O
EG1AgeWqVQxXKXoMpojdW+svxirdbvfkgm7D4CQQiMbx150L0f9DSZY2gI/AKu1Rfy+g2nRY+xiV
pLatEqI35Z3HDGMPKh8bPgyLyXKnWLjKlfUFSf6NXLM2yWjo6eVFAIBwogjY1A9mSnTL63VOFXlX
1yLFXiERfJmRV5ZztPGLwb3FzoHbmIq3pwTXG3M8Xwe6ZbBCc4lbFMgjaLk2jJRUvfYxxBYJliIt
Q0/m4+mrjcwD4m4jyu6KU2FKC5+1S2CcUQjFpz5fFb7HKMzOj2biVCrqnPo4kv84XBKSbWvZ/0v4
YHF21knWsX9QZ/IvFMsmT3slLXNc2vA8h58zcSgLOSzo2mfRd+omPA58GhU9DTYOUdClZNxJdfyq
c1cEsP237ZGUt4l2QHBfDRMh8JK4uVfFj2fuTXCDrlSGX1aFKU3PHphBo5HbBgd0jcyrqEm8ewtG
F8LEIQq9YjM7ci3/lKoce3cZNpA9HiPAZYzSlULr3DycMhjbNs0Sa1E7/Xwcqf4VYJXG0/ts8r4R
+dz0S5YQSyKyorVPDXckfuxJYgVNUhHsQl4+QJqksT8fqiEFUkRu4I0UE7PA5Eawr866zNVcK7wA
SoI5J15LvyyjMAf00gsODDTSZ0jBByTFt1HVE+YdKI86dxBl75K6TOvnF5fQzEI3ExVuNAOMVu7U
ShIZWOIoJll3+uq1A9NC4HRlEaoGYlw/Ahl0lkam8TaJ4pNhMuGYQWqBCfRlL8XKdwuJi615cIM3
h3Spu4LIsLYPG9y/W9E8Zg+ctKsjpNns3RQI/cF6X8qA6vCIM7LldtzUs/5dX5EkqKz4F5lrvUqa
NDaotQSSt8E4uxVrpOS+WRXHPFIJPpw6wIOupLjQNZHI8y64FowNaSbR2sg4Lu3CZPnbFghP4M0h
l6yUTh/JxzNE7yi6zaGZxS7QxPlA11wYwC7Bu6CR/CQ/9aLL/qyPKOr2JoLlCJ5T79v7o1v+GMBl
xpl5N135ivCrB2g+bFjVduEecDjevJN85LreQRmHIMGWepkkvLb3+8KKaRfSLgfrstrYx9lYUU4D
TISXfz23ObK9HXfezzrjmiZLsdebsUH3dkgunN+9ChVO+5nn3Vi7GCQQHEqt7bvcKxyohPICk9XT
I0vDwlISvCci/taLuzN9H2BY3JbrIygABmw/HpPEYOErUnFP6kD+PpoBC0mg6CVKrE9uAgGHi41E
loGDESSgMmkxr87fyetStSgMJgmsTVJpdWYhDwEosat2wxYxvysT/jQAq5xL0moklxJDm1Lr+KII
UYsDJvPP0+3OFD5mxjdToTzQFxvWkuMAL9/CVgQb9uWdOsXcugLmOFp0zmjHPPWKacFx5zjQBqXc
Po3Mn2bEGXfws+dV5SfNILgOX2X+SqoYFTdAaY5Gz9QjTPmQsoUENbr9DFOIT3n6oa1IRiNCVNxw
rlTmu++eYN50qWK5Vy+6eugOu2FZl+o6f+9yB3k4N+6VxRWm196enZ7QYph8xsWAQtsmUDikJtAo
K2QBM8iKWnaneyj0HPv/V4xNa8dOENP+WjIO7LzdUWn5POce5CgluKT+AxtK6bUqXbxBhA2hXZ6t
alg/asLkKDHvqih18I0NntiGaSFl0ICV3odnUTO3qEv3H//mBKlP/jU+7fGi6IFy4Bfhy5K233ve
O3fOVMXlpOH2uF6ce/p76MNYmNjiYGufGMc1bM0bF25jZUYazpns6pTr2TeJHwzbGO6dquK7QTBR
3SXwR3YkE98kV5JNwgx4JAkGfe7cRQ+WfVGP58fbJFIAdJixIISrCbVsf0BcQo3V1Tb/UUHYjl9r
8O15dg884X5MdTKITyLzzMdfo+XPWpKETf9Pd85wD9m7hfOw6jT5ipuj5iO711keCSQwf9Sp5G7O
o2VeyISrz80GWV5wi5oAy+c+hpDiz4VN2N09p4+0npOHlvKapk5U+wPOs18RA9vFTVFRFY898Lfp
/Iurb7HW2atP6c4MhcHrwhQ8kBNmodctwtMZt4e6RwDyEwH1BH9UM+EsvYmxe6Nc8albB0S0ibUe
DVrEbJQOSK22maTV4EbMTuyc39KLxRixnPljdRZqrv7KZn79jHki7sI5GtMP/dcopNEF5wuowO4d
iXeyO3zjMc/OtTqgf5y+rklf+dszs3eNw0TtYyejDQCpFT+ygi2A4D+DlDFsOuQavR3C78+iBwaF
Ws2UVab+eJanCmOD7Oqlb3G5K1tW/ZtXXO8VaXFLr5bfcdSho6GnNvabbll1ANsc2h5frwjitqLw
0eTP0655W3ZeJuKKesBilBXWsbAtLzhGVMnLQGi9cqUFnQwSzh6EUbbSFLnzO9ojFxA354ALuu1j
6Bqr1a5TnDMKK/Ifu/LBX5PEec3pzH+tfzexyQDEVTZSfB5hsjrpe1Mg4/SspTQNGNyLtA93ktO5
bMVQh/eLfU95tDizDabHzFnuUotFrX/lI++DWrG3tXfj5dnwycda+u7gL3QXln1Dx6nHxJt4EV2s
7Mgt9CQIMSEOlEdNYroO18klhZUEzXFtca32GuXU3cMdshoxr8ZRORHU2881Vx9honoT7nA5Nvbw
4XYC1NjAMU7JPfwln8Qa5uHhkGIOo914haTASJmDhg1ijBElkfuxQjiMw6DrKWKSFFS8iXVxNv30
cROzNmi6rdEecWm+9bkeSJBUsUhWWXN7JBnit5hEjQMPMMByR/0RyMWdg99aBnWXfGyGqWcoYMDF
n9qEhn7Vt1hun+a1r72GZdbQK4pyASaeDbCsovrb5SdfnbwmVeHLTj56mcATKIKmUkbrIik5Zx9a
N1O+xq4XSWwTrybWS0Z96ima/sQYs2plyddusYU39aAhA9OsjO0jjOpZ2eJrPbv3V6qGjX7AKXwe
M7LDFu5BiJJnFOABOXc+BDcq+uBoLketyHOF1xQEnKH6s2yU3KsBFxtNvc2ZOiIYD3cM5yzJZVA+
i2Nybxb9g4desO0nl8dIkJNapiulTxmZuQKHhpa8x4DFjqJc4q3jXikAaRVXuMov8JnWfUWIX8xS
+MzRTXNGiqOLK2yRfh7TnSURjaAaT/6gSjdweU1rKyAvh88Xg1upBJKt0EQZEw6wSNFj9jW12mGZ
6+bXk2LGXJqiOplsZK7FCl+Pcd0LGmE+x79J1UE5tyWKuJku68gYAvE4UitQZ65YIJ773/d2G495
/PTaNp9uY1lGnfL4r6hJrYnJ3nZznHR/X2RO4rwnXHOldy+9oOxbe9x3PsKz5EkK24lCaG946JEK
U1IIBskp4olU86QEo4Y3U7JRRhytVXKNL6LyS7Xtn3Y1EMwN6OR7PuFeOipayPvOOciB9/5MIdj2
IujsmAl5B64qxYKRaeDt5i5uhtKUQ8CHfDzrv/RZyqx8fXJXcIx/VBLqQkpd4aTQ9KH6hWntPQ3b
inOaPlyEyOF+mbZO7G7BKkexHaS8rDB0kMsr2esGRXYs+3JwJ04RfcXaS+/H82v42+W7nGWr5FDJ
hduswez+cID9UoM2sC8Ln0MVZg8h585RXRCtUfhX+C74rD0tVlvCRaJ5ozvwkkuesBji3YPGG7yA
2zCtX0OlfH6VyrJcurVxCeUGVujCOFQAj4/0NDO7h9ojhyvGdmCWL5/WxQ7lgwqw+OWSq0/Nc+en
a7DqhRlz60Qr1vdnOD83+N+xl8+YNWCWhsHhaxvgfydWw7A/oc3/vuqS89ysAhocio4mlDmV9mbo
xU9Jdoymiak5OJv1Wu1mkOqlRNg8QADcdnDbYT7Pe2Hv6OXQUHxgKlozKtJYO3hQilfUsx5QHWwT
Zb7GZeJzHPtyMV4lJajWvzK5pTv3KBgPIMROuqdG4GuuIxPeNZC9V68i7nFhaaLlZkdQNjjBZI6C
cmLptFf7fqTr4B5Jh5QT8PmlSlhZGox4sSbws2YyTloF21qbw+W3zmiB+0bKjrvzVg8SpMseFYjx
VejNx+dZNCvGbyFTPWFcJpAvdRfI2Ft17NhhXqmnBR/7HpA2YIuIzonnAC66x0jmpknEkaKLlWN9
hNNJELEV6ygyivSeWApii4SurUzfGOB8/c6tjC/FCWqcPBQcfGKRcVJaWdj15FBbEtu3WCm4Kky0
jGii/B25bSdzTXEUtVHAftSBHP9ORpzm8xSYJBXIWPJkHemBOif07Z/rbEMko1cRrq2UXMAk5MgB
wHgPsdD+H4hIKoHWtw7PAnHxgxZZy9HzPiKCuOCvMbkfElKks/kxMjp7TPkJy6pU+qETWyYJlZiA
OknpzjCJ2ncXdJGqypfsM+lioErfWTWT3MW7UPrakFAjFcwkd6eU4t3RJVIr1YPbOdh9fTCbS2Vk
EvdAY3vrQ/z5i6Ard3Ea0PdCybaQGKwDJds0laEgFUjFU2Q8WeiEWffuUZRzV0F4nOd47ht7mPnf
E7DqxEsiNuR2qPrf5HhJX20Xtu2Lmu9KKeu0XcT33kwDlqnBddaaKoaqGlzs8qOEDGFSsvmBQ1gN
BIWY6nt5jh0L3Xr22HJJDYF9getWm81P4mI4lN1cSD3wWTE4itPUd6l5bqwdsSWDn/0e6IfSqyUL
y6C3qiyMKV/eS7gwscGYOfbYXyzVfPCSJ9weqTiRFor3oXw7oWQ089Gvqit/4tqWYp4SZck1lSdN
qa/wri4Gh0X7xdZGObiDKuKe9phppLjZTXFXCsBD4QGDc+i0GC99mKM/Xoku1JGo9512lJLnDOCb
u60t3KjyI2kO8fsATyNjM7fjzM8SF9nEPfq9kesctuIboWNueW0HSvljaOSri+mo8YDmDNhjLDGl
cXKWqIt6oqU1cq7HTkIVDdKDD9wQnGm5Kgdutl0okQiiemtATZWM8jQ4MXFQPwqsFVvF+PuIw2S1
4aDHKwWNDOg2ZPhyk86EqAsE/jBxuBXY3B0UA10IfWTlcRVm0DFsTkZ420wvLQWbSS9nhPYO/Efc
SO5mJegNcyqclzIfHNhf8uB2fXWB6pxRlH0mlSia5WjDjG3HHyt3Yi8HNgM8mIumlycLYYTnQcS4
vnazDco0E127EzQ33s4QQR5W4e740z5UmzSON1Jd5cDsbyKEp0uuUVlHG+mPGXOV3Cg5S88TD+Wt
z/pl5Eifi4Vq+K6MQ3feDQPeLwnPPkZzMtIUddW5ToBs/EJUv5e3QkxJ3NoAxZPHoHp6J4hGllPp
9xdOhERW7qmFjGCOgysdAvkYDAsdDXf73OGLAOG6JLbpXlyITu86UtKWOvIJZ+pl27nLc/Km51OU
PSWXuCkJi1QesTt3mnnvBvKHl8LpkcTWMHwyGvlgwTmAeXcZ2V6QZ+fe09RHwEBlVdd5RIg3I05a
3NXw+p+zrKuT3QlJfX29TmpJcDveK1kwC9Ut22IbHewn+dhyvAlQWOGh/Xddwax9PQZ7VG5b6qK2
MXBCfyQCjB2JSlWnAI7GIgNXmnCauXQl/SOV1jFhrT5X9EMJlJaFjA7q5ypp4ZBUIADm2WAhsbtP
JhlBfAnlqQttJEFsHEJJkKqWSltmB/NoPBCnf0jf90V7/jkGaiOXA1tFB0Euyy1np1CZ6rc8xuvN
IEGVmTWr9Z4xa8P7/q4BWMFaXkYhN2GUx//Y3o/0OaVqHP7Sdag9s4Q1eBMpiHiLWtoS8TEN9Aqt
ZmLV0r/OVvwd4E8dHKfm3WnkqlPQPjR/r9A+OCPmFYJInpDqcQMXeBWSuKS1QgcpGVs4KFOJqIqt
Koa8uzkbjB1sUiGTBufkivbz/N75u6IfMVbtRUpgK+AZ6Q7etPDmj04X7yNwiIuApAp6vqGt1iVy
mizB04nGTJy8a5yi9sG4/2ENj6rGv6w8KyLB6UhR08b+EXruG44ts97WcSm1Mu1txHR9Nwleh6er
6aFm9CgSGITZjFaZswvKOqM4FC/fplGyTdBf6tB7LO3739YXijrn/IQ1QUHRiyBTmgE19x9spaGn
SfH2Ki1FuVg3m1v0tAku+D/9iaBZgfRPcFJsc1fk4nJu6SWYjzO21gUG68lWdhuIxJwLCjAI7fXq
cmuCKNKajnA35AqsFkof2NScZHldxxZH8WUCgwIDs2gGebmz8zBwl4RJ0eHRXkinuhbMJ/hblHgc
5pdNqUO8mephEo5iO/Nxi7Mv53mX+0YiKmEMSa9Vvaz+nEDChh8trP59/bdqIDd2NhSh5WsIpTeF
4nL75wJyJhyekjEA0nOVAvGpN4zFL2h2DWJr+CUvwfq+h0PSAiDGAW3+1veu1kFO7QXeeFlvJKIM
eaS6izQnId3Wag+h620DBpmgrmuhBSL7tBc2bR8k4v0YrGJJmZt/TXOsXZxaJL1Ph1BCS3lFq7O7
Eof9Pj08mg/ni1A84g3kOXmmwbtC6AuFNJ5GJx99E7KHEE24MLU0a5ECZiTyO6g7Y1iZ2Gr1PvVm
lmSR4JQ4GT+fjmgKLJK5YMMPrC9kvpjeZCjD3+5bmBP9CB2M4dltcA1cbxCeb9zoE42reQfVmXYB
T8KNmqYYaXEPvB9RKL2ollWnlWFO9Wo86AwPHf/NhYdSucfr7lGLmZUnsMJeot7py/4Ppe6+VAqr
+wcuidZqZroRDtvmuqYnXir37/iZUT7LRAmtfnQ3vSJrQ+T01iEWQ+UgQpLToIjAhnOHHKnsoDxm
MKO2hPchnu88FtynidcH1lURvdh9Ltri6j4W9j+SnFv8etd9KoFQHBrjfGP3r4l631JU9ObDsk4l
fJjROeK7QLLScnQ/qJGzlM+6+ipqE+Iuk8bHszsiqSilPLP8rxrKweYb5TBhs5gHe/5p7UzL5+nB
C4BVsEaGfY8inZ5qBvT2S1+AN+tRH8NcfIuSFcCRtKqAIYth+LibDdvGz7tqbN5dpG4vRTGfnc7U
DFoJ5TZo60qkT//gAGO8W2wMGY4Hq73X9NtmWOcUa2yUt5EGdv+Ir/cJwttIWTdlxw05oPbbQdlO
3lAjw1n3j4m7ehTGQGwngUAPz3F7UWbgV7MNSjgU5/oV1zBpLzhq19wJfA/SCFSZ/BhCm3RI3JYM
nETr4T5NlMPbzhcR5ZLrDYF24D6zPlvDpkWI8dTE98L/FwUuQfhYta9X1P5nHiMvBWZIxcjaFnT4
dFHfoVDqatL//Dl9Eg6hpkqVsbtr8+mdi3QPxZjApfUXqq28kmconCAA9Yq3AVoyOae/0i9qMA/g
FNutkGDplQitUCm+4CGV7xLjDIuoLZyKRYTqPXfTIsSvxqTFfX75m6d5/TwewIz3XGV7ATgQ6WqT
50EBqZSZ1RnzCbRAx7kf+DdC7lnmn4oOwv+RpqGc2E/aLuF7p+KD+xDJPZCXAfGqbna27FnMt26+
N2Xn1HHrLbBOyuqWFLex8mCMM7uk6AC/Q/RgHXaI0B05iWYtuFi+GlqVAPNZk/CGzSscSULmdO47
c0qDRDp6EptHqAEhlL8Y3BrT0UR5O+51kMxEHaZNPCabcccD3TrjDDJodsEfkrReaIwFYqc3Hfza
bFbJk3eLuWu1C/OgNwmG7562+iFZT2InK97bd0JKgD1giGY3YgE3PS2riktRDD0Od5xlubbYykyX
a7/wiVDYfNs9rYcW2gTihIroeygXaZfUV/dVi6pHs+jj7r+Cvi2q7xZM0F/IlNbsaffdb8RpLDmP
xHpafubmWqTSHSn6Txpw+8UDOu53lYNHh/yhiy5jh/CDGhhWYSnr9zxg2cAOAGajnbvDJRE8QGcW
GOI1D56ZVjZOmJNVQLhqDUGq82Ph6XzNpnBJGs44aoMuAJlpiE3e4lj2en7LDcd6wOy9Lco4pOZ2
8gNmbeC+s0PTeUyX9inXFn4ynoM2Cd2uRJTMEVOHPY6idMKI4DX3O+Bd3nBvDXoJKnzNkBrr2tvW
PpHHev0SGoJ/ORG91lED4lbwS/CGs07OuwvPdpwKY7LaerXooV2CYk6rUDuadjZNcdRMIbnFHAi8
7MJU7OBKyio9S/FeQzbzfMHKSPAJpiEcP0+TzJ3E+HMcZ5v5AFN3zricroCD0OVbXiF/171rBKuY
fGzaph6KWJDTibST36gOkNMIrkGvsvMYJKcYgUg9jIoW6WAyzq0V87dnIFXWI5ocobIn5oh+/1Ug
+kXqP9NnSRydXhvVzSE+G31KKbvt2C8iwlPNS4LCEH+bs3GKs8TkefVnfYDxoS5NYmUDhGPO2eTY
mYV8XIGqvRgc2gCKHSf8zSSDz6IF00C9J9h7rbg01f6satIqzMfMbaioLkua5o/hjhw1hltMZezT
INA9xkhe2VL4roBXi1s6/DvIu0NhcNy2Ka7Ay9F6SF3zWXu+xwu91RHj5etUdi1z9KAEQiZBMpS8
xStlvRb9rqcKpwfRL/wnyEKg0vPt7qBmbXGbis4hnrR83KdnaPSyJhzH07WMhDCoqKmVYKXaTLO4
mEBzBT7f6JywvrKqBbcbFARsCJGNWTxsDb2IW+2Mq8oZ+NEAK3uf17cUGlQChIKGS2Hbq7Vgitur
T2fEZlVdrx89LBQ9XGyxQZA0D+FibXyBvJQQKS7n0Xv+c3uF6muteYgHn/VlFx9kzzFS8nJh0/01
1zN7CAx4LLwy1rS029mT437I9XDAXmoYIXCWD467Yf5XwOJ0Gz5iYYqSC1/C0+kWo1WCppZu41RC
AIKYnuIvLxtoUX06U9ex2zhu4QvBkrSvlrTlqN4JFqf6644T8JAB4KiuiqR5kjYhYkeGvLN081A+
Byg4J7Y/4uisiGO5tz8/hk+Lh5P7xPE9LAWYM+PiVb6cEoXKYwqGjuxk5Rok9WJQP5I5MbKYuH5A
toh79/qNYdaKloorOqlSE+5HTP/0fZL8Toodc5jHCkPkNB7DN/aZjTkKVi2ZUVCz5V7bcwqjmzz4
lecBdkfMe13yyyU+ZfNoW99cu3Sqd06MDK5eE0myc+Ql3AuMRilWAwnmnh93BRaoMGusXMo/Ix+3
XAdvhM0KsxEvkuWcW6fXXIUL+3whJ4BWDNGeB6Y/W4Bp08jURyEKpXLBPDuF4JX9emIp5Aadb864
gjtPf5PQm9+53GmNGJMj2OXX7goBT+Mwuf1znuAOCcIoqMEVZ+ZUVXlb72vA7HfCNeXxyK74MM68
RdMRbJsoY1flD2iqVfe2Xj0O/3fyBUCKd0w2M7ijsBWqsyWDIbv53S32jx7H1evUmAWZSBbsAmg3
uSKS6ngW9kIwRSh3+OQflP10MEG6AHBOAKIIZbBkjshi0LMXhcv7utPgN4F4cv58K7jTl3Gem0M/
msNcJjO4XqT25H9KLb7DN3GLf7W1jk/UN+9MmFvTwnJk3DKHyThTsJHQ9Gz2t2Al0GUFduWoFJjM
rqiWoC0w3BvnMdE3PLr9yVSyvBelxluKt6UMmnZp+daKsLQHV1iP2NQe3xLlpOYk/JmeTl5NMU2p
4EFvqK/AkKlpEhA46i0umXl4zXvHnPFhI1qt+jCT/Tl6XmJweyDmUCJt/IathsKwq0Cs6aNo1YyJ
Yq4m+hMi3fFqkRKj+GlLhyjcwiRgOSnNYJPkbLIaX4HN050CxdIpoDP4o7WAlzE4ZrcPaae8JwPi
fhlRTL17biOSjM9R/6Ffuw7sgM9Pvj2aXXNZBtjdJJLiWlKXpJAQbxsrq51K5mtATEA2yMywGA99
NijyD7xj7KuhSYBDObG9hShzhIOvIXfgKOLMeJtCK4vgrhJjR96Yb0VCSWhqRfOt959UljPJ96eP
xRVPWwYkhoOu8nsGfd2hnhhjZVsz0x3VUC7hNDW0MqDXZXJpia5LD6GV9AjOIDHEmvodf4Uig64h
VcaqebLq0SXF6TBYTSgU0zb1t85VIytBophIj1LuXg5KtlMo8K092C6W1UfjXwxlC1P7N/OEKTpc
ngs3pdFduVu4mwWNetYpRsgiykVb8JSFtKVCtDVGj9QuDNptEcpmsAUCb+QTapTitDXrzLYJttIg
7WFQMGzyxZDuo4D4gkoCy+U7h58g/iNm1KDN4Tl2fodibCsekCFfjaRpBMXetDxuHobv4k0DdOWR
OVTeLYFlZyfD9dmZiPek/1aL1A/ajTCxBmp9NTP0M4YTzXajLt2d4iEGIGhQuqs2JjNVasuzzwTN
TlreGtbr2/w5sbFeIXD9Nga+ozqQiXow9K1OsKR6ZV8CEyG787IP1IqaFMczxyaFwTg7F6e2vDDG
76nxi32k7TuGE5evn3l1XMW71Ul3lzkcjTxnyj/bj5XOtSvtFdEeua3xbcKwuFXxBYk0thPcyPpz
Zm9VPOpgabhQG1HQHnoqq6fy4Du+ajFnjEmF353U8H+yKdIn8oZsEsGfC1yxYSvo5+i0uAHuxJCQ
eCYfcj72kKQHoqBn4R4dEEsBBG0Ybwv189ogDX/IJcJg7gGORNq8I0fCFuEUaGmqH2gtL4WK038G
qQgLnEs8OuTCzFUY12bKJURwM0HcfW49pH/5dshC1zXTbFs5PfdvZs6TQeQ5sntWIV79nOghptsS
QVmdmASUvavQHugl/JrgqPtbsq0XRaiQaMJhYlKBKiqY245AxM/DeSCsw2k6i9im4ZyYlNQikGZB
UW9FeKBk1baviKwvzJVxVKeGAgwCvnPsAizVqHaHKhtFk70FGoibcT3HMORerjqnXjow8Sct9Ik9
GSSC8e04mmPvU9TusPnzy6sFvyu9mKJCwpGE5pUquvSpsbmchWpWQI1In3RBmKb0PNvfcfuDqMKk
LGfD3verOnwOlbnKr2lxP70qfVySO7pJR+2bHA7Wf8wHzsfS4FPkFfYtsfdwah+pOZMalgMEUTpb
5CFjj9Z1dNBLHli5Os22BBZZXkcz419u98QvPSlnhqunr/xS+F8fGQ822AN3LnqbaX+ItyvN6WV1
hsZPdFtCRvaUMxHMLWBoU96pTE5fC+Gj5UBrJlHkzbMG21opgCrLTjxCulFIbRC9l7/v0ujqTYbO
GF+1Pb8yaoWHFUxdmOfechGSTBAa8O0DDiAPXYYW2z/3JMybnJ2DVFukLYIUeAE5bKYoMq1yd6z6
dBdaDMgVfUETye4q+eIGkZUAnyx35gje/gqXrXOVXoMzUHG9ZyFU9wfZ3OcD4YrBzB+p3ZDnSEiS
ukh6t1fHxoTEpgJyoXgMibige7ZkXiYkxQikQywtGZNm88+wzEMN7IR6sCIjjGzeK83XVzbl3HgP
jBjq0Rz1RaDvOAKclnG3H7EGp9Kb/U5CA1oKYf9fPfvVKgF3CjaeePSu1fY/3T5WOJMwZdMaje3H
/wai2Sst54wCA2X2lFatT+1aZ/NHjXirT/bdtxB/DZs0jcMzOmePRGsyBkF0m2AauUGVWteTuLzM
HFVsiZol+rMbJJKn5TWXIsVkCt6TFrMJ0Cv6FQniylFwiKap/BsgJ0FMmWYSaMS3ItqXge3w9Lse
0sAHYMcO96rWw3As+vlz/y0Q+8uAvOsBjRWFPQSbHDTCLDnN2OfF2x9XymveizMoSeHI7HvYVpN8
81EPCVasFfFQPL1NvT8bGYadxKwUnGZXhCtYVWX/eO67Yvx/H1gSirhWNCDsAW5g9mhE0h7l+V6y
XIzemJT0gYwV/Sof8QKv2U+e5R/w3p7933oCEIP9FNwpoBQZHxsJxCEvB9/b3ysJkD2xgNkHVu80
jdH+HaUXcwbv4f4luLeFCke5pogd/s+qvapVA/jSh8HZOK7GxSvCOro2Y1mHeHEduzJpl2eBOUW1
2xtD4wlHwLe6EIFCilomod/VY2OpHnONLdTK7gREzSBjh2XXIi5i48yhR8dMB9dJ83G++11KqrCW
20XY/v8va9obKnus+JQXdx5tzfMJY7yHuwRV6mp8Mzvj9BpLVvSzxKMV7edBxnSG6aJOpH89ZPIi
1fT33JjMf3YJp2WcObySZmzETOZsSdoGlmWyrRP8jT4+9sHzGhlrJYjdH+khMAS0AiUMzVQ1v4uV
BLWIt3BnSwlAV1NAHzTl8lqnyk/rdSN18Q3OfkXS7f0mWUtVyjGDM7HLM0q5rybRijGe6VjFgcLH
yA4775b0rK7i85RW3jLel4/7+/8mvGmZdqXmR9r1WsnTT+fQR/x+efUBxElSadM3k7V5CGE0CMgN
FveKYk1W3FZpwjL2OX+aRx/BB7M/CtDvpncPPNKSg4iqMWIueKEAA4HrQXYQUz9MsBynrLK4p3NK
WdYym+YAYZydy80Tze6fywIDKQTVx1/VvRG6pT6unwH0AK33/0CT1jP3E5g0V1X6DNbwbz+GaP5t
wTP7vrmspyGWV3vPUWa0b0RN2ZNOCO2MuqpS5FkXY/MzX9X8sUNYLaDuekG1xP6ktkVJpJUAUMU0
8f1Qy+fDaC3edIhLNJ4rX1W49ntDXojhcLVZCoLoPof2Gg3B2BGGyl0jvqEWeqcF58L3ROIbU5Y3
6FFYSkRO9zdp7EbNpoOEUCPW+4zfvPlvX6y8ce+RyHnMVCkL2S23Qp8fjDxRVwoADudGcl7b7bbx
eZY6kMra8hlkCNtEGov2c4OapCFK6PLvDNsSnT6GqNRzvmR0ygJz2Fhnsmfc2rZFUPuXsDQi5/u9
t3WOrxSR9awEPAhjtFQlLCY3mxIngzLUAVEdZ8snkYCvIFz+1LWTPulcisAug+DkOr2DJUuU/E6p
yoyBVBzgnyoXMGm67O24pnrG+E6Ae6gvBAEP0speEgth90vfMHtTL0+9/R3zioK4A6PboBJ8xej8
FmhY3319/UZksS58PhFELmgesBRZc88cy02mocyPbQNmqkegRNJmytMNeHrcn8DATCkDw3z4jYQQ
uXkzlw4bKxsghVOlRUXSdP0eypzgntmXQJ9kci3+kY+bS/tjJL0s0wuirYoe7NgxIObTJ+0MTyd/
4ZpaxaHDCuoN2e4smST3ZMsKWIixqofKQNNJDv3E3XL6g/NM1DRj/nxj+WcACkI+KkhGZBvV/kxg
m/rydqTgNCmz/uohP9nXdYZjATv6gHSXD67AzQ3Lp2QrVMfNV6gXqpUepLtjrXAFEaEIs2dSNT1q
+dQOLofS5M5Ct/hcYaZaaevKDZbHTA9AuloYxnJXDpshcuXKu3SWppDQRG1gdsI3YgZfTc4agJ11
oobPT7LU/9blO9+BiNUuPH3LsWIO8gGEMGnbSfTPJMZaf4FXGh5IVp1Gp4K7H++ZfPjEtGllx08D
vQNyUo4DR5cnnU8J8CKxSsJdvRmQJO//2o41pCUurvTyHzrvzvDd/Nd3wZP+ltiaXli6BdpUG9so
lYzwhhJlmbCIe2y4Cnhe7G+/U3+IlipFlWDFNmBldq69hlybxJ8tq+7tYoFolnk/qa2034W9sFOY
YRRBCnVioCAPA5CgzP/iV8J11WWcHoNPhkQNLcDxZZpxJCt1nv6LByR6JHfFBn+jSH37XKJfR1xD
c8ZewVO3OZ5Xwl3X9MlZeSZ0qJqHAXzsODty7yePP6LkCkzx9xmXX2a3S9wXOUgnYTiEgOJmRgVE
Q0ymB5PEknUXvdScVoiX4SIsuh10YgJnAHkeaF+Br74Wq0/ebT5zjukfMm316cGooIeDPSOLNL8d
af3VzSmGQBR9qEXxBSxICzJujZuNRe9gpvcxSyr7VKzgQFTxz0d5jnvQMBLQ6IgbWPf3dYlRdKwr
jcEKzpZd6uvo50j0D4130Nd9cKhYcv1YFF5v8Ic9bltxapY14F/A4jEZ2F2UHOaHhNhtG6M8R+om
cPHf1WSRVpjmLVL+cM2t9bNKmHRf8eTDDIKXuV+0h43+VE1FIUJzW8jKv6jyN36y/EpYYq5+f1Tp
eF2QpG59nXIQFk7xId+XiZr8mjyZIDYhPkyJUL91zMb/vmapCPAfXRfB4XnR8gvNUBQs2l4SXKBH
+cTbnx7SPj8fN6M0OcEwZzcMi5v48RKfEPi9J2oK0hifQX8LW5p9wUrD0rJhigYB8TWYOFRTOsft
NcfJwLDfOVcngV4RXV1fyETc1qayM5JAfHJ8hl79SXqk9oA+h//oDPAnVlyGO0l3+Ys8JKIYJ1sD
K/PqUtrLy9B777k4Mz3N8Fff3UvUBz5E3Ea6nni5pUsPx/L0AkezSw+MwzuBubRwL6nKK4HJf/sQ
dJzf1cYw+m67PN6+uFvee9UusgEDeugfJI8aSMDws9LP24pIMSdj+5XB59IkG5eaQAUkGABwHcpF
QvqiX3vCl+yO1Vk57HQhTrULXE64lty9XSFYJw6n+H9Ut98klmKaxZOEjgEcBF0EQwbXBjNm7IPv
/vjrHPCo/xIhx9UzjqZCRPrYes7tzumn99cIU/ewRvCvTD4035oEylz3miwHIVLLgN3NOPBRWZIp
LfRK/NIztqPaECPa5b0mykgcF9A29cU1e2LFWzyW531/ZjzpoOW6MrVfyloPsBoGUC4GehecSpxD
HSA70+orrzB8qOZHB+3MoALp9wnOI1H2OKeuLfKZVgCBt2QAwztuDv4ohinxUaG1upPLl/MNRrE5
gXaoE+Oyg9ne9POGUbpXb2EdwTlk5ZhtHQhpa8gAR7PZY1GTZMMO8t2Is6+W4OUbhuAUVqShqy7U
lJqbBFfBOZ87H/H68Ax0hOm21I8NK2CD+XuytRVWFyJD8IGPU89hOV4tlajRKjZ/r/DUu/nBKzmD
ToGgbqIftnFZdGclTHOIZ1/jt+E9talYNWbbiBjE/xVRiLOpnKcH44QiFHrjraJ9r19hRAZlIJyr
++4mS2Yd3mXVRoG19WBMR5dVqfgOCvlum4dxw2Q7R1InAPKhgwOxvp83obBTs82/I3W3kPwKor4p
mGc8GLGmjSYs06SKyP6eGzutHrfn1TR9d45W/s/eFYP69xiU/uNOK4IGtDXPGkEjHtZX5sVwIAa2
9+rhj8NlwK22i9f3AImholUsE0k9d0xoHuiRwkEW+BWZ3DNUs6Iwvit5EW2C3/xYvhfVuMTXsl+v
7rOMg0p0oeLMi2b0qzHp0rHdHNgawL9fg+7A1rFqz5B3UW6w3WkXTCfr8HdvvYtZMCJ23dzoKhXi
GH42Len8ZBmMiqBFzlHso7PbwVoATRSAsCX0u7egK5oXanxvBelaxfyQ3BAOoaDrfMG2jOrhLac2
KpQYlt8lx9NEKDYATJkXwbcNv6fbZPoIXQljAZlQ2V33XWrpn0pEfUZwR8Fck9i0akV+ioTgw1/x
ey2LMKh77qeNl8QYGmylBOYto4QRE7mniDtYnk3sCo9QOKwheDd4Q44NjqDUdCC9tRFee5sbW4ZS
eo7crCdwi5Yi4OVuTlq5sgjKS6xy9hMRkEZe+HOihzzHX4cVWQBRigZj0zaXIGA/zr1dxOcXkxXO
iCJuOm7OtNwaxIlR3U4OibLNnlrcT4B2X23qMVAgSN38HMjiheakyTI354c+BFMKQxsVg6HPaNND
fyKcCacYB0NX4F8oOCCOIBnKad6tBj29bTh8grlz85PmQy+AOW3l0p00FOKS4XFpFjBPSksSfJ7s
adDRYD0H9TwMxmbeIyKBilTinCIP6JJ1akje1xAqp47PczAFI29v+NPgoVVgEyDEcTfmmu5yKSTT
ofV55HAowUkj0Hg/MW9vBjWSld6IaLqUbEE64+YAoFm2ztV4Xv6eVY9h0Vi+eDBWhTMfbwk5fRhA
YS3BtBfs+OwvDLeJsYikv5ld9FziYwn6NBEsTjEkks1IVxf/WN4DCYq8zPLRxcN7S6/ah7j2OXLo
gBDuhviztf26lTOXjgZt4ZR9gwSygVEUW94pU+VPQYtODUAJCkpYr2ydjeD+383KK09X0L3ghviJ
R+yOhyuCmttPjhtU/E6nz+MSHyeCC/p4pWXJhC4lwH5dJ6ainBMIDGrA2YNVS4tqy+ysy1BlG+sC
2rEoa3xGt7cDxW3NBH+TKLl7Fe/3ncbPu4XgL0sEYcRGMvzj94Pm7stKxxJFoAg8rUUOooXUzNww
ewSke3SsQu6DLNlDUW6/F4+7y1lIyG+m6ABWSlY65qqzFCuvplL+Y+GgJrRMVmRMc8sHw139zbL4
BsZjLkT+yA75Izu1ps/DZymwiFRbFJ8NPl9Zbam6CyyaDDT1JY2stFj1Kk6PzU7/8IGDZnbG3kkH
HU/tG7cvYrrjMWN2lVNeKVDkeDINZFD9jAMUJUaq8U+njjvRxZqGnJv6rHX5pK2ivCiXSFlyzDnR
BnjDp0CN5joHz1VEBpYROHR/04AZqjkgTdKwM6j0In9a9Ow5KtA/jylTxwlOjBE703QVuhVraXqa
QDqPzUtTUmafZSkwArlyIXJ0mMxem8xrF4XjdKeeB3Z5a5SAmepxZYKaOzhLrrPQVKNzdm1Sba5y
uFUQ0RsFkERl8xohtgBrRz8zv+zrB2757GTlPuWqD9w+vjx9LM9Z1kWYafZOoEthFzw1umIPwViZ
CddbU/UVy6Y5JkpZ9C1wiYV2r1UJBUTvknBjMP8McDPEzCKdZCr5TIjBb8mU8C2+LjgysB9KqyHm
jKDLmTTcFQLvrkLoZ16bB3Zm894ifuT+/b6YSgHKV7ShGzvxW6wOqikHEwwle33Q5rEcuE/OOMIG
kEWH7cLTDCXuUwycN3mwepzbOidmMNRjq41XSATv3ttZW7S2WTTsAxvvcE4kObshxYW1UytYMSyO
5QpRzrQhrJz+FlIa9HbwDuhytFghaG2MKt0FJiC1xmwanH4pB3o0/WAtLdD/qiymVn8PLqkIok8m
viPEcDXercKquJ4eBlef7lCzHBe6S3qEqsF/kXXf6qCqOis1Y2X6/2zTFakfbH7IKutKbeLBmpnG
uTssuRqhMv8Vk7e6YgEoqRsmfvDclIVeOFk5FB+kvnJuSu7Pm7WPL2adSnOHV+aI4DuF+EAr8wo4
VV6XWYnNAhQ95Ng/PlwCTaHKmjoLbvXavdAEqNH/Hel0gtFHFxxPYyFDgC3buttC/kwVjSnFtPFh
6l3bDxq8kP5APppF0zDudZIvgNysVqBHKCLxQbgP91SNjcqGCBioxMskxpwLBYGqUKpfotJiM7He
b2Y1SY5HSEIn0gjBme+EYJiUccC27F4AmUEjy5yh7qdaPAfLWlq2MIX2/FP988Buscx/D1q6o3FX
q8vTl4cJYvyR1GotzOIbp9UYEPebrYW68yEEzl+H6QBnw4u0PUOxZZwXMfDW2vUnRcSfojpL5tJ4
wFYcJKCbR3DUs7rFjbwHmbTN9PRGL2Vi0V7ejw0vwu856Hwsi2cOwjHui7c4qJkGyCDnvfjLS2E8
CbTPK8bK/RXRWR2fyXBvJNGBUiTGn9fx9tlFdSJ50QF5iu0izTpLJlAPId5mxaPqpGKNSS+cBOvg
uAbn97VkXilsQEBe/8/UjIvCcIwW0cFTLR1p+J75jibyIl00OBiE6EefUp46nB64WGVQOmgijBti
AjamxZ/CCsWUCue8LD3yH6tQgtqOl4O63qRb378wly0VlRrGVxND1qy16BHV0xq7KwqOJrH1UBsW
ku6GdT2M/6YgduUXYgWbDy49P5c3fRuNpY/XXggWXR01stv6HxkzAXTRQ28NMbdbT9K9PmbYVw30
7j9ICjR6RJIXDuHbJvP9mDkpQRdgdK1yLAq5J2pDamT29IPbCKibRakXBCw2PxAc3aN6rYIcWHKG
83QZ3HIJMg6QNB5uGLXXG0ewNdONM0RxLzLCB+3pl7gWfHeLhrxmXGDqUvlJCaKHtOOBGIgPPdLe
/CnnuyH+6ecf9FnZ84icFGpZmtkuQRGm22BoM6Cb6AQAFJ/QnAYqZzLccaxCRwUGWuSLMggDUHFT
GRJ2/vYOq/IVB38IwUu4EbBlqKjV2/vifdWRfU6y91OYNROefWlwEz45Ukyo9boVIcD1aGLOaPHg
AYge/IGHic/eoQKQVGeQ95jp4cRj7xp8fRlRlL8mtZX7Tise1YPfXVyEA77DfO+tHWkAAJN12KWP
bZNoAg4SB2suknY6lLVwMHGnFUcpvyY1+EVvobAA+lTTGTxo07hZznTaMwIszN9ii0FssgMgcTqe
NxKwkJoWmg2GCKNhWzeO8rXCwbBcNYkNC7dxx0ozPCLIKuzpIKh8FYPiRiYxAjYOQYUKEl3V5+ST
wPMaQbEsIOJo/zXdgf4risABBCAtvLta2gj+KFEAK/SanoxLfvarzXOqfOAqAOtga1CwmeTyt/Jp
HoolSpew+q44hGSPSrRZByMucBEEs6zuJ1GLYjVOFruJLLScmtRpEuREl8TkuXAOxp8ubQbtp3qk
YnN1q0b5dV3dcPox6z/RcOS9EUwQKYEqchxaVNEJrlDTcsUl9cmSUZ26nuXOyBmpsgUpHdSUqMJG
VDGrRqcBx7Dh5C1qG0HlFcTYI5cNmrELsFCKuqjMrvRKfdvme/EqYZzlC8LpoQAFvBxuW7LAF2GC
X2A325Cf0jFc0szPf+dtl1Eb4nDZWpnin14GiaA/kawKxrrKdp+bNZEmMi1m7ZkG56Ar5u62B6Gf
iU3ldiA/OkTwTNJQ6AUYjZEBxZQt4HwsUCVXd+n4fcNc6vu+A5aY5mv7mFdWtjaI6J7FjK/xZw4r
9IACf88x7xw7XebaAGS2+o2M+rAgChHtQFjjeRhWjVIw7QrKakUfutI0w6i5m7I0T5N31sIabggE
e3QXP2tjoVvz2JNLO7dYbRMIf8qsWKlc8luJarhKDtsByDVyObxBQAU7+y/eNIPmYBGbkxhhkEf2
ElN5VWpzIAZpHtrpnLPXX6QLxTTWGR0XQ2+4BlRzWu/5WgB048PpN/vBHtH/yQ4dLd/AgnXyOKfv
/vauedubzEXMkiDAdI41FQ+CINMR4ZOmJbw05PNBE89GR1erTr6QnAFfjDnrW/EjeVRp9zoL8nxA
4TTEv+P6/I0ozDb/pzY4Y3Sl683V+h9roJtSZgoCs/tX4nGDvB9g+7UfGkjOv9jbnTnrzq54+YCo
3Dl//5Ffsb6TXdt7NCVwlYEB6JjxfTVOm34RME2WaGBgcBCdmWLPmAotB1MYyw1sTg8S3J/DbfFq
N4jZ98qJod4XZnzCJz3G2OVBDlmIO2UGxV5OntNYtNRPphNUPZFQ0MZIu9YVDqRDjOCWM+dIH4E7
f+kjpBhIrozqw/jNvhstGWv2JgAEMob6bRK09Z/koay/PHZyvp06ajW0a7TPT05vB+dYl/hCGAGT
LBJgqm6jtcoFUuD5WD5MmkbkSptR7MwXLVfaTEDZF2o3YhtIwB7cHY0UFc07+NjIlHpIeS/RgsWP
MgkU9FCctotFygLuGmD/SjMTml4HQlbyMCMYRKqEYVSKjYjHqsKb1ydg9QZInLh+BiNZGLwL4OQd
Vgkr3MueeNy8i0Bce+9xrhH970reTYtMEIvgCDLLtEsNYhoZVXFqEutzqln7oq9J+zeRjTRIkA5r
TKFZgoLyP/7fC4DsZSRxdMc8KG7sBX78r2KXuihFpQ4jCACBbjV//j2qQv4sYFUfeSnj5nS8h4Lo
Zdc/xr6BlGA84YdNH09RC5D0gcPxUb9Qj2S3z38GS7gkttKxurYDLc/b/cHoUguW32316eHd8ulU
mK51yz4qB/GLusCJ24fmj52NNGLaUDy4RECVER3b1bDOF3bK9vbpmcOoxY8H2pIcTUAWXmIEj4Wj
ypX57OPhT19gaagl4G/fGEa7efKx11k8GD/E8htPiRA98uk3NyJNYLV4yCEYgSzUmdXgSFBdjoCe
Q9dhJerNUHtEEGedXuhuWO56sfUBpmgM6WCk+ZjLw8xCtaypjgQu7r3nl/tvFgFK+Yceojz7qGII
jizeyFfV1sllKcFJiHNTdTIZ75/E9fMSIzzTlwc4cPf4qBGOIHBIuQcoWt6yJxzyeumDJRKYDq27
nQ9TXgcKfu/zRue/6cM7AkhJDQ5ncTpOsFEGkiJjUoT5pGJ4cdL+lHEYLMqetUgtZgrZOEX0h9jT
o6AygUJJhLQbVjLFXKhYFa3NlROzd/Jd+26aC+EH3Rr6T2kQb6y/zLAWe+W0rW3tgrI4efyvqmn1
srVIDyYOtxZI6LtA4DqyWrG7u3FFYq5Q6xgYECgg5JWaYsc1y8+bx0uxug+JVaFSnLJHVMGCf+4b
DuUu7yMESA0+RCJvnLtne9CxrOCL+pojlMu//Y+ddasSgZHPd7D8Xe1uTUENShsCYvb69hRmOEub
zWWClUJt0ll77WPQR7a6pKxL180FGg65+vygRgV0kA35dkAIKJr0JBfAIC7kAXNJpW28CKuQm6Rk
TmmAV0IwoyoCAFhnpN4UHhPn4Xt1BxjGGJNisIiZ2TJGjz/GxlvSjjhDEMbpzLpCDpv90ZYFf/PP
a2+Tgxoaps1vWp7eX4iAD8o6rJlhOKHbBq3xEcuA4+C0uoLmUQzftJMbjI5kcSWzJerRuLR10F1P
eaTQdyrGnLWWkSLME8NOYusmBbmuMU1J9+wG8HJ6Iq7o6Qt8PojBo/ZkzqTolOf832Ihr7DU244D
rGVCpEBygf+f8px+6ZImKYPw9PH4qtw01ZJQBDkr4JxqdcR+Z8DvDhaCKKamFR52NP9HmdmBPvyM
zq/RwXFzQ8d/8y4BLKgoej58qSjC2bcy/uCzKLSkhhu+LW6YWMQQp27spA1AOyW+MBk2o2bSGXAA
D0VUP5lthF2gTJoBsCulAW5SEwaelTNs10oB40c8luowrK/eO3U1nq5+xGPDNojpFj6+8xb3nz2N
KgmgdVKkSmHdJRFrT4EGHZz3OlFrTABXCHwY9aJ6konueEkz3Kb+4mr0dxofYxGtnD2hw9fDQM1S
VEI/pybLR35Y3fFjbOSCRq34fdOAhE8y6jTAeXtgJt/XLdDDGSx6c1Xi88+N9wBh21PtJeSU+3hl
JwnQKyJx/XjR3LHvHh6gY/UkqNIOn1mAStPBCkqgjE8knx40b+CQaMcqOPvxCAGmKw+LnUub5Kg3
hocXiLfRcYAEynu95MA5RWoq1PYcSq0+W91VfdOs40pxG2906FDE49su0swy4Uw/I9tVLt0mx0PU
2xdjqiW/sRSobb+Atm9t+1AwDrgNiRQdYSl4uDXkULu5U1bsodvXuJ27S/UH0lXh5QPnVFjrtaKv
OTGQV0vbBimGHsesw/1l7oHEW6zpQ/8WDY4C5keFUlWlhZHYj/A+LLqI8EHKPbs8O37bxBoLwK9t
6x+401BZV4BadQmcdP4ZQTUgHGcL6kxBKMOTNd+KzzsgAmW1NiXlH+3MaAx/UWffjLmjU7Lp/rZZ
IeHzzys80NvW0+d4tVxVp2UCk/DCANkwscxb63FL/UOIbJgzzvuOZcTIA+7UTwBEiDXeLYoCoVuR
tSNI+GGXq8XYpnObIX2YBu/JwACeC4wMM0KUjZJ0ZJee7a0vN53xagvbXkpWV3XgL6t2JsK7VUyw
0jPG30sOszM7qkR3u2xJbUz4bl/ZhxSSoaoco28qv99+LKOoGQzCk8C2orF2A4uBYxbngaTbpbQx
sKeHD+2dOvl8IL4n3yYBoBydC0S/4BZcpw74B+ml/j8RqrmBmkj9hD91pGmOgE3W7HNu6Dy/jl1f
HqcWaYdDN1FODjsydeyami7JhzM6/FCt7qLIwcg1WZbSRQQuHhKnnOh1yPYEupjMSglv5N7vviGD
2xb1NPNWtYGnz5TpiJzVgYWzwT1bo2oYdf3kRUf7odzSUGm9910L+6HexrN02NRgG3iG8oJZ2624
DV+/HyuqFmi5jqwzY8WPbgwhPebQIR4ZJF1I3+/6Xrnpsl/veWO0v2gdfsqVJGLrkDhkMn+kTi0T
AGz3D2RPQfBs4saBQfPAWqFCxgHUTkihntN/w7PCkHiHmWNZLTY0qee+LL+W4c4h4kdXX8lIPGiW
3b/iTUyFOV6iZK1/UXx7A8NG+1Nu4BLc0QL8/3FR5/0EVXunXzUZEuT5eutUyS2gZvHISVb37r5c
aZ/JotFkfFEeHifmNxXF7Nd1hEZ3FzXyy2qbu1KYlDAOxM8+t/JqS/d73f/ijEm7o/i3CfQm2MpS
QTrVHita2/qzrtGp3r/PVzJD3UevULQdf6Tbjt7s1wi5N3Rw7jbQCUM9zaQWYJKb5O9+7QpL1Tz3
ZL4e43sIr3LwtvZTkr6ZFXd1iuHPEYi2GGXB6w1Fv/HG5xwrMV2XpPyLnUSF+fntl+5RDaJy4+Gt
+3EVe/4GzAqxsyfanjkC4HfkPVXXDdhlIR4Gg+He09PHSAWvbvu0BiEdqBEPTfbIYiUbBW1hrWAT
qPn2eVvi5AnI4hBmgJrnxzxR5ik2BxILFg0wnyyW2OcgXDHOiFINbmqmFQ5l3Z6f4Fdp3iULnTm8
1F9mwlTXJJ+0sqnnDPqW3qHIN5fHx4g1i58wagvh1MQZ6khmJqszEuAz2wFIplZWYX2iEWPuhAA4
lB6cv3kbiSMKZJNIswsqRNZiJ7pH/BM84I38F3o+gAJP72wGCvgTqYvTo734NTLnfmY8iGU4yJti
pyYyfwsVVjxq+65i0iVyppJNa6yBrZBhgYWktN934rwTTpEz3n/zx7+Q5XAcpLJ5iukX8j0AZIYb
a3+pIaAuksm2gOPT58U5s3DSTpc8J1+1iXGyeqKrrFigoBGYIpARwhmAOwUHkuVkH894zQIt/MJQ
XYOeIiFBmLri6NH3HexxJM8v84yg/r+NTFcavVN5f4f31BFmX5Vk1Zo24PVPNqOqE4qjQXfg4Pml
wlSXVKOS9t7Bgyz4M/60sarqh0yMeDKakB1y79W80OEPZTVp0aqe3j777F2ANOEwPHZTPPdiclQs
u3NPQYcawzI+T8aqaEfo2pKjpYfiKw1B+AD71WIa7gIoEkIIQCumkcefH9fW6MMoyE/XdHAWD9WK
7SkoDZyWloM5KKwOhnlmGCgjWzYXDOcM5hm1K99hrENpZ9h59LctwX1SAHYJrxCY1nHSItJ3VZP/
Vb0lvel+mBX8C4nrT+woH1m/95A7xzCne8kog3Q3AwBrOhKv1UhQsORFTZSRq/b5UTGk3wnmhnm6
VbauyAh4nDOaw2fDuh3AbrhLWhGLCEJUYoPoCzGXe05/1NEgY2xxC+9CpZpMjSPpDbDGaDlzMK+6
MGteoK0OOovYzhi7LTXJa0849tZK7bP0BfkRqrNyrDg2rWdhESjF2ifKwcJFzW+m+V5GSxVEwZXX
mpGFRbRS91AUvzt2GUeGCp/QSqTE7ixWgALOBPQzDXMbPsSFLEDQzht6tg6tYWAscqCqwp5PrRh6
2N8LEvLiajc49Ks4NqsofARSIT2B4b3sg5q/fzPdjnDgesd3DSca/G8K23upFGeh+V5w68uiRISi
FMHc1lHAqJvQNxvcJeysndYdJIHV7ZkV81vniNLtuwPeZlGiHV4A8AQu+8nU/1EArOciSBDlkNKc
N+BeAjTBKbXM9WO5gOTDTzbC4Hob6ti2D6CielgAQza2GL0TbkPBcHmyYDT3EPXj9qUBfW//jK29
iRlP+DHLKwO8/JtDwSe8fhu/qKu9fjkBqfM6AH+R+i1wRxR3Q8x1dTutFoTf7SQnPbVZnjnvlhZe
R1VxR24mp/KS01rGKEG6GLd6uXEbE2HrBOPklKxOPjl0YzmngRNIrD7mnFdNBebtaC3ix5yeTIjO
G/yAyV/si5rjXA62kT4iGxPjLS7CrC8WbyAH01CJMNcSn3GsgEnmTRGovSsw/j38gmx5L5aNFY2u
hSl7DfWAPt0gDcJluKUNMgNCIja6NOXgV5YU8qydHUd5yg/ecj6J3Uqd6BI5QtVsgz5W4NZbKaVW
GjPaEnYF0fnzrDiE03hX3jCAQzzmk6FHAHFa+ezlidhWhBsk3Nm0rmmDeXsplWaGHO4vkh7AMXqO
Vk6X9qF3ce2dNpIDduO9ogeKGALzZbnPcS9BmaoiZOjSQFB7WVU8BX/rWa4cpKTej4gjFFu5GbYr
DchSa2FlR2rKM6CmNot7KzrFBbnPOEiuLAaqPD71ijp6t4IF04rTxbsjI2meSfNFf7YqTikBR39P
hSEgbwcOdgd9mUy3F1C6GqGt+kQBGCQ2kMT7ndaVHrOcZ8OGystT/LAM/N2506PApENLx6qLi4N1
VO557jUGZfwffnL6yUA8d1pmdJhMbkA1NNIps+MG1sE+UKDVIz4K78uZaGFZ4JcbNWI6+DkDkEbj
yTGSm2/HlWmo3JjrImvrkLTP7ymHMFJITltZN/PtsxE43zmxMl+nNySkZe6ot9IQMnmSgFsLZx6H
X0R6sRoHi5G6R/zD69Q0BAD/57cQ2C+u/h0CogNwcR9Vyt4WwWw2YBnI0SdNJThtuo6ZnJSIwisu
/Ec1p1gPtSPqoe1YTnqsqJm2N+R1LOyoeJq+LOtqBKCtx1S1o/0NS2cHAsrVSG/SKw9bPJWUNEJc
1eUkhOKT/U2nOXsJRozO+xMjXUvAgyyOUhVyHubycEq2bmF/uwyPDP0QEyXNe7HgV7f9ceW9tmIk
+Jjl5UszPbXpTK/SHW3zDd+u4vYeV2MOUt8DKnMZAo2Ru6eYp3C5isxzdszNcbc7eNXxeeoCVQ62
m9NvuGiMmHzmulTR3GukMWKmtmj3CLGJlF8xrKDhbLWeiookECPGQKoGdENvhc/4RnqCVeEEU7iD
JjxoQX3H//2zzVO7FJmS+drKczvre37meFYQ5PfP/qHT4yOveFiqFUA+N+/u7wsAryStd1kcRXgL
0Ko8VK1kzlGIDVfJsAqlVsbRkSCEg1z6DpQZl27S6hMd8GtqCxAWzOpu2/9qbsrhe4Zl6xafffee
ULZ6bamHgo26zgHyDYZs9B5eVJ4A6IQrzXczBI19GwFh/6kMH2pfh14kRmqFT/YWg1vsct9h/1oS
F7pUXnpw8QTLAOYbomIQi81QUtjXeGKyWv2X5qvFJsdbMZXS7SxOTt7THVJ6I0j3J20y2P9Pgkjo
S8CVgpKBhZqUHoiOyk4jyIG2fEscmcvEqo5JsIWbJZp1kqO651M4sStMCT7dGD/TUWeWyCresGvl
vV1swGIdTHgN0fSmUaNhQbwQ22IWSl9B41Nurz/DwG1OCrPBompX5b28lm9fzQ0ZuUjKUabO6iIe
uYvtCgS5Sb03ydCerP68T9hEFe+Q8U5fPYvOhE+oP/+jBcYEoeCEuKq1rT0ArO/+0lxJoU3+AweR
Ati9vPTWP+xbCwBBiJfutJDEq0A4wyy3wt2mbROyuz3V50Ee5K6aGOnNX14Eopl+F9qBKqGh3MzF
YzguLWnrlA59LatUdlqqnI1ZE1gZJw4QOOE8wqbCBCGYb9LdyMQ1b4cTYNDJoIvkBgwnisz+Y8o2
Dl+d9hxP5j+uw+C2HDA8jZfrDLOUjjpD8jt7VIPNGr1SWKv3V5BJV1kbnMjpOjD2SHCFhRM3mdix
IerD7W+7fyXTLNjRJFUC9zRZ6uzlTFp/R19bd4favJ4ssY7NNbTE2Y3yyNxAfWjAB11lR6aEm85U
GLZeHoxy1dV/yUVz3UjTtuKw0N6ve7HKRQNg/pMI4mVw539KkukyBshaY+4I5uBOjSIUM+zGpFlb
Y1x+KC7fQUjE7xSXCJOVibR5QkojO38oQIiScrqxpxPPzw+gi6dFxomJjj1XSTCXPwBBi0eZ1eAx
f3wr2atjiuBghHvfV61l8go3EfuUDHR0WQc0QfunmCJlf98pOGD7qpy5nKwASoPBVqFnQgV0Ro2S
rg8LjQ10NjSIAVSGnlXWk/l2K2DqiKDouSKnNP9Ws53yAVfA8l2swxW5Bxd1nTADNoja4v6uf8hj
w48HorkzY6nnHlR3X5aBl5sTJSGlA4HbP7dmC9N52Dsk5/dANkisLkbMf5T+IG+xfwVMhpuwmbNA
sHP0JS7bZX1j8egMSyy6F7tWgksrmuQDrjksprxxiGLqxoOZD6n5Y7ExG94wu42qh5yqo25p/nC5
cdd2Bh3aUtQPTtacR/Zs1dMy729/updpjVAKQioWOWJNWM7U2YNeVBL5LnNn6NW7EHm7Mf+fxdaF
peX3hWC8Fg/kzRxzIrq0IhDdnv5ZmqZX+KBtewdOKk9MecfSIRSJCzZLJTGBTzm5NkChJSsuSzEr
u8LInR/jz3stzv4JGN+YOUPN2iRkdcRGprocnXyTchMqmptnHlsSX33HKXc1xrW96H/zNzt9XHPR
FYf8SSsOcr3YzyVbzpfZe1XeKK/D9z+cEFKv4t2Z5AtN9HW2EEA7ceywwkkQC9oBsVk47N06sSOp
T0PJu12z/7bZAzByoGvA03IPXV6kuyaNeZv4GAWZVmCFAO9x1HFvcIx/jo6rm0NHDvU/xfoG9orU
GKqMK0JVz1qyj04Zo/Kw+VqftpRkvQ0FJSHSzKh3R7ZCIqxJBna1uvOSGym3zQuOZpMIfFomjJ0v
h7iSLq4vKAmxQ6yGyyi8CmVnzVjItAa6CQUCLXSgg3cahwCtG76orf2Bz7T4WY7EUvMmyoBuhpQ9
ajCmWcmj/HRyJhnvTf6aiFMnPq9ypuXc1VM3lRE7O8UwaeMzdilgwuIRQ3y7JmfirK/kFF/3VT8p
FH5+hnC53FcyuGZRC2wW/J2RV1a1+GrYUgtJIwVi9LKJTMeyMYiU//horH6vOIIow6b8KoVjmQu3
7Uee4SsBEZ3Ck2XgLZcXiKTlFt9fGkmJg1WaYCu6fIgRtQ3GbS/wsqzzU4CBvEh6j9GK0mZbxy4Z
Fba4NuV9PtiuIB1YRyLw4rs+6i/v/lPPULou6cjn5V+e60jfMNtU2dwfm0BSY0p3I7yDaIQ7TRW5
rI0RtWoRHNm8F/UlwEdnXgQl90TUH995dV4Q5ytskF7ifCZN0XuJc2s1sak5HUohooyjHoDmFFV5
ZiHsDyjabIQqENRA3ww/wBCOrJe38Pzx8rI6YMvuhxOf9Fgww1+xhngiSLVLxVChWAnuJ6eTRE1Z
gBzS6iKnlezzR60AbRiU/4BjYrz1mIXERQUe/a4BeBRRxiy5vFKR5FnbdjUglF0vaPfCjwF8NN0B
pqbILrd4cQslO5IuxVGOhmKFOC5uFEX/WTSnIVTHtotAPwD+2IYTq0Q1p+fpZhfI9aY9b28UZZuv
42aZnQpvsHgASPurRP3H5Ebc8k2Ds+3Fb9X6ZNxIyNIX9oPlPLZlN2TZeoTlXzqklazGjzrKF0y+
CQHi1E28ZhAAL8r6t4A47jKiBtpRTq84DnY2MHjBhfdgk4GMKVpJ+i8A79vc6YFSPh8499f6BxmB
qdzPwio+U8yXGYk2CEmU7cVOfm89utkWPRbIht9cTthvEjSBxBLy18jpAllkRMDrXrg+fU5+TSMU
TKMoi5ER1m7o/ZowyrxYs6pX7CQLTGRqRVlbnSDwtuEwjkQXgclJ01IxQsJifXKofs7pHaV7NzmZ
w6Tr5qT5ccFb8Rzw1IRoQP+mrq+vQzSiHXGuyxNmwEUyLifE8aR/8/K1pJnmBe8ShdVbNzgXjhAR
+2nDP9eLfscXg1o2fXMnNeABE+gN7lE97PHqAIANYIw97wek6ivKhxac1+0pxoR9oWSzmRiHNx0P
GNPl/B50rrIgGDRw+6OHTMcvEEcBiKzbpL3jlURAGNBLpWCsWi3qgNPN7xQyYjgWu6jqoXvTKDfP
cnkzt257Am+t/iU2loaAV2OLkW1Gf43kO4GWSFJevje/4qXAwi4xxh9Rp29AiaPja6/tcqbrm5ys
uYgzME51JRhPe+VDSQu1c6MR2orkRBoXbo8ZdSiiwgFT1VpMBBbTeweDt8KReBztI2W9xO2iQxHl
dBe6BOVkd0qcbx1/8+Gfi3pgPQZoQn8fs1d9jEECf3R2whTuhBgS99l9IRmL2bfnnOEVVVlKsshh
OGAiW7lYfu2E+yMilikVUE3t8aCdO7MlyXnyu/HYuqYDbh/yor3ngteqvIaLht4x4aGGqv7I1YuY
GYU6ZPtJtJM4QbtejNNdOIoGInfGs21GELcQnnd1zAQtlNd43OjNVuJMjeJ2L38nPBb/FaLtJ3ic
RCC2JAXiLJb32X8kJgQ6YC8qdiH41VQ/F9e6pNR5XuU/aqq9yjeQoOrJ7//SgjBJk9HrUErC5CsF
HrI/V8vkv3UiT/cdF+NYHaW4OJjVbCIi3drY7HU9hgAx5Ha8mXLRS2i2JmMO6BtTMqDbxaGQ3deY
X7BYXLtmytEcNV6ijxUUIVWp5Vq24isDk34rJApBCT9E3q5+9D1TtS2DzxEEApysUsUNANnLc7Tu
LztniUilsWtFaZcyTe86YE2EHxr86KCXL0f9SsN3ooU/1WYlyyZu7PuuIvQkhPAHcMHhXk6CATsF
DfDYUgUd0CHcYlX4HnWCUPuvwH+1BJB7ddQ6smf0+3uobYDJfJXBxp34EaCYI0KgJv5JU/I7Bu9S
wtkb4loDt3d3JOMGNuMOMfouUkMzBwh3BsOQor2pfBk04Pvke5YCu39jQSqJv9DJh8S6AXHvhKl/
T1aP4hFKLkYJe3ZA/+T4ScuQYgxCsFwsfprgo16K5ypUiX/zErCQaj7zKpDLxqBN41kLHZ6p0p/j
03rpFsVQTC7CTlEGXkIzv2rbuT0pIMOPSJHc1omkkeOsOUOMSyikssT0qdQNpM57kU1OUJm3hRXr
94uS6N7Uc/zsYJ3J75AhYyjhzbudLx9fInZ5SxAsrX3JfS9/jOi3OphSOID2EzkXdQhbEQyxi0wD
Nr3+Ihc4ByP+ESWveIJkUn18y/iHZntcrz3ag3+/tuxoI+mBFlG44KmztqE8BYBAlg+ewww0/3bV
sX9DFdaxXyd1OydD9Fwn0grUvSO1n1dvRfH6lGT553PA4DQTZXSLu/cJiHakPW1Mn3f+4E/J+yGJ
d6aEMmu2eJZ/S2eMuQNe6g+abP3F2axZslBEherf/MqvwGubnGfQpKc1fILer3cNNlreI+RdaAF+
dLF83gDBdkzb4YIzkrJVP1j0dm9VXJaqbi27inlG4DvRQV+ccOT8kWuijUnwxzpNrlvVK6Fm9Xn4
A5DEMgDsdmlPN9xsebNFllY3fedd1RoIWxESAk8X2O77y2MkJ26BJjjUsx1ma319lYHPoGl3FkZd
GFyT0AIqACd+uBUVq2ZqN2tUuRuu/p336GWHS6cnJgyys3quiupTOrqF6fDczpP1LTMzqmif1DFT
dxuqabvPuCwhvQp/uih7gqGH7FY0H6pf42IMLm4dBtoXvD8qt2vgDuuCQSBRuI2wfuMGMsYzaCWp
T3NI1HV/egTNQLzdx3vsBDGK79/152RL45ttaCUL0M/FbFYTmFiWo2psz0JxCgVwO2Ay5f1sk/W2
XOzGtN/T+qqvVuLBZpFyauzWCcGO1eyMemZIUvn9dOyCK8+SSR4V80psYgtxajmmMS1tPwGIawN0
M492HgD1QviujWaZTOIAf04lHaGDMNAKCc/mh6d5kk5KXlpc/ak6QKbHmAmHqwRWPCqs/ZMbGx7j
nVpxr3i58DV7WcwfFzHIU61LKjq441OXgOpLH8aHVGbchc5t7qLxqlFylmuMR3+/84yIfTzad0kF
CwMwA3pVrtIZJk26F3K/afpcGUUZ4/2LNBuTURw03xaLYtHfD0jcYWAxQdBMRv6Di5bM0Qab3uFk
JqFSbiWpu8GynzN4FE6qAsMUDNcrBhyF1+mrju1VwotoPtLj0nNOhAA222RF06T44awNd2B8PcY6
iLPvy5kLg5Okg2gApRE1ze9nDGzXhhWktBZJiIBaRA4L/GRPlQU7lasErKq/52e5EuaZkz/JfCX7
L26BVI8PQqc4jhcIVr2GlyliOBXzXqcRRlK9KJ1fDfxV28SXXOkfzq5mbsdG6QS2PLLAbOuTB1OK
M4Uz7Uhio95zXMf0xPj9XR/D4q6iCWEvvxWgbmXoFzY/6AR2gjybY4CwVyNWIsa9jziRaVR8tW23
u0E0YdFfcC4EfE8w3Hz9yaz0ukuHdGpq/JMzHkFVtMDQE+kdLhUU7tmmdHXmT766otnojw/s/c/T
SAvU9l6k23OBCJvOh5s8d2i4nVxA+KVa3NAfyaNfGULPOJS4lM1GkdbDfHWErh4EsOy2m59GQUHy
bx00dcfPHxOO7+ruLhqjIsuVn2ArUafx8nND6crHjX0asoSnqOp36zGA5J7BHxEJv2o4gWYOOMxu
P8yBnNLuoghZ7/AvGV+DXeWnB6miSBEJkpE42vBCDEkxcGdGyMI8NvWHgnHhQUO6LYrgrkd2WVUc
PTcQoiOzKfeE1+uDBiq/hRRkvzRT1rkcEFiRyH+cNboVM1gXRnWqP6wRFB5w8icoGhTNLPgMwZLF
DP7FlqRdq97g09P1eNEUN9AGYticN5wt0/WwFEq09Kr61T2KQdpfhA3Jcz2wanGIJFn5nyRF9CoZ
7v3m17apVsrz4wcyFyY/a7BtPWA/WzI6iSrURdEGCg8hUkChbSoFz+5d/a9L5aovPchS1SjH6L++
FSHZeJ2nWWfXNlie17gE/15/kA2NyVUJmAk1lKRa+Kwp3IvNZKf8Gc/fCF1M7/FG+qxNOt6YcmKs
+EVOQDItDvYGRdB+JW2uubiEAGxwPw6/YRRc9gXwWTv+3dd/IE3TUTH9t8FBXF5GaCoZdZsDswVI
dSzwF0aRF/oQRIJIW7IC4UHbL9YQgDo6ZzSQ9mXKb/YoQNoZ64RsM2576SM1e9RDHUr4LQtuf+Kt
yo2g30wmyW4kyMAmiAW3xQbNhSOTa2uik3rw31dP9Sk7a8UHSbbR+tsbu1vZgHiaIXx3p8hThIj0
ytooFzABQCkj0+w7s+2FyBt/2FKCEGk2LCsEiaAC+1X4ivgZwMYJZdZTtdfCs1K6jT+iFP0BkbEj
0/OWxqvdRlQSvl7ggzk4y7o2KNCaaCcnQ8N2QyZeY1+2/DkI8BRYcTem8uusCphGLomvPYUkhmmM
HqDqa5h1+zozmPnAAE364w2v0iiGhAGgkGe9g2Tg6bYx7j5t4Hdh2jk1fx701jes17hqtgl0w582
qEaEI32vejZVF64GTrLP2D4xpH3CCV5wi4aFBkLp2e4qmDQJn0u76ONKI3zsCDTKRPhdDiMtOl4n
45BWm5Iv6x6mOXRG9mtAV7hIu7L2mMttn5s90kaP06cHehLJZM9QQj1YGKHIsYJ6sXlYHUjC2Yjx
EYJxAyvvrsH6WYD38zKGoWW5yppLRXdx3O73hvEWuqHEmoNGSUMaMrY8FiXF/zeHf0lQLOmt4DL+
aihH5w/TukPjg7E8YMwENCxMAE6uLwy/oCr/NtzJXYBavBIBdbD4L6AhEZBn8euRn1gGhEjGahik
KSsV5h1ruZUYPRwn7Qw7ZFzyEavAluvyf791fkqVLExsYMZsDBgBHFURrRFZzCyMXIapQGF7Lm6d
OYpj8tIjJnSKDTriurlCialrX1q8F7pPsUQg/2wPeGmjaijyqUyp8D0w9Y4ucp71IPlp5wUa29fw
UINomYVNbaH7ibVRepsHBcfarQpQC7NnoLtQ3GbX4t8He2sfjR3Jd2HhBiAm0PjD9g3fqXPvdptE
biRo9tqv6HB7ft+w/iQp59CI0YVqLFTvXgKS0dIxcsDpZdSAA0M9YzsQpeJZ6EZQtIetcXcznQ1S
x3aa1d9Ayod+HLV7b9JoCoXxTqasgrrEpRHipzNijRfawzg6DDf1SuxJeU0arzgrRIhW9J6n1JaD
RrTALZi7Xzh9+tyb/5p43CAqwCEhN3nb6PLHSy1fLU57g4JjOGEaHZaD+9Deq4A4U5UZ0n4Z+dTA
ItXohH2HWmpyQ9pizqum0pPL1pXLaqrrJVw0jI3UMd+RmMFZ4yvCRV5SYkEHH7dLSbM7jnELBfze
WjuxpGW2RDijlv74p4hVdk73479EVPEpCV27HYaTex6dUh7JOErHHiQLfWwAub9RwT20h7VDSu4w
3UkUt7Ftp/f6Be4Lpt9oWxsyzZpcXDExiRbyYRyaKQeysrLnPXkuh0vUiqMAG5JhA/dyFkHIwM96
y0EB4dH7L7dxFe5zwk62wQPSi3b1to8za6nlmsjCjXEzE8iwyFZYzDZOygv1CzM8uVNpjX6VMFl7
x/eduhi21eQ5D1/51tixiNrATjmGyxi4J8J6O41DZky1PwwrOLz8SDEAfYAqlCwDSEddAoE7tRPC
1FMAf1tP+ORxUz1tqa6lpqhIB4aPfcHuPkNmSFmRiZejbJD5kl9hacZ2lRHiSCLkaQq3IN6E1oJP
YAVMsA+mqa7JlZ13nD4l5Yseu54X0W6PYDC1A8tKMeyV/n4eQt4ixCBVdqjrn0gKWGTt1uk7/zrS
Ekvv6WlEgW9qYzeFCuiAn4zmhmpxw0efLfe28ARuDtWlJuJdbg76fYR38siUfg0ABztvcDRykkMl
EChdR3BfOfnmWegwl3VNhEOIIWOhMIR25Ex/E5s2pI7C7gM5gnWl5Sb77md/Qm9oTXQQvDWvbJ0V
IngKUOnBQCCxqW9CPPuXkAgXFv3IUlrHTPSKWL/PvebxYhrPj8z+7piLGzGVwa/utNESn2oaUdpi
0RYT+elbKmP50vEWVhHDC5x9q3w6ZY0/bb4AqXnb4UwnTr2obXIezTE7y1aahYs6dpsTIuDtD9k3
2ofJeOcPY9XlJkxzuBsfshXKYSjeq7O2JoEcfBqqYgTBSmg1IvmD1yhm//iUY5qqgSAJfiDEm/G6
PFsPXd6odMWSVFOK26Q7fXv+fI+HaFaE00TOkjO/x1EKBxUVlIIok009NlYqss6D/69dqNPrKYTO
Nz69mHxRwnE6HUbxX9gz/8Bq79bZ7UFR3G8wBlO3+LmFZI1Ug7FNoHjSR0DHx5PIw5zWNFH4HagL
c1YZ6DvPnDRoK6XlTz0woDbQL15UTHnTete5+y0ECEjOcCsV2Itik2VyTMCxShaTU+7hCXOgUCCH
pv0QC8FYM44lpkpEmvHpVk2YIkN5NNeg1Kr8DAO35+bhRqTYGo/NdQh+xBAyzgotzMKff7Zw7LcW
zINxbZuuZVvaT3s53VemL51rILM3IDgbFT0/lcNcTlL5+14QILK9euBexmzj8RUmrl7Xu87VQ+4H
jOOFrKkrghoiwF7G8fVjkA/OZukK/+8Kgkz9EZqcJKPugYyup7yJv6ynPTwJ1+k8kCDowWWtzU1v
kRU6lG5T17dKZv4IDGKEy+9s93JeThj+O1gX/TgeKLwdy6P481iArVkpIfFJgo9sKnF9DX3hoVaD
M1k8GEPdUI1/9Tvv4CZzkIRPcd4yEWCOV4J4cVlrsMyQwyvoVEnkWAG/Q26YUW2Pbs8udIxSTEsW
UHPj+7rqx5TIM4yWW0pjINzg/TBxpThDBe+FGioHWNBmBjdUV4thVqjserMdTscYJzi5CSXN9f7F
XjPOGRTyBaGjFkAk6S8Ta3ETjT3vDjMMemBPzoAypNlrGuJID+jYlc9PoVQ2EdudkzjNgJjkmicL
/742HJe+9OFaeXzNzrS6IS/URFCMPrvBcbrvFxyzT8v/3vwtwRnOUacPpyGIuskc8zH9+A2jPd8G
ogCz74CPrKcx16tzonIIMszPO5U5fes5sa9Bbpt9Z0vArhHPjbzm4d7kHPJrcZAXJSYpJy4aQiMA
Q0uC+OrSAF9t59SYkmiW3LPGPeIrGYOdptcBno/1wNab919VPWB0SVq6z97CHUzggbZ4rZ4PGIFD
twWaeNdPhfqGbhYBOOIN2ja0faHCIi+5fn7/RmZFZHUJURwzY7+bhGYneAB+yBkq2yiU5eqH8bSj
1MOmOEd7AxuoQho8amAALQDWFUGURbyR/pMCsF4VLlSpf40xLTPg0XoJCcsiv9VkqZcw/AF5LsxU
KozFn15Dd2NovOpP3Y2Tv5xnkunXK9lUK0g/W2wB4kKb2x5R4mYAC1L80cKHbUGq1ARCrNBU7ZRj
4lxWbBC5gQSicQSWDNAwoQUWbIYmC9G9Dd+NETzcpqNL5lADzYKVe9xV+bbdNomM7yWaA1dNERkx
01Zr+1AG00ay6ta7Yz4bhlowNE7EXmhYz+RqRUUzAvHXGGiWeFRO8cE2SGmH4PK/TrCaYC6v78rA
BZdTOSZM2CNmkyJuqTIRjcl8h8qBUG5ndq0bsvTaK3Q+1z+dVkltf8DgaCRdeoXAPzlxYOEKNom7
2tNS68YzxHbu9wHeNWPl+OkLcyGFuhZUfCIxk7TqW44+IWtiTrA7BXfmo4tjFYcK2/RRBApov8sd
GbGlerZSJkHSYZdHdcV9RQwyzFF0ffVq1QHawCYlvtoCzb6RLnxhPUeXNC3qSwg3MDHxGV9Pn0Sv
+d+UtkKTzJaNaJ4kQlIkXQ3ZoJ8X/VcK48DoGUKn7POa37zCT0XzWlYKp/nAIcbO7JxvqGeDhzMs
L3dNo7yWeTn2VVrOWgBNRnxrmoRBtRG8iRKudYN5MaCw0QZIxjq0K6BWgPdoFryz+JYUMALqwBa2
Brh4i45qBe3TTGOYqL5RMGMK9Q+cZlo5SfmXuJAVk01Av1rXEw1QV0v4fdrK6svVSbgrEjhzYZ+H
LTKOmE6kh6MAMhdFcWKc2BqdOeIJo56bRcPFIJuxTe/T1254N6cKy0vqNq3MwcSn12xePsNZlPxS
1b8hBoYUUod1L5ZoV/7iyO4lBiMKKkRkhC2v/uFAsyJHXLfI/DwRRj9Bj8AusQdpXnb7KF3s8ukJ
Yq1hNDsDTYBly7QIgO7fkndqldBRHc+TyqgElvN3qkb+x9EjeM3zPkGCwOl26ge4JctcdEp3AXrl
QwhLNqMfEMNXRU1QbVl1BdH8zWORUgOU0Bu4zzFdVWfmO0JoS2wea+JXayIoWIgDKqjTEZu6pCQe
JOzS5kVMANngftWqn/eoOF0iDNq4aUdOu76ChuXO/0SLQu6ti9yIRoilTf4IxvZ9jJFoulMBxXAj
i9P/3HHPVmzn6cJKZZ3DeEYr4odPVDJFdRiu6Nu7++suKnPVDT4PWGKylqaAWBSkfBGbK1evUapN
kCdy0h26lP7Lj3Kc/VbXyEo3EYoT9tn2G+/DhpoFz39OcgXmgaO2Zozj/Ykw0qh4a6QGzAD+J9b/
NqzYa/9+4BIZRMdEkO3hoyOG9yycQTUxbHHwsDe6O/oo/Lhq0dB/h4ed0MCTZZX3BMQRprLaVWN8
+d7lXvo68KXLJL27aIpRZcBy3qEaEoIyVJf9WbV+nekR6LKksd8Mv50AMFE33myB/o7yI8nwVzV6
mTRUlqZbLStvYWqcXRoMLCNp6c1S1OnoCX9HJQNmkpDI+GXCsjS/Gvr1rhvIgnh47RLjz8zm0zsf
Fh0KEwlcnaV0BcBr52aAhf5Vwhf/aLdzQ5QRUh7JZOS76aAOI/43pMWflvXNXyhlDtLXyGoYuuHn
OMVdz9bMPdFgKZkeF+PHnfxtiReRvBRANF/M/9IpPvl4u6WAn3vw3ejyiySecDrnv7LCtb8U5TaV
xl6cb8Ke/tfj8qwR0jxMXY1tb9CJc+TLsprYN52uNVtX4KG7j0i5IOYq+iMspR0vN5FaqwbCnLas
vkXFC9nZmzAcuKKZCszusnquerdx7xULtbSAH8R/WRq+4mfubH2bttqim9X/PrOfxmoK0JbEZZva
9GxBDBlRQiEzJPdxSMMWs54IAc26l7b7xpjHhtx0HIy76RMEWXf5VWY9VbN5Fqjig6uS80eLwhS4
61ot4shDtoBSdClZdXsnjVBPLemhGGqC/Obr8nkCP835pvgae+DuZZ93ptD9rDJm0sfJtazzieb/
6CrLhp7LQ4pghr5FJXBq0jOfoEbncimiwxzvfEEHY2xQr62tEZ+FaMBxCwuI7x043Wusqz2S7dVo
wkGOdwCNP0oCqiFJNqpIIN/50YPzd97hYOVPFAV63WKnkonAlRkSOVrhwaxlvTgVFGhe/u+SH9SX
sk5GVs40m4ZMWjcN3XK1BqJO/zVmIqAauD+OrdnFkvhcozdrbdx4/x9Sea5Tg23QIXozrNBpz4bq
gjBxqh16/GLaaAbY+nW9PJZhwdGYFDOjE5GNS7Marp8tdZOkmTsfsR9y3rzko1S2ZKygJ/kvSx0l
amGpzolOBHC6QKEPJwaHy/RgKphw/KypYSHk44EKuulo6OV9n/bKoiaR/o+kZ/iR6V1TFeTAVm8K
2Fp/qbdphXPXQD9S5GSoG+IFgnYVrqSaWo6DE3j+93kCZ3w4xQImFsRU9cKBQECSPH7s7fznrlMP
GaFxafciwzW+kpTp399dVdEUKoFXicRlb1wjn00WnQziHlshMVYnJxYnwTkiB6GEmDSirin8wrxT
U2MuvEJ4YIbt3P8HYOWXepHR7XtcHGVhEK2lrDVq6ElGppH2F4d32E0j65Ll7QxiRObE4wm653MW
HTZX0+0/E71Bo2kMQEXU9sFLCFavQazLodtc1kxEOWbHMZiRuCIc4tyG6gbIGc1UOGxOlkvmEq3C
X//RHdMUZvZEqRZEygmb93ppK/l74vjBATOFJ8sTmx6xTSUPlld3T9l/ddc1FfoblIZe1F98LUH5
NDw0wxDJlEbbE+p0Ja/WLmAt8nwrqf5qAIoN3FYtocKtS4K6Y8iXy2NyGrrvPiIsmLHDBQHMLEg7
LPw2zD3B7MEYuEsxt+oEcQYKNn3o1V/T+GXEnnuI57nQvY2egBagLelxNtCdv9NgILaxgjs7Adjh
Cw3KiHJDTMCgbSlksoPcownIUk/6jLuVS0l16RAnWmDQcMDRtTHju/BAnIYMIjkoUqZ9QV0Vok7T
WmqdpKAbb9PHHNpd5cVXZz1UM2spAiChVwTUMth/Dh9z5PvpgSI0tiO3bt3WlR1bMgr+s84mP5yT
PiOMBqf/xvZGH892ibCoKsJvEOZ7kAf5fCcmdzSXUNH0HgNYh/HEQWj6XOvm48uounu2v1mKavUo
x3eNapz149RWjG2cTdTg1vXXClJ7VBAlY87iFicKbLI7Q+TDoagESU90kdYx1aJtt3et02ceUaIv
PGlH8ktfRdjbfQmxkeIjNGfuF+WlHegBUKdNfgLu3HdE43vmDWg5MMnrYjm6hTEMCKkO+auhk466
ObvsjRCrg6B2gXgAfGL/qKyhkdSseeB3fUGGaLMriKvHRMngzXwfTENgI9piwYtEvFAzjmwjIa14
bGwUcpUmYySwRHWLVaOR2vwwPxsrUsb2MOJ6AOFMYSGBJUWfokEOO9nx6uCubjdk2cH6Mh36wa4v
+pZMzZgF70OfVoSu0396u0YkmohWxKLOgUpj1nCxKgUnaOOhtNckNu9wZ67IWeHIvTx9wmxqHe71
rDlFXtdyYIP/rUG3sHKvUbGIY+IBmhlqmP0rW7WDGLDJJ1v3t15MfVHmNMd38KukZF1GdznOzJs4
EdYjDhhUIgKqiTbHHCi8YURmtYmfa3qx//squUi0kQYAVSR0O6rgxafPbF3PyVR4DHhSeHv8u9MK
VimW8XrizWxcaSO1WBaPdcAjoxheg5Cuud9nCSqzTnU6OuI+JzBi03wc5G67ZXC3P9BzgvlJbkLW
KojiY5soHBtHGaaFNHZq2ZixU+Im+O3BBvZ/ZWpr4XK9ClLaR8nwuRIBXlp4n6rUa95o9lIz/+9P
8yMfYmhCJlS0So0HqU2z+AUMaI0PaGTA52rjosMUwwSTDG8ZSYqYlNy5F3TeKn3ME1BjwTB3UQGv
w/vCv4DDdP+rMmYVP2aFHMiqZ36zc8xagqQhJff09liki1DqD5xZJjb5JsLidFYGW0281ms4Moh1
LwRumDAWOWwCXUHFmv1g3pjmTmyrkLqGCzcqROe2y1PQQeNPydyImM2Fqd+J9J79+xo4M4LCvrYW
vyR1t7voBllCaATbq1xzx5dXX+6Wrlt4+BVh4VnCMwbET7A1AjooiayrTwYJhXSDs7LkljSEnnX7
YnjJdT4ENa3Bc1akj2XexxNZBBhscQvUrLLRLI7P+9kIUlyGDVLNWtQRTMw3FM3qnJKVX8iHnxI4
go0eXcFIzf2rx1fyhx/rTkfmLJUixlxuxBRhrDehHu5b0auUCKRcf+tzBz6LB7L7gpv1A1PYKZAp
fcTn1GsAU7CcetUeih1637UN3FYt+S90NDcqMB9L9yEVs2Z31kqIBTtAMSWEMMwla5AcICLv4Tmr
QaCjC4zBJJYUloIQIth8Oi/XPBcYThZ/YFmeoWigX/iyV2o9pM2qNH5oSO8gHm0Gm0ZdQfk8/oHW
1Y6c8v8RS1J7E/osh1Vv4JjXhWcaM1YY7RYiPmepepia3+XBxsaAts5yQR67M4rGnbJNoHvBp7MW
PFnhGP+ztDFETASK1nFfg+bSUGR0Eez+o9K+QJx1KvfEKsJbHH00EI4Ga5aYGu33+z3EU9B7o8sN
LtS8TAY9DwH+mf7VsWuz2JsN035rN+sf4uEli7SH4p9C2BC948s2YDOeAMK8+hSTjlMjL9b/+Fn8
3eoOSwQ/X2QtreemQFhwBei4F3Kfze1Q3vZtr8edei8vLaORmKzbs4iYLXTnXjoQjjIDQNA+iONY
k33Hz6wix8MaRCKea4I3XKCHWJBRVY4iRcWkdSsSo3Ika+aLrfXTvEmGEXsXxR2OdpBJlhc/1NIz
84Hv6pVpNOQyV8M6OD+1JO+K/z+4ci6nbZL1dBQot12QNGML4rw66/y8LZFMmRlmF+Ry2a7dsizF
U6PUVpp96r3PAzgHCxK0HTI8bqWA4PLLoYgq4irzqJqvtS5xIRdTq4w2r8sCq6wBQk65XEXnJXAu
1zJcVkBF3mAradCZkzkdsbgD1JweJIBI8yr2lJMDcSwSSH1Gd/iK5EiPSD5dv8ElKYQqIEZFop5y
WKEJRmv4hssk9waZBF0y9d9II6eW/zYdzyKiFqb85aWUXbx08+ugslONUhpkIDwCHhQAxB0Ha4zi
fdJ4poSWIJxuGYRjLk1t/gglZ0dTxdct8jGiRSzzvSbJKnmj/ATcAl83xLm4zbJ6t6w9FEdJaeGX
9xEFBwZaHRnzGn9rhSShG4C2xn9X3NxU9Y+n7yXkkLJmYSPq0gyKLWPbWRVm4FBYFNS4qPeNMzn+
CkWjbOAXYJyTBQzK+sMsmVH8E6ztSPOnY/A+Z/pmjVrmWXL5OgjcGY2zweqzruDuKmKeMHfuvwfs
Em6Y5Zdi99aGuhRZvC/+dk7lSTwHmVyc/6j99wTGAw1ERwThszbXnT5iglqcKF7r0kiYdN/frE9/
wa2+JJr6JPkLkwumThN9mFqWnVyxLFVAvqGs6KXzCooOCVNZsEJDs98QyYcEP+H40PfK1+f5yHJu
G20HeN7FR2loap0H0DIM7Qjp66gJKmVzBkDWybXyCVAyYYgXuvRIXwooghx958HNMmCohBfBoRkd
7CPsjmMh3mCcPkCuYaJDp6Nw+WhlXUQ4OuC1006dZym8njxF4nSXrrTNXzYtcMDHkNdv0fbG1aQ5
0k+qYek5WX2tTxMR+JQbCGTD5uov2xIfraxoYxvOx6Ud+eUlh2yR8STcz+UIKpJpR5jJqebzP6dl
ejs1hZEaFfIle+VI1SB0l89jqnmePrJWyROd4cFDJ05MsFpWqfGoSX/51ujPAzdQrlZ1J5hI+v57
YpOw68N0tGo6A5p983fUEUVOhW/qybczTcuF1+6+Asj8TMGNOflWAhpZIWUhLwZX5S4gO2MkxpxE
hmluBfNYFFAJsXsd2sxLf+Nth3vYds5vHRoT+86HKArO0ghUzVF1OqBVyOF45R6o9uTzI/VPV2V/
HZwpMC3FHkNrNMbK275H1MTNmpuomsPKR/aZjAUDvQgaTKwY/vbEr1xMJNVX/GdJIA+/NC3XNWAm
l9z1ZYwN6bzPPuD0/mg6dnoQfQGPHs+XHeLfHQhfuh8VkRC0eHmxXISo/86gp9TyiAAJXhNbM0Da
wyg0ptakJN2xMjzmZ5J5tNxai2jV+lI2i3Eg5mMQFJGA1wEpyfY9MkBX+zqg3NXLUURluPsxhflM
/ka4xr0oLm39/UoDQAa/o89Cy7x1ZCHid25duLkAflskwXxbPcl6kd2nq7Bno+XbUZCCR6Bg5aRb
DZEDCyRg6FAZRjIDzICT9yUD2OcWYXrixd18SzfdR4/F5oHsJNn6mdZxqtgBOT2vTkwPVt/cCCq6
mXW5+DC06lPeOXWJx8QRzXFHfceHX21/2Ar1WoLbAvB/BAQy4jWvlD5nyYDXtdY38ti1D51BWcVe
iD59kPp+LIcovjr4vuFHExh7oGqt6BoCZl3+W02REXvdB/W21ULdeWWsIWOA0ufQFS256ob3HzM8
DhTckc0Xk35TSD+Wn1ni2lbzBVyIOV5dwkQVGUZNaTfXI/HchmWmKVdhBMp6lk3UZ1S81VW0/+hS
etlw5s9AaqDOEQdCfktLkkoKaO0692n1qaL3H8wQBbZWQuC7VcLjMhk4EYCfF+OyAYSae1t8RoPc
3yzFpcab6UW56RsoVPBsFTcG2mgK6jJpbeWWj949XmtqB7IfHTu6YtKNFUyJ98jbuZPg1oqg5k3U
0CU22bbRBhgDv1eMVj3Oek7zWZhb58uGVDytzrGHjgBM1UQMiZ9RLMa7ZLzIspEcbYVcMvPBw3bA
b755OSf+mBwLGXI1SHvRRY5m7lPcTboe//OUc3eluvsTG7OB/t9p8+SMLTFZBhfaPPWP8JbM5o3L
e7B9n4gb7IQ1uo8p8CEA/FnYRITc+5MfYpckaXt4a2RKfS7ccM0wddGpLHi3SCXwESqatx0s+LmF
DY7ubmcB4mJbpHhTZnnjOgDnBx+LRjG/Hkkbvfsfzv3YK9KZVHjWG9yHYlPojv83lOBJb1KykGSG
IAElZzz0lUtT/l7+S7MtIKWqW8xKUGMgFd4NysGqjOHOZfWWMwdcGCNUj7wXwctJGw9jVsPLNiK7
0liYBS34M63+xVlvbOzHPQY41BM/47k8yDsdJrUrCxp9mCQuapajg8G9edp5h+HUA6t2AuA6p27E
roNZyBAm+sa2xt+G1KDpsZ3FaFkJbvShYrRJxrvGu+qlodJYZWsW+SwPME3w3+RNs9ey6dprmXuB
5x5ZQMMtNedXDaOdFiJZiq3xTlnHtBfI/HyszUCRumfHoR3PmjJ7KClxSq/SqbzLeEhK2MU16NaC
Mq9bPf9F/6MSN1lll7ffNCi57l2GpqLK5TMcggx+WIYej7rds9Ovn6bsovT7GE0kjW9OtmgkJXOe
U3g5iYKKVsCOpt+9Hpksw5wEvpHruWxywJuwj+ipicOtAgvesSuNcbaKxsAkFv0FBR7LEhZhwPz4
Dg/0KtLCvskHuhAnZFRETFyNE7rH0YHytpEpUrZYSUY3+nXJ9L6GZHvuvT+t1lfwCjFr9RoXoXdn
A1PEa2ythCKgxUCIGic/WGaOGN4bwycR3Sw7jGmdvKaPLOd8iCaUJSyFC2QRb5oPTdlpnm6J3neO
p/K75LIvW79tW9mjxeNhP874RVsyovd6/5QHBX5q3Y1ptBzHGPu8EgPPNY84nQ4WD5l/NFteOmJr
nNgI6a7XsJyjo5uK0znN31+nav3DuHeqIFHwORpC3UjfZVfh8YuvtTWowhWxyr3rKG2pb2l0T2fi
FN4QkiLMA9vHNS4tUeBrrpIgSxZUAz8BCfneOj+Urisuf5wpZK8ccGG8v1yKbt457O46KPaxo/ki
gogDFiW+ZXLM78htWu1qN2JKXkPkzMcHq2yUNugo4OCWvrQh5mvX5fKD2WcyIijXo4daEZqz7nkV
CH33lpYrixQMD/wnv0a4z0NS8eFxKalzLGcISUuSZtQEq4O0xno02g9k3ef/oMRNOupk8efTZwAl
p7r3XWCgC/Q5i5ZpUzSDJ/+MAKDbKMFpYT3QwBsoIedTnTVrXK4dszzIyOT7zEm/FeVEn76lVizB
WbBO3cNVowizNsjcrSeGm2QLWt7EPyvK9q/ndukME5XADWa9BREiOVymAOucAPyITgh5lG1O5cu1
uVJJ8bvKYM6jBzM97Z5SqdDLhNc+7Ipag+kkMJQKfvFxgv9+s5Y+TJLfHqccBqomAVQ7OCS3RTOQ
JRGrtjXgBKscCrH2XepDLGwzPwalx/sg9hlH+0zNl4ZRGBFo7YHv9VJQzWEUqu1cusGCTU1rx0vT
qPgj8FtY1fNvoglMCn5gBnbI0htEhQAFxlvLAd1L5vi74jt8w7jVpbkAbpf+DKEl6EUlL/hwOAR/
i6VhCanxGLflSxVwX/Pk4Qbx34mFmHYk1CSnD/ipOL/83KbVgROih14T3u2DMax82IBrIr3M0XRH
Q+xQVWm6tqeHVJt1JjMMNLTmUInUTNUWPXsY08Y83lCvkF/PfHPhqYYa6HukCq5nIUHfbW5vBZ/N
8NASLJxeqMKULDBk7ncQnB8ij1Z6I9RhNZ//Nuy+N1WvtyN5zUp0y2Hr4Fe3dDnXCZyU0LebNkxP
kpLC0G//3IJPdXYPrhQ20A8gZnrnuHB705+EmkIKmErY98aEeSqn+IiUsOXztlbX0mI9LjVf5CsP
vABaMH21BCd2Q0QT0mR56SI/y2tePochd+QB77byFtS3ALz1pUXPMXRaLQlnM/lBkCPH7DcAi+5j
CPuMikXzrmvMAObfazeB/+r6u4xDuLW4Rgc8E6eqANC1oJGn2T+x/eGCwCb3Au9xsHDDFnoc/Tks
IM5faQWbts43+La3Yj71Kdqws2SqUUSawZcFY1u2kZIRXqHGBl7ZBoIKUt9AymNdFBRaufOxj3b5
809Ebfb3YfoIetzBorV9o6bM5UPPfYgJfYbYUSa0F7oWWnqrnaw0HDwf6ZOYBqGbGdm9dPNpaZKn
YZ8KheSrNRsYHLdNCQekCjgzA73NtsT0s5O13nkDb7vhmtCBXLbT/DJDZOIVCN1a2ClLVUBc4bLK
NCJqjBbghK3v6cirlS8kw5OLe8F8O3yc9zRhIN/5cX1c5ZLEsV6FqMwEu7/RzNao7jXm9BinpG/w
IFrQB8Taxf42//lv1YRtVaiUcsBO2A6J0JZRrZ93nacDCnFLwgqI+wWA2n1LfYqsWBXQpoiBSQm3
WhcJhISzsSRjPnmnT5dGIVreRr+svwRGQgAzP8T888GNmibZFH/zwbmakz7l8u3MwAQkl/R3Ihjq
M19fkgNRxSVak7A7coKZI2+wnlZSyTJSS+xpVhKM+Hmnxt8hq/IhtTaMDv1K2rKVZQVBuJW/2UvX
soC8XXoNDv4YIPqGUp2IyfPXlZT2ZLmqRJat4dVgtVmtWbSBD15Cqv2vhfmBU2go3H8yEy5EI4s5
Z5kn1bf0B7CDCGxVO4qHfB4Ylqh2omhE6YJJV/Hp2OuUwV2iMpQaQOQ+le7b/nzEJPxZsnXhgmw8
VMjNgARTXmV1do6l7Z+CnzS/80MaqrB0WaVvKRTBHjXtXmHKE2jJM+vHMz/vVzMgqTlHH6nh9Uza
MMrZ7wcmPkxJE0INH/fROMXpXhoQ8Zcs0wdAdGqoxdguPnRGiy2NXcVQ07N7tnfApo6iT17hyPCO
IG/IIXcGT/KqquJEOQjDYD4jb46n7r85yrwBoNUjgemAQ5dOozBmZXupAWrOGJJn3rQ56uk7dRTh
ZYjRmz4g1o4g+10tDalrOs6UljcnW1x7sQjwVZjqLMlTCKgZkvCPk1xmwUHTfqzZQ6BLhLguqYNy
CIzBtSlh5MDJWpfqkZIQZlsbso18cS6dDNm0MXlCb7asTGbXqE9Wqs7Vvw5rq8N5+eNcZtjZHbV/
Pu6QxdtUtniQb6I4scIeahbB3/sTtXKK4Et/rv/x1DjnaZP3Md7hDrzT2GEeAFfnMO0EqfdCzdsa
Oxesjjo45I1VmCeREjRJRil4XvY9uqRRASibR8cPgeQM5wHes/Mr6KHpexviWQDgEc2klsMXsqB9
kkziJyQFBafcmcHPlVl6sdB8Qo10HEZkiJ5huPMGn/3GxNMbw6AiEkYV4/1Fd8MeJ4WFbbbYCaVA
AvsbOWS6pa6vXbWvDxP1AsbY6wcpcu21zdy6nB3kx9AysOIFEof9Xxd49RL5C8H2f9660XndFGeY
2UvuIVg8Jx7aIzi2S+og4HsyQdoDaKxJzx+eU2Ch/ehn9JdzIH8Je1Fn1qkFdLeRJwk4bei39qSL
YPHLEAyuQ6A7UBzulqJLiynYYumuOAXPyNJYzF0xpolXrKiB6yiioZLb6x8RiJv88sQAZcO1hJkv
6BO4tkKZ+QGJnAXdpL6EFamtutGFwITgyAMtBi95jsDe9WDWY06GIg0sklnJ4vWsTdEs7TDdS1fO
V2J6xnk7Dg9oico9mpeLudAktqDUziCSeGY05OqElmpb+Hw9DvBMNWWv8K8Oc+YpOo5CElw6MNWm
6P0cZJLUoow/N7/SDjzpB04gQ0IzHAtuqLVja0DMagRAv+Edz2QZuNB4iofzVck9LY1fUoHY59Pt
XzZ9IOgNzdBXpkNfAcFlpGmtGJJSbeb89hg5dJBtNcyOH4Of/1UhKeWFoDvRt6ADxSIaN5qrUfuD
IX5c19X1y7d2//DrDmn6MdWrYV8esDG78+OCqxqQOQ0fybqG4XNORzRB3gUme4cMbxAGEq5ERqVr
D8ivaaBaGk0gqRb9P4JulZLZ0QCbU+c7bwZ5VMVu0GPxLSi7rDRexTag6oRjkYCRta1OAxJv8jui
HjTME3WBM9bzC1A4xuDokiUP2P3LTla/E/7U5/IcMVqhixYpaclBvwODvq7jS3xzV2LVYPfew34L
339/nmapSWmaRqB0A+AAoU98b/ubrUoRnNFSWBYLPNLkXl4yhPjnixpShxQRKfAHlqTig48ckVyv
sTZkgsVJC8SZQwJJsOhJHMGFIepIFGEz/EJ/n2jBjkdsxSlG8TI1wAI5kdjfh+dlmikE2hjwIbDZ
tZld4tpZJ6CXyytOGbtZ2jBeYv1JPI2mLt70Whg7LBkWNHCpzMlg3oQUZYb3Hly8uLfGi1GM/kE0
+reC5hQS/BNgUgDtR5m/G7GF3wk7JO0OuDeVKyuda7qhEu37OT39ZBBLRgSCSNHNYJZOIJJh2OmK
U+/r/51/+FFaLEYOmZ1iq3SJaATUNgSOIzcBjGLuoPmn7il0/TAA6zHRY7xokJNd5AIqmBPJm7Ip
KsYgck/L18L0i4tfg3JujO16r7GDm98stB2BJH63NUeToEbB7boK+gK0KsDXPCVSOFCdIZLJg/lo
IviXhQ80UFSs9dPI/eeLQpeqC+LjNOg6ifDzzW64G5Kd62AUlOcW5gzBLenCf2QtOnB+Sz5X2cua
HQn7v/SAhBEFAf2TLaaMxNsoCjbrN+UTPWaNuPrldRPJ6bM8v9tFxdUdp/F6A6wMegg8J59mk+yg
dvu4IKr6uy7N+a65x4Uv7XZXqdMXsAxP4weniR7k4xOmqRllcOI8t1ykxohfWH7Yb7Dlpzwfpagt
T4Zu9EEIOX7e4xKC7JrGm2HpU0dCLZ4fF437JM4Fq4lVf62ilAHx2EGO225ZsD0I6stBUoNLDnEB
HBUK/vLG/uz2gATlv7tEIn8sGd8h+WSagbx6YGejmGIEW85OIjK6J/klb+O2DMgBS8kIyY2lEglM
l8Zt0dY2svV5qOUX+aIv17WBWysnpdx8AQ3AQIVkRxEB2IAlJoIFEBXOhENiSAWLE0wOusK/gN6O
tpzu2Sspq5A3QbRUMgPZqvTEyL+mInfyIDd1UQwavzHjZ9b0Fof2xzWUjMhduPLvA4VBVomiDjTg
It7dqGADJKclX8kqKnZCydoJ1pcUq3eib8PBTFwIP3dnsWfI5esZ2+ZMOjfnzLbvioxHzivng0TH
UdeppaVOdVasjtahH65CPEoIMgBBehMaLY6tkXHmmU7X+nnS+CwolnYUTMLyiMJMGChOIbadN0Ty
aey/YxmlV9PNeRfPmBcsmemhlRt8xZi2hznL714VecRlhG78BTTCuZJDR8WmmB/5BC0Hp/ZGevzy
2xNIadEtAO+Q/3lx1Kty4zHawUIrm6zKbVZTBmNw/PXRF/GYrKCKPIiFPWWwSyktd6Pkd3H+6l9k
BHMUUeFGGhtSusSQE7CqZKuQ6Z00L8hps8BtzB5f5oJRBOCTVkJK8wKB6vyJ8z/npFgamoKdSpm6
6aUNdCWAEZcJXHA/A1BmSQjTFnpVMZbkB21bHQ+2rSiPXQmkS4aB7hg25p0tQ/jqqLOkeSlf08EP
th7zUhlx8F3rZjhmf2OBeCsD5dx8iGoaaSqt4fr5THS0tn8GItxGp+fqI1KzUCkqYM6qJmrohyAw
RxJejuthM3xZhuOpwB2KS50VgA6GnS0rSxXAJGE6s4iglINlKKso8Qcjn1tLmgYay+ruatLmSiwI
lCvd0MMtEjJIvnA9krCkTw+m0oXFUaU8dXDQjrKCdCmCDsS0SYHL+MYJFNzFzzMOqKmixnnFfQ+v
CK+BB0EQRJWApqYn7a97RCq9id05aNKIl29Pt4m4IHnpT9oNn7Zo345wd1f7HYaLFTmZ/jcHMPuJ
qjQCOJm9ipyfleJ5XJrXrOyPfGxbKBaOR5NALkRa/OLAamFNP6Yvb4zD6lfeA7klJso2CVSAo5DQ
+9wYATsn4ET4uPlkXyRvQ8ozsg1MafmU2NOI4h3W2+PNrwzoQteCfXbkvDVeJrQ1n6s53q+d0YGl
PhMRXJxju/ICqZfHZnQd8zrblLz5k8vhg+e5FDejzbJl3yJXocYXinYqROX9d3b2Cc5f5uctUwBT
SL306zS291kAXp12AaFiqOSclLKIt3gFdVMyhEAFDqchxLSoemx1TV/RteptsuB9kP0oIOR26WAR
3Li1j2w/1afCz4kdgclAij6t9bLWAzMmOKU789sayzvpz6WTpaeSqub/5BwNuxAfsdKt8cB6xq4B
qdo83ksLVA1Wf7UJDyC66wFPYwBmC3x88b99bTOo5V8YvTG7ge1y8snzOJIAkhKLehw1/1/n1NMo
XjAbM3OetpyQzGcH67R/5tcy76mQQ/qRvPVrtsJj1V50QAxZ+uQHAoYnAVXQb6aqrPDeCFNE8mBg
NUYJccgs9g+lHMoxhu2dt82Gix1gxP4OPsYKsPw+GFqXKkw4eCv/8PZ4ttF1oiyA+QdWxyGvw9W3
bN5yVcsW30LH11kA2cpD2+9RqTb1FEYwBH/oJGdDj7qenPY5fkFsHRZVlt9wL/bHtNw9GhnCRR90
gcBC1fdKrspTLIaqUVlNHuuS7LQF1abF152ByPFadmade02Gk21ZFK5S6RQjkU4OFjPCZHIfJoCh
Ydpz1t3GZ/u9M2uhE+yhKb1no7vQIS8FBaQHbeqhT9Lsac0UZKzPWq3sVOyGx2+0Y1HPVB2P8Vi0
KXvH6PmmYrZi8DzwcLtGcyNqgKS1w9g8DyckULICk2NtBsOtYBQpqcx42YgvML96YZcpE45TC7iF
Vl6QtXjo28WM6k5mhcbrfECHVoYC7nkwz6gnsrlde/cgcuq4tJaoXHLjdUKeSg8wCDi9uNLns5Li
/muGoCrw/Nl3x282KGQuxnhR69Eg+yUj+sbllG8NVzG8rmiwmb3sQsdzYBF1klMB0A2jCajDNPHg
EamdEp/bpPhBKiEts6iqsLBwS3WF54c8wrcmp+mzIkRYnMIK3w9gfr1ECIHvkRyhqJWJx5Z7QHTj
hXxTm9rHCazbiUs75X0JzFokd4MCV6rQl0gq2dU/+jnu6e2hRVWW3+AeEm0eHvjnOHuwPvR/sEZH
7+75hV21cXSyHYCSG90mo1NiuMONgIRq5gu6wP16noVnT/DlxNA+2n8hnCthQjVSvQ058ZXrYTa4
jMo2+x+6vDrFSz98fribMfGO4PXliEntKcGpkHCjOnBc2beH/lAB68HZK3XE7d7hYcNQweNaPLMa
20/6z6oqNuSfMVva4Ev37WfPDQCtLoidJPwWS9h8r3NHAcuKscApppuG4iYfRyUDocTIOoBxV3ZW
ft8LAeG8h523U2PryE0vQ+vCmBfjpEWRlWblERdjdkLqAuMlsGdUN8os9peMSEU2ADOo3T39lAuS
6Da9lpbAYCv4ruo4HjsWqFkSl7YyKvyaSEi5g0G3d0ODNmzis1ODsVud2sfLJOxpF26wkyce+rSr
7lKzvabC6jZmzmleHf6nQ3qzyEPjLsHX7MZazxu38TdrzSSSjGzGyV6otDszpDI0RCgkhZ8MIF5h
1fZQ+/LkosW2+pysZQZNOv8gqD2YyWLiwlCQMkIeJs4EgiBA7qOYYXxCU+GLqFoHDNbZS6ZahWi+
6IgHcuG/UAgPA43kjrPMsydmy5XeA79uyDGq3js2AjDnJGIaFkqRkTEM2dhVaFnAAIpKt4SCv4RJ
0WHrFtDh6eM/cC5FtrPI2i3SmG52s+0Os9CdcN53VHhBH4MtByw2L5EeALL/+AZDZFH/sHe0/gZt
wZaQIAaOWiyXGGval+sUq0yg6CEMYdvzC+W7FQuz7xB1K7S01vybI59ncFk/hX/PZYXWorbxkN2O
Y5hXfoHWlpwwWR9cd/ZRGzr8f2CG9b2iab/iM6UZ0HpKbL7dDxRlXEPGdtJhTOAGOlaQqW8P6NSe
Oh2g8SIwVJv6AwSIP/Je6XJ7s1jD+nwwGolPidVMqypdRIuZRBraH2TDnD/BVsMys4piDQvoTeOq
c9JU3ZwqY6nxrvarT/df0u+uOT1R8NinsoakJ+TEpFTUMddeikMRnnNHsSbezSCfFYwut2rWKoax
L1Uc7D2ChZ66sA4cb305RjtO2k33TRg974BccAXvvW8mhJuJqTKw7GRiJjgY2FnRwYFfAf6nsECJ
tPKoFk1kgROA/1Lbo1+i+YFNTd4bVon6T9sO6vSP8OXsr/mmL0k5jEqadvcJMXsctJvNvyARm6lk
VhuXfuBoQv+VJI8tklHjDBa2LkOLUnu7i9epiPiG52jEUudU2enHEhWqio1LNQgtOklqJdKlKr++
F8HaRoOU8PIdePqCwZSLJgqMu+aZ/Q9WRjNpp4Njyc5BnpB0OkX0DX6wEYfC1INLmueknJ+hd1Xk
/cSv+OC3GcqRUUl7FwOY2Q+vlOgtAOmuUmwpmeNSmSb0g2yy4YPqXQTN4mSkW6nY5J0oX12rKedh
MyODm+qmKkrdF3Lh55yMqfXmEZ3hYC4VOE45OBNw/qKq8fnxcVFo026gzXj9Ud8jJMqFINRK3tcp
WOPpgbdP6C93f0B5yWbC/0GUbUfRfD7XAkzax8I298/cHNqWXOYTknBqRse/62Vyi8Hl9xd+DSVE
4gZfP+W5Kj4nGvy8rYTuGq2fczUEtOv78cOt0XcSpIdPH/f+1uxmACf8fCw1qRu71cMHG0PYmKRg
SRol1Vua5IYQV9jU0RNj3KU+JGmOZ0gV00yG2y8sTRAgH7yMiV2VnTt0KxBgOEXQ5snHAV+qiLSq
3F9+y12Jn+5agOc2KwdxGZKQFfvGWymRPMfTiQRKMKJIVj+Ty0v3uxdkgjZh1VMjVALSe+URmF+X
e9tOypk0MHtwcLtichtFz9xmDLmHBtmHMLLsjhlgQSwWaVD1Hx/v7Av7XhJ/jAeYh6cFb6NHrq1T
rmEw+h678/p9eaBq7rPA8bU10yLT5m3jmnIohD+gqlF6/tnRAzld+ZIKGQRvU6FjiieiGbfYpu0S
ArUZKVNVmq2hANbu5xrVStjz2WW0ye6klrf7JaC7MimJL+E9KfQd7NM5h5Rk3FZJSr0ppAPKXN8K
4YQoQvd4eCn3nBZAEy0NBhU+ZNzTT2fOxRC+Mi+rBrOp/iOx4zI8L61YDqslAqRKYQqAg1KVcdQr
ZpIiPc5PbyCzRMX+QSh+eV4vVA25gvL3AT3dAjXfmGRlMedrn5OBIR4PbP91S2ZOBRdTuY07MX4C
ZCrcRVSicLENZ+Po7+dvLT6oB9e4gkwGWwYGE4s/STf8WgeIP8xnp5oXBNk+FrgcqFsgGls+/cLk
uiQo9qbCVx6U6YJ3rFWcVLTUzm6as+XTbVckHYOREawFBNDC2qntaCO3S3BJZpzANg+icgx8bmxh
mDpUoZFFFt6mYB/8O+uq2qrHlKnlRHKa9MDFa88JJMTnGezvecRvMMMrm4obHCOAFuPQ00WLoTwz
20PBVYBWm5MiBYsyjUDYbW5nymHTgjryERnrURdP4wfjek6k8VZQC+4rnw/QgbXDQmasa52x4qsK
jOHNdC8m2aDy8U+apQPHOG8YCccSKcs9eMJAMuef1vNsY815uuN6NdODuEOp5GoSq/3vOVSDINvT
5snEqAiinT8Tkmu5j+kSPO1zq7yVFVDz3HiKPnDnfdaRlzb4PXv+X0GUNF1aYvDg8tsy0qiHn+kX
lk+4SvPNGME1Mt9WampD4uyMXNBD0WlCf71iMbQ893B0BQgJdjN9OL2Fs6A0Snq08nMqCZH27TWV
xLOowSbd8QI2Iyy+NDZsImIp4toF5Q7qvCt79E1VqQNEkbDUSlEYg8MNYwWghEBLIYzDpkNlW09n
ZvdlCmb9WVGk9R84HB2R+YhZHegTFLvTABgKY4DXpAJxmXVkWTcsElalDP24aueCIIXhvIGQGvPX
IHe4SpdYBFQ1pduHuyctVPMB3henw90Eh4mgE5lggkbVDVDfMRTJw0ldesz/79Q+yoC5MLX8Mde5
hA00949HE8h7R6JVSiZBJz+SQbUYVxbKi89IPg+O53av2ORlcP6kD5Vjqgr3gVmdLMXeMCXgf0K5
MPnFbnyyKjkTYmQvDwykNk1yVnjgtSx28etJyYVIGSbDDURcn4GkopYxbhm1xDAcetIEGaYvXc8n
ibaIbExxKlOo5qV/A4y2oqv0BVUDky0esG17wzsMp5RpETej3mgw8NbxL5VU/hB7LYx+4JFAn3fQ
cfthPKCXsVS04TnbL02bPS1NuIiPgvscMSp0PR0MOj1dvAfpTB86GDGYKvat/PnNw1vwtDA+Utju
EioYaMp3vuhKLpuVEPfw7RLZrroxW/+JfFOdrgIkk2CQbURhAgyqt4ju47pk25Thg2nmRq61mFMW
gLA/qu4bQ33o7cqu3SK4UeVwx2vAvLKCz/QZhXadUCaxmK8zNGFKoVdsl4SCneYz9yAXSl1xb7PZ
Mi5PlEzV7N5KnJz78eEiezHIbq5mXGDamLPVjFuh5IphwJBcLgwFWiDgCKI8Hre/Yi2LrmLxB/xM
kNRJMd0l5YXAvle/DaAF7hZUz1iP/9ar2mA3AIHQDFd6Pwf6nQKOPaIRTEI8NCpdDSFr47jfPHC6
VgLegUxiAgee2S7Wxbng9DFkrkT++a1QKFrwbCnhyXYVGqhEsKQ0gWmUiDrxbHBAFTUDJ4QBJUyp
zKslmzEJxFyyheFqJWwPC+3ICknsHFo3qwPzX3mYrWswUpsptRyiIX7PGwICfyhuAoAPO8xDZVgq
cDE3ZVKmBEHjhXS7b2ONYnWs3xGNTevOvebQZs8bNjYROR6bIuigLekHNbp8i6WEJcJApsujXoKN
3Yot8736iIIwwM5qOO2Ce0FCMTmBLDFWUcYwjJQVONZhgWzYyL5TOdWI/2ikY1K1f5kpu7pzYhKu
lpeZ7wxrUk15YWoCk8BoTM8OpQKvXl6grD2csN96nm9xl1dGx/tbr3i12Qzhps74ODSuFGtUENEk
BMyPIhMQ39/F0wkxoy9d84K5MqG3T38pAH/YEqfGZYFHRsB1bdHJRZpOuzVaFJGOp3K7oVd9Ajtj
m6q6X/4NbJPd45zotlbvSIKcrN/eFP82b45ze0xgPwotVz1pzcZDkf6xTUw9dU35Z95KuES34Nc5
hTOjaOJpAyUPDf9IEcHISW52+OsEPMq7gGVCoUU39bSAagB/g5fuScp5MnxaZRDEUwR+d5060ZB5
281xvJjSoa1gLZ22isrNdMnACxz43NAzR00QVZ+HcB0a1LAXsHcUsRC1L15trwLak/36oPaoTCDi
dbC/Pxx1YpL2+eljum68Z6731z4tRgs4CiHum+SEvY2Otc3+1O7w9kCSy4YTtAS5+I4fXmFBCxAD
NpAC16jaJVidi9IxrgJbDjazwfshfa7zaT/IBN1J6yhLvbELWPq6A2pw1liKhNpCJYtf5YHvhsKz
AUNIL8jiO/6f6dxhiMLSar1GfXdoX9PTnggqOgCjSVVZ0mUOhTScCmKVpUREXd0Cj4ctLNzW5AQF
RRsF+z8uNyFeKJrfMLoj1bZZ7aqvjPcWNe34fYNa71usE7ItWKFIhMO/wKYcIhZkSLX4UT7CBI/M
SaYOYUtDwnblIrrg3COOnNN/vAknOGR2dTGAgCbUb3hjkn4SesIpyDHbKXkrSyP5/dj9zOpbdjE9
Ps11gPIgnVD8kejN9k+CRq6jU/uEkGQurOJgSW4TrYokrECkA/KPMmrlaGpyMVRXT71Zz4W7Oruu
ZVRY6cp5Ud9lGKTzVFDL9zSgvpppBLkos2UCzZ66W4bZFTUcp5FflMSirA2eZ1LVx+gndX7NS6ph
a0ZYK35/7fnZr9JwcXhhAEYgAYQpoqaIw/ezEf0c4OA5fLQVWx2Ee9NwYbAdrz7fYZK88u34R0Hz
XlOtFek/oO9uiYAt0LYYV2U3iaccD20GNTdWKtSuHhiIwp4yb6PLk3ZD87KLdyj2KJ+3i3e4k/we
nZh0fS709QcIS7xqKOZ/6qZAK02YXlM6FeZsp13nXR8XPCHJkCEW9TbCCFa0CJ77znUfDpNcCZGr
NJBtkgw78dn65TcQJ84jPDgNJlAXmv7qrKhWtvFj6EW0uEzrT1/kdat8V7lqM6AAo2ecZBqvKK2H
VEWU82h6MdsxTPnOJkACpxd9YNZNJtWbuZz8GtIBOMub9Pu0ZehS6hyVrtr7xl7paC9twVuXiWEY
8E6yS4wlUW1uR6bUowEhuSh3JeZMP7yO8shWALrbkGsuX/cn6v5nliwfFPWV/DXYNj5WiI+5ajLX
1X679dDPc+KT/46UeEWifWdeR0E2CWD4X40oTMJiv7eAzbCjY7Z4jcUavEndD57FNp9Uso2DhRVN
Uon+ytOnZxWTQilgNY826qYUea0j+qWnjYCCSUZGPqUqyFMTTZ7PAxTh6n9f5mUiPKgXLkQLwQiA
apb5j9UA2eu3vxjVjS40RLysUVBxSB5TrkpmAwd5Dk2hVJUuWSMRPKML5DtXrfq6DmJFlwyzZNWo
lqWqogJFKloFFLObUfAVnfY0waQkZfs3QKBA7kAUYVqYpPB9f2FEBf9VTyhSopz9AiohWfyNnnih
p9OfvXvooDgL+YFdg04yBsLbKg9zFScf6Ez+ZSf4YqQWNBmRv4kkt2GJVjS03PtGtBsTOJ/+mj/n
IybdMmZ+8WEtDLvRpqnOP055yHrO5SRAH/4w44SLcIdPdUtSSNg1bmp9K0N96yBJbJ7xcdol+aOv
7OoWGGfibBNn28WMeuew2X/C9iIBzzi9hGJSf9kx8bV61MiaxCslKmNt//qbyAH293THHxP0Pgsx
307PdjOdT9nQRwJwXy/0RvkAdmibE0jwlmDQJnZRBBdv2IQpLbCUHesD/IewB0pGyV1O1JJTzsjz
tYQ302hjmxCVxiP7Q5s9RE1x/oh5UqoQCCjGtBvQ37k3Ug/T+kqX/y1KifpNj0qU8z51QM2tj65F
kgQj4ifVkHUppJZYh97Gt7ygL/v+emP82ombt/gPBv8Q7DZ4CEzum3jowG+HasEaAxecyx5H36B1
m0RBuxMPsZIU1WhD/8OPsPQlJrgJLAIUQo4xf8Ir+1jVrzveb9JpnSplWoK//ga2Baxqk7GnGIr7
wGPANlUJppeoSKY5R2WYKWaMpeNJ/2djkaHKFIUAXnhYUCSMxa1U0gj5ZRFbzSKq/s3N+rFvXpnr
hkrJpmL4LRwYbGAWEKrc+Wzvy79jraXdSNDkUjTnYft+rBlz00s4oV/nWk54xtyvwrn1VwTcMfyO
QZ3Ym36iyK8O3o8U2biiXMfx7ZB8rvQaeLwMudqVxZTLQk/l/smL21OVhSUJImydOOpEq7DZRhXw
FtmUpbgJtkFIbQ1wUCRz8cBNQDMgK5zWcT0dfEIl/InHL3MfZcopPad7/+NZJ8pFptgGRFrTubuG
jNlfjFju7Jn+7lzR5nupLnx1YwJ2vU1KTVDbuk9bFCw+3fFbCVaY1DhHibLyxK4a8zIViNO45Znt
iiQVaMPbJSipeZCwdFNvh0baIE8u9CmgIC7WpPWQA4Aykdw9MS/d3RQ6Zj44qG5MN/saE0tsD2RR
oZhSOXdIxCxKZinNe7buatQonRveGg8Z6+PJQOJmZ6klOHOQ7+rEa9u0Bcpuy5Z79CCPX0VvYlof
oLGZxSm0mvQ1gWlW3RC3o7cTDZS8sG4hCojNWfX37vTlV1JE32dbtXclG/H6iMeDZ5FXZSPcM1Cv
+MwLl1MMBn896/hciQqxRWtozCLVheSjaIxQawXuiQb1GOCvEG6X8ZVC3ho5eH6aF/nVmXPatuQ6
1xwHJZB5FKdVgGgf+dgmC942KR9KFBkuHaeZbbG4sis93R+5jKBxd9B7ZpcqNiDjxwcIdJw2JG8p
KtR5F/5pJaV2xdjx+BS7x/4Co1m04TIM/VrvYyCLp1oAsvqkAvT0kZvTRQ4ocDdxtSTIa53bBwwr
WlW2ldTRE/VqFycV/7K3FgpmGojTEwrxZ62PsSfkq4C6dgsbLA72X1k98UwyUra/baGlPJViqFQs
5sYze+bXYhlRAK4aHVh53hzpGgpF3DMtGxopGPpjOjDETVb5VeHthsd66mkJlGpGEAyks+65Izsm
cdZChONTfInKHJPIPFnhbiQX0yb7ibz8xoXCLXIG7UD7Q1QZSsHxAkJ+wkMwvnQBklxsw1EPFRXD
kasuRZpzo4brKKg25QFPMwdLuknx9DUvvB0JH90l7Iez93TIfR4GNKaJlD4C0bFB6xGZRMZGXxTZ
g7H+hNF/BZt2HGlfAxpbR2WCB0eUIrjQl1MDGsyNUXN/7vMoghNzac5OM5mv7XUZ1dpuZkwziJn5
ZSIEtb+YI881iFON+9RYH9BNYm7yi63UFUfzMO32ntKTbPLV+jaM6FuOamv5e5V0K9bdPMmtFblq
h73mUte8ndrjz1tdkKyhCa4ELEdC5NjwcYnp/cDGsZZFaPOwtQbtMyAEgYgPNcXfZ60qQpYUBkIT
i2PklXu1i407FgqQQQav8/YCZEJyrKV26IVUBFJE2pmlNWLlkltNvS3B/pE9yBbqHPs2GuJKA/Nj
ixNPFSmpqTeSHp5nP1pgda6J+Ejhgh8LD07kp1bxRBU5Mpt5jiIZHMgWVmz9n7NnhBId/qqi0D7g
zLuDqDffHuOFEsyLnDLg6AtmO98jnehwFv1B2JRs/rTxEib8YwD7IBhkGq5sIugjcRsZH7XHzm34
sasWXeQu81s+Sw0JbmEGFD8yXydjUEPYsrqhXu2c4ZLGSL4O2b5gXI534v3qwXe5rhVc1Z6Uc3L0
kP+iDmGduoQYbioiyDHWfgJUiQGkRcLp77vzKtAhverKofz/hJbol/37w4gX2d6UfmdgZUFW/YUg
7rJWoqTu5lr+pY5AlPLAN/azHdq3JcU+q/ef2PWm6L1Bnt/ajtUYUpSkEclT/jINMOrTBM96AgAN
xkHHh1Ogwdi41aM8lx55E8H0cQXqS6MRyF6gARXvP8NSicSrolwA+ukhbkTAQ6LvucFdrUJbKkKo
ga6DlacMckrzUwtT3EIuIdFTsNUQyRpF6dDq0N+I2RTrR0uM8k3mVCB7iDdnqtHn70uRVM64wE+N
QCroZrNZCXQF6kGPiWjMaX8Gs4S/MBxbFxG5896lnApf4cQm3aP+wmyo3WnWQD+0+RaimimJWxMq
cMgVyNevRAl02VElfZ8eYbQeeMKKPgcRZQcVvWQQMDy8OdHxG0MyNpUfi2NUgYCYZIT+bfLt/oyI
Harq9ig+QRLvn2vlbmmwXpw+vLE64aFKq8J8EoLePwRTRRQmB0M/Zcei8um+8DI+ZDTUKvFXXtu5
EvFcSbLqUjHMjhRAevvnr31vxuCjRakZm+ZDecOzlBLcavdhzaV3vyFt2NDQaZrgamuLAE1Vrl+E
LsKNumcHYUmx1l7uyEOK58Wg5gpJfMuJL6R+Gfjpij1WYPpCG+i7KG8UY5EtR7qMcBslyiyAEXvI
RsO6fSiwhqMjniVlSc1G1Oy/7GlVsaO1nXGYBnuHX7l76vFSZpLazb3v1fW3EomQq/eAxevRgUn9
ENtRrDHGAoawZASQ4Tf/vkKJQ9JWXZyvA+cmkd41jLvOfU9kTXvw0tW9hM1VSE9pF1fNP9ZY+nvi
D7AcYtTatamUtx/LLe0uXFCStetsBAH5bXWejpRhgJ4Tp2Tca6aEtNcnL/D0Y2kBd0DwXurifl9S
uVQT5F00i83Ax8x0najN0yYI/gifmHVrX8JYgwaHzwZbpqEkgJ8mk9TGcwPBxmpjTt5RcAsaYkfW
QWjv1kb4KGOt0KzxK/o29/xm30/K7DRE/pc+kRfI9OL3f6w78gTLl15sYaUgirvqPBoiQfwZv2no
tbrNu05qpmG44IuLtvWWmQOGs/dCnnufgf7/laqpab2TLNor52GSRXMWHzFI9HpMMp90kGPqhdyZ
3H4+hSFo1xt6ZFS7+MdsIl5tD7BVE86iqkM7RWyyS3HrhI+2JpJ5/+kj1BHE5V3hBWINpe4U/fw3
660R078p4a8AuIvlWaD9fhKKepL8Kq2AlxH7lCxWQ9LW8ZBUeThOh5QlF0Kg1glFYleH+BIZBeCq
PvZgXYDR+C5OUAVpnT+qlEmA03ZY2kJRAof4FpK1IYM8EHn+U1Dx1Gh8sXu9k3gsi32EaCsjYJHF
FxJop9rAsxwsQzJKcDbxfxMPrXYaxJ8CET3nMT+YeBsK29AdnkeALO9Vip11Qqi6FlTDe7rQRsuh
sIGlFs9qauQbeWHAaNC14MIwoGMRSkGYIPf9QwY/+9Am3tSJs9AV+c0V/VhE9tORy2R3uu1taPUO
iL+PcCKiHmLq7L1/IlwyQHHCvU77IwLG0187NnHjtsMOFlUi63I2MUfjnuiAs/3/zMEIdePiAGH+
/AP3vZe6BtqGGfoYzVrTRtbNRXiAs+lO3yL7cUp/45mhNkPPk9NnAxGB9B39gc89Nep9h2HZQh3S
L5hbtmmMHdz72AY3LtZpH3ZLyB41caHfzDhBAZY5XPFi+y80i0NAp6gesntGBxOEXXyFkHleDh6b
YMpcX7lLad+9Kj83v/+NkjEE+8avOEUJmk4cG7xkQL4uT2fK4kA/1caZj2L5XO+5UwNJi73m5kVe
RwjAuDS4F6OV31YbTgzPp57GtHjti3/HZJ8Z+APJv6GtfPXSPisnYqisiT1NYS5FKnlLOZROCUSR
C9kJxcdQm+Elnc+SpIi4wERAdHgRzB7dhlVniRgme3QK1CZmkQKFocce1tT1ujEsxByffu7wI3cY
bRJ6PCIBGOaidgPZd6oY0XvX3kgKuIrpLajPELIzyjYjL2gmQaa6csZ8aZ1LMhEtjRIFgLrvlCls
cG0c8dI6vNR4lpNAdot9oA01tc+yT8gTfVmUuqLXf8I3EY7TWqA2oPwIh/vhp1fNzHk7KWlF9U2A
cTDIKXCT5UHeKqSTCqDNZruXwk7qJW7rqiU9RKpyXPQZiluny/rkhbv0ox6QQq9FFZ6wFXjJ7lo4
yJ1tBEndSUWss/7uH5qPl8cWGqzNDRRPSBhGHbWDxgMU57mDC2O3PzC3ESvNXGLH/3hzdzTxeDub
p+I229DUy8LhWs54EHcHlJuvq1a2xL/g61jyYetr2/Eof+Ezm/7u/90ztt6VeF138fPx0gqA2DL2
aJhM9Nncb3PXOYWevLTfvpDT8dTNH4JQg3MXv0Psyzo645BN5ZCU7ynPxcCLKLyRQm6f6Drbneqt
98L22jdRXnnT1ozyWIfCIcOt7lzzPprHTS/X8UjOq2pMWgqqfmlZGXt2m7LtoCgyP4/TsUxuR5WQ
+Ouyeu/XhqoW9mcFmpvd7ZwRuXFbpTU3jfi7C4qvd0uXBcO95s5UMzGCFbtUesSYIlWQvMDbqEMJ
zsx9bqTeUFuyuN9e8DRMNrjKAE0OgmDipbKKzCC2MJ01VJnYM92zCCZNffG6PE8JuIc2EmAr1Wys
bSEoWJndTsMoucEAuHAaOITollzK0GXhxUaOZPQH8UrggqSmYN69Tm01VvpfX2L+u/pnHJsFAEsS
7B1CCbXCN9t6/B8j5QW+ymHcZ8zCYea773ImUFhTXKRfItIZh3THq5zgscO0NQvL4ItBeYDkpxdW
iv7Lc66ttLmotXt+Tvjl7IKUAWY9BNBef9cFUr6DpYtPXXCGYGqXU5Nxy54bD6XPFvyJrHiOjR/R
cYI1/eFdzVHC+2RpbpAn8Jx3UPLLSipkl1wTBJtvHT+A93QceNjn3BA9u3+cy2jOFOC3E8JalozF
knTZdGbG3q5DUECn3pDkxh7rTlRFS+9VXoTGKT2mpKLD2j+L03lh9SOecPQTbmQ8aurMlqxUJSww
+F7fqe1xEDiJgBT0YW0jnNZeEoW0CCDwxJDaf1/RgsU3/cTEsL2ZyHsQPfNYBBceKDSE4NZFubbG
n7IFTSqa2607Hi6PtQrJ6efwkZ0FltnSJbH6MQUcjcvTCP2wi/cUJknvWUbp1uRogkjjLXdLpnGz
hDal3LUUDbB1HaOxyklMJHdSyVVSJhcO2KTKhcAQb8yFEzkwwvB2s+60V/5iRw/YHJwlwXEWXi7S
9N1fP33wIXZRrB7lqD9T3AQdEIrClF8a7Vgy51gpQtaF6T+uPdKaPaow4TMrXcYPUW8admFoWv7c
sxIKQwAm6IX4TylQctMXtcha4By9TlBlvLMuPoVh2RNuRKcXLSf/qNeDsBKfGFrHTLiRj2PUdSvZ
bIi1AqJ9VlK8dJ9IJRHk55GRNr1mTt2pXPnxpuaqYQ+yBio8hQGgBdT5R67RZ87XjSRllFC3b3Qp
6LQAlepQHHTX5E+yNhC/4TBg04+QPvbz6yNP9PY9POp6E18BL+2Z5rfVRPxprnPF9/moRejRrwou
X/1XDrsCSBMQ+wKq8gm3fFquDTV/hA8FUKwC7Yf+qCUUQexcWJt1kEA9tri6VnXtwak1d8xh/8rd
wlpwJ4Qn1Q3of1phBs/JwPhZ33IcQN1gy7FoUiO4ym9iXU8qcwtMbXjWjJAglT9LjqlG6+roVD2B
dTzWe7y/EKPWo5Xkv1xHy82MwNfYUpaBnAOETbSXBfTEboj+SNZwtA0rHkmA6F2pTJpCwCnxnPHs
8p0kNlQqqI7CqyVpWzBqP01rRXGo2a2BeIh3VrY8/zXEZ3jcx11qXVSUfnLrdWtyeKMyTVufG4Vl
LKTrWp2zoI3J9H4bHmb3bpBrZUwxkTituIreSXGOmnfkRJ35lwzQjf0BVQtbMnL2HtukQZfZ4FGE
Kd8dQtHkPD29lp+iftZ5U9zAM8LiCw3FccN3kvfQfhdb5aEQuf/EZmqTpiubsHpyAKUo1hJrJrsr
3jzdS0D29o+TTzfFOE2kaKsou5vkuG+2ia6OqUfb5gJ4dNnJnKGM4mZu2+9e7K/LcqZUdRUva/C5
RS+HyVTw5ipJEIKf5jU5eDAShL6myt3StheRV77iMgVddQbmU//IYh/M8RY0fwOYbAbamw545EAi
ChCMhVI14nukNcSHDS042q+BplxliLWDta4K+jfWHcbORzaBrAfJcqIXOFhGtCWJqdag1A8hJ0aL
SMf/EuL4WLXOIr38CmsHkKFohC+EmYaJze8EFPjm9/0e7ec36rfuWLH6wZ4DywwpST+cPG2VLIuN
FoD2wK/E+eItVLnYJFVr1oyh7/ksa3QgEhdIMIyIvkO8PfNih0mz1ULepJVW/FdE0IH7SS7x9Bnx
pUMy1amxeCWNk23jO57ecTK8wKH08HS3wWNHpnEauVaSxxMOJHKEkIDSTTaEtsNJKY5eqKPdaIxW
ojUb8Vd/MEiKmHgJrkaywu0kRsa1lKtTNZa0xP9O425fgze0jCbcxF2lggi9rGUSXAD51OQ8FUwn
ClOCDMFGHP+SeYBybO2q30EUOk+VCT/cp4tvYr32gJ8JNoaZJLluBRTjyuD7V16ZLkO2R7hpSOYN
Db/lQP89rnfsXttV8pBkO0pJYOhcbXNPfTxm7Bjl01YKfiynVGUywr8rRB9zgHjZ8AgHwHAEts3h
YJEqsZNmZLowMNefEA/OWjzfOA1rPEByuPZ5SZKBZ8yyHx57DBJ2Wa0Zqb454JoeEr8ZI0qV2Wer
6z+hAfPSz1V/lC/HDZ3AhwhQrrtLrej3nq6G6oj/X7fCBtk6jpMgM61wgd5rFlURZkZXR482FeQC
zObvA2tfodd6oAh82vSUmwxmnpmx1ljlvjUlvYI1Dqj2SUXhRCHr2UfezmQvQc0PQ3gczdXmMrwd
wE69q+QyCSOe/1iYr0WWS+DnBMgu1nIemDmtuEmgXgR52TcER31Jbf4nR+iLY33rCyLlZ4GlBxLX
hHldHeFrpTMpzii/RL+yrlLaaAuFXfBxC82mMOUmrLTMrXAdOvMw7I8SORaTRlFF0JoVcIgr9gqt
JLlOiUkwlwbLdaHypcyf5A4sy2+IY4/hTSjVB1o6If8/T8X23Ws6rBrAy+cQCEOm/tkB14tb577c
tbaSrj3fqEzkg5eQhJ3+l3HNkjYI1HF+F8xcCb2qSebb6Q0rpSsKmQhi0mwxHWfvptKne3TDLGoT
psnKJ8l2k6fHzfcHEPia0AF1w7v5pABgWxbJzxMsOitgnC/TLd+EVgRMD9zaTX7uP6525S8IOR7j
agENjIFJaDrMME/DE6LjPHD+FR3bbjCPNtwNd0Ml0pyyPozLQaCA4oYMfCbdacC3k7wDka0P7jrE
miX+TiKwr1mwfFanEWuE/A0elhEVRcboxnNDRJi5b+pZ0QqlsI1O5YE35ARbckgYAtAcluup16bQ
mCavmm4uHVM7YcI3MO1e3QOKVRLTW2U7f6t9sqAj0q98Z7y/B19W17nbaydBIQ6FOQdbo0ws7IB6
CY0S2d9OQgoCqKh/uM6+8TXZsTawQNj6eDPiJgnL195cXNEajHo9ql+H7wv0uFJH1PCAkbuLIePg
rXi6160U37yG8KOOJnIGOlIlUlBAjrtbZ9IeqeEuIQ9XITmaNf0e8Eo1fVVihpkC1BDad/mtyu3M
BQjzGEHyfNmW/eGZH9FMHCDq7+Iuyji8XH344MTYlxEx8xh6JqnH2gJ9nmqPNLEoAaAGZkr9Lizl
U/DtYUNW3K+QKPr7etvixTOrqjqWfZtstE/zG1fT2xL4mg78s7PC86XrIFMw2IhizSuuu+reiLk8
+bhMOKI73kSbzIsVrxsWdrebjyoJbB1yK8EWA5MJ4UWtj8rFUufy13KwNykndvmLkXZ9JrPf3WA2
HaW31adyitgAeWsKPZRHaahvklJngzWcm3v8wISFWtmWbp0brraBnp0kC5FwajhqUxJtGAqaufg5
E3NgOokeRb1xm/32Xx4DKhqpIA+6ynVx7excX8OyoEJV8mFGUwawgXNmI+r2ZX7Uw2saZHGpT8QK
WLUoBYy0UPvN+14KunqZQBTVQw6Y8+bG43anF5ES8/6qbcJxdoBs0VrA+x1qjrpvYUfT/VRpwNUC
3OXVtiyKyusf1k825B/LR4b50WcSobps8AEFWmg9RiAophxuJZ/KSU7OHlBBzGIZegEsvzdAT0cG
tb9GZAeGBxhCiZowseZwXk+WKeaG2KSv/HKUvkL6YCmMnSucQEJkusSp6X8W4CzS5VyJYiT39SLO
kyWKfD7vrRXp6j0bSwWp5RU+ARdyyNQxbP+8o/fculv0f4XfBkO/7+MRPPpN1SEJv1otNnSTBPeB
Rk1JDKDGYPJR8RQw/hRBB4R7zwU1axi3VMOnKRc9zLhD+i20EsI4XYQ5SUKAryK5uYDE4Qk8fZXd
Dqcp0vgq88dtn0C+4z8wwStyLxBrcLej5azhnDoC5xGCXZppz6hkJAPKNoCY+p5Uc5nkMhZVTJuJ
w8S7brz7C9IrKMnky7J3IjpzduAKTywRnIeU5/UwEjeXhjtRexKw17q9uj5fabJd2JxGwQUX47Cl
F5RAt/qFSkMKmMCnoYEukXkLVCtFFCrns3d48ofRpgqSw+7TVzBYBhhHXSs26Aw8ilmlBtm38eBg
yAIrVbKUiwz03SneEE0TaWKCDGICo4GH04fO/RKBuWToYyDZz+3BxrCs+0kc3faEvpxG0fRo+HN+
ro2GgT1D0coVkWDK2DOe0HaBkSQ4LMIDhootCxEzIJBDpeaXjcJBtCpxhSJ7lbab4j4A3F73yxW2
ygvJJLl1uKSwlQvz1SLuS246icoRNutnShyKIR2E3HpAdO4aGX5fL/KzBr493XopQ8UWaK8cQnY3
xdOl25K8Z1ExqsNwE0J3KfSHpdPYkGbQT7RMiiNee+5M1Rx+UHT/prTl3CNynuxm1CiB7JHUy7xp
oh+YyAgeoIH58b2yqEgZJD6/a1Oxl0A6kE8LFVMSqUsikh4iL9LxBZN6L8P5cqPjLfKdTkfJ7ADs
EBok7BecMGoWUamX0WjBjqU8g/X3XAwx94wtuhR0SovCc8MS+ldeuSdVYvSvXcifJ10dxYMZq6q8
IGHzviU+psguUVMp/lCoKScRNG+X0bfV6ZFzfDvidtqKjuLAwjeKh9GNePGDjRDiR5XQr5hc6CIh
ZpcrfNCmjqABeSO+597kl9Vft38/SIIod8lgirIu20scPMh5s3cuyu31sNMLkHwTy5/0f7fHnBPO
cefYAybEN9EIf0KyroiAXn6Cvd+SlZVNKDO5PCEbJKeT0IudcJ9mDQoDzQ5Wvllrg433frAcNbeV
x4fhek15Ky+hoDtPECwBvP0M2XE/nRJlp2zPgd1FYR6Q5IH1P8+u+axRS/q3831ECqXT5Ym5Xl1s
4DAr2GTEE9sYg1BpYCh5vLhUKOs5UU+yx+ydYKw09TJNA6BBnPObbQ3iNrMooWEFVfv61/l4FFY8
bPL+v/tLn/zIyMFi7hRq1N99iSdtfngofGi50eCae1I1izqPNzF29y/jTOCvy1pK6ECoQtbmXY8g
Via1oo+f63a6BnJGEeU06BFHbCqKEAPwLClJRQnPCzSVmTCSAjcFNTo7KwQKiFu2GhQqOlPis1nj
9/0w74uWPmsKt5nJwZJ9Cbox24hJaHzvvUlaVKBLp3OEMExaf51/BLG8E+fnARyV6IQBo3HFBFVK
JRFpnDUXpFvPGXwAY2GMmSr04u6WtqIzbmD/P5o5XnRHMy5PT/KWUpC56BO8MWmCL1vML7WgMFfJ
cgw3NXYN+/Xi854tHFVGiltWfprOCSBpnutYjkzqF3fYOA/hNZPepkmJHBuCauFvUEU/krj3sSI0
sjPrdrV83x5gV33327uFWQwTiWSCIehbPOHJJN3horcEdsbxQDeZ9lvKb2klwvPxK5gbVgy0l2ZW
lNkVwFVwR74h91PxCdhRY86tn1029Yj4nMZBBxv5IAQqkZwUUtvIVdBKQ/1ZFz4BsOAG+BBlq9O6
ipiedjBWpPALSQhNqFr/t7zdzUNx7Fw2CGZmauktiglfnI2LTEGtU2vb7Ku4DMQi6ThEf1EKsL/0
xF18WD7bXNerLFtQsMam/I3T9VM8lY/hqSPniYVbfgdtxCFvICnfKi7Htn3V/JDP9eZvE100ghmv
NE16Z6GQC+SGnCbNSKKbEkF4D4DOTtI1c3ppNPOCDfxEeHXjVF5ScoQzI0n6WAvfUbfma0GDPTMn
QN/JK85lJ+GTKwfnruZe9NYxBvyKhmlTM9p/EQGTbJ6QaSA8XA0ImqJ457+/oFcmyxCBDAi7qn9n
hlIuciPVs9vbt7ulwQ+rAYH2DQBWwqcl5keG3LWx4Vr5jXqdewKIppcgRvFAvyuPke4cUZJVkseO
l9+AsKwTo/45cnllu1aWkUOAS52OYvRs68j94rcKx8c7uivUo4pYBsDXyr0OG79aQYLnQen8qedV
Hcidoi1zm6b5nb+FZMAVMVJe3II+wyEhsjMYNDtcFjF52kWlctC8JHWW24GLGJNsI+8xoTAiFGYE
sqBNgly3JNaLZWe8yFbc6R3YB9d8GatW0zF5jhiilLPfwzQ2XFogVKqo7ieNZZskjAqQT/lEvPki
WwJKQvL/Fi23DXxR8BldnN79uBiANL0TWW+i3iiyVlCTlaEJe/eqh5AVYJ17Bc+jEgQVgC+c2w6B
fCzsUzj75uqKFZG0NlaHZ6Fg0DJc8UGKUCtjjZoIXMhTDDTGAXZkcjcT9RfjXNf5VCQmRItO4FkV
mZsi0XkkJ9AjPumVJqMGmpgvoEcsrRImSCG7JorZY4lMLBxWacLzKyftGVFcQZHvTIrNxxS8Wxu8
MvwtbYVx+TUL+GNRTunaeGLMr+dIaaOExayWdMt3jLdE/kVPYdNIslaOJea2sUVd/Rn9dzRWBhdn
7YltFFFEFwfViCJqDOFPjEAOeh37Qpt5ttl7y2x5t41Zygb9GzyP/+AqfVJR4Aiew87WpW3E8GBL
A6tWLhoNqjPQpdOg8233jQT9eTWSfRozecSI7YrnE8UIrvPuxCM2GJzp7MaJg3xe/ffORXWGW9/q
94VICGq1oLyZRNSRyMOyOqli+SCwHkOAv/lYl3rMmg3GGknh5CRJmzL0Bg9jHWbYH3J4fsamUZ6W
Scj+HuosFqg51XEbfMe5k/Bk9G1XXZaOR/MQvkqOzPnlki8jbEavEN2ypVFYARuNU20VSfTYVvjv
5lIM8sQncuogGDOCz5r5jJDcvp8jBlVUs9svFb5cVIgn+fV5K0oIK/lKhRNPWO76PLg2/6QJdQou
ZBkaJoguEfmaqn0f30SfS9YOxiyowtldpTFhLkQBj74MPIt7aMfILPli6l4gJNRtPg/T8tQJAvgx
E2eNHyAGXefhP9/DjQTqWgX/Yh8qWgEKgoIDjhnFEyuXgZDhN2Klw8ky4db35v+pamrZjLS/J60v
ilOhMZX4xlUKFwVIf+OfUtKRXv3iDQiMU6q3xAoCAZMTVHrFmlmH3UnCBiUvNXbNTeYcfL30ixB4
hXroC8HkO4e9g9UQKtC/hyBOUYQjs6ppFbu0CI8JehsKVj1mFyE/sl6k0vJ7Wp45KMHcDJxUbv+9
gNR65rfBVsTl+xEsXe3NXZhcJ1Sdq6g5LKW+iN8cVc8t0LoqO7BHK8VhDDQ6diRf3iDci1W+25LN
htmRM7m2mlfXWqyhO1ENIaEaesqTs67Pt+FVSttUkVt2/C5Qv0cFtGlmvM+E6hCJmAzdr1++WIfJ
5UxUExMVJMxcNy7n1mDBBuYpnQ/3cRfUc2JI+Qo0NKaM6GDxVjkOXH24ri6aCn0WOkebaO5lFBkO
L7mbi1TM/VZIFSCoTaby1tOUoZQvCQW0TaFB49F5ISFka4+MRN7pG+X28nZ/aYPjECNG83jYbnWi
f1jGSHGoGbRMpXDTC2bGDOBaVnq2c4E0STebAB4FtKpbCnxhxIg2zLmM81u+OtHDlJxNYoMqwIVl
PEQ1IRZbu2DBbB2YT4ilmvwxr7Mijxn5zVoUgikFiCE7uagi7k+f2u2p4qpII3uatLlCai7ZaX9w
qV91ppti7lXqYVKtTiQetAvxkQFFRNdzyniBkVBYlBTtHPfbGi3b66eceSSCb8lPCO2qtO6rbAvE
+t0X2aojFTcvnsm0BbyALfJTo8zFQQS1eEBppae8YNqVV/VCcbRL1p1ttm6BV8ZKBni0FZJcRilD
Ly/+cmpwQBqrjB9TvtyELGt0lK2HH8flfWFjdf9/+HAsfJoQGSX2nTmW+irKJyV52tU/7lm4bxA4
UDoCxbTs4QbdXercAQJvBP2MPCaT+63g5FNT80GVrem9j7XrejE+wooxU0zT5uF9pFDWtGr79JBJ
q1H3CZX3B6z9GzKQziy4oi16nwTyOQ/4gzcGzrsSVqVgqO/8ePAO9mUTZKQFL3xDDDlYrjMnq8M7
o+X3hqsFLajzTSjmN3Igg6jGrBCbPLoTeAH6Qt2Pa0WoqjHYfGHAhDSjXvoaHRxjspt8s0oMtCr6
ZuhEMOqVKF1p9PmgDZ2y6BBCyJdApcsvbdTGLV2vKXhcmIduqf8Lx6itLQT2ONiIWniznLi20dgg
ciCGIUgBlU+JQD0c0AV7bkbz1nAOU3csPAN/IlCv2X3Dpv8HPZgMjWNUvHFKuaHB8JE4OalnMmt9
Qr89sLjb17LQlwSKgfpom5wdJnNCerasHpupMS14JywmmKtI7tgFtgAwF8SUn1wKDzP6ClU+mxIS
QHTDs5kBoM1GU/OgtVSsjd00hAxlbk5k/tVUhYlWRm4o2mVaGAyo8MsaufqjLJhAjbK++rFwJF3I
QwJt0Im4mzBvWz7g9nudyxiDWrphsbikWx0Ne0eYQn/YOGWsm0keOQ7WpuZPcIiqESd5Uvd7FTZ9
pe8/EiUFQ9xOyvfZi37JreXEtKjucJZTL1EFoW9IlCMrl8dODMS5cVKzQ2eH2kWLmrN7NrOgDa4W
aDGLju/cVahydVVthA+lK0nep9J88WPSXurZNdRNcZzn03k5fZxfkrxWFEtF8twBmUsgkBsYjhO0
gi69raWDSexBhotl2ZXDnpv/xreD0lT1AzRTxMh6o3DYpijk6Yvf4Uc9UzBYvVFYmnLXqpo3MVZS
iN8lB4sOoKXAADOBUFFstGG9LvAMfCEvVw7yxuVCpG5UMNSnT8dxEheZBiiA15fINBJa4a+rdPjw
U8i0OxATJ+WyRXNK9dmdkIy+mYle/s7Bq2Al5thZ31Nu3MM4rCFrBSCoQARAMvqsH8vKVMBNmabD
qKVU4cK55hSPfaAqRGp3YVI3MKpNfb52yBcLiowZME9HFcBJXtJIya8V2GCuj41nAr0Y9G9bCLzE
HUaDocVJY5yKrtpK6DQ6xfxVyhhB1mb/ErrwYHjlJJKpwu9b7yKceMGP2GWdDZ1bxG5QkwGlOJhJ
oxQ9V0wAxXg01pQqDmrmEOExD/LI5FTjMbrOnWEUEb/H5oAb9bHy93hg1C6acFZT3bpmkBZUgQtC
GF9paxGr9kYGY7cZHbCcLF9SAnwmI0ykZd4fG2Mc+LzkjkyRVMeGy9bYzmcMCZc743ULt7IrQ9Ob
j63I2m14Oa9sWrUgODzuTVifrpVwSdRQkUVuzV4Bi07hLjRutW6J2VZLjdwIUgACBQ7M6xBSn3Zr
W+v27LLSoY9OSQsOrrJcuXyyEgAaUFqD6nqr1YPCaJzzhc65IJeEE69w4EvJKOkHJA6JrEuJ9Z5o
adWo4X3Kx1BllubH6bnOexmQHN2eIz8OBUs0pBuPoPqfEnOl8faKsAYmR1phJI9K7jfImzZLTu15
qAodQIbWzn5723jhxaelX+2hNn/pQJ5o8J0j9PZ1Vk46kLMrDIgzHVlBYC5+41febPUlFK93V4xZ
UjmScRY3vA4Ptl/DPHotBP6wBGUibq/aWLCNhZGWdBul/L1ZstUxjo3usZlEcLEflDTf1B1IYLke
KNl2cfF9R3Jc2FVhkFDw9pnVpEPCiTFjNORj+l0wOx/aTVDLRuHaMvHhPLVhYBVeo/jpQXqYvPDA
7F6NI33wPt7GXbksxVyQsOAFsOZWCIIhDQ4GAFF2PCsON4HywCbqTHaXVO102zL9ADU4QMqCn3pD
2vvVJO3V2eS21FUukHw6sCGoHVxfySQirwWLgO4EIMS4z8ruKarjx3ZIJC4BNkV9bA3dzd9u2NBx
noOeRwcubEl8p63gtnxknXvE/572qHEZ7kQZx+1l82HX1aw1QpfUOL+LSldyDY/oDAhcAcK6VzV+
j2UsqddEhkZQBLEqobDGNA1oL+2jot9Eg3739tlU50H7kvebDQs14GuDbJMzRHJOSZBQVKlhUCSL
AfQal6kCbpk5AZMs38gtu505Toa53BwpmqRyYRFpv9TlriZbZqnHlMvCbcAHjmbJutV+mAHLDD7a
hIVMTQfLRl/kMVZpYXA/LxXX41KSzG4g18hl3U3rBo9qEsiPbrChquppT99rQ+O3l4PWA9OG3+hm
b2gcqwoFPwOmryk8evotG4iwx8mYBLrgfp0O59dWY8FI9En7DBYmIpJh08lJblw1wVcMMeLPHZ1i
MkQq6F5KOFkBpUtfvk9lJJvGfiQNANCIirXsO4xPIe3Tds+o3xIWi9uNGumf+94RXZQbeqOoDtJ2
jrEx1v7uBu+Yq5+8A5IHBmNGz1yOvMrO8sbHu0wl+wK/4O18l+9lqZelUyVw59pwIs5vXWhWQ0Nr
bWEOZ67xgMoG9wY5Ir2iyUcA77HudXufoDd6EU4yxj3fA5eE8/nreFxS9F3Z9rrQUdl7A7ce4S70
2kh8w65x3Yz9IudF7wcNFr6a6LmLUV7Hp08vM2fispbiB+NA0kt3tAxC8Kl6DZ+AlK3pbZ0PUEnK
snAANIzgjMPkRE2GcWKCFlwxqmI0il0/HSeKhLtRXs83n6Hf8b6RoX13zFaYI96kMNidvuitsEsS
oWXLtF9z/v9QGaJT8efkiMG6R6aodjG7+wqxsgU8/XbyFAfbuqB+rHluUuM4R6Pdbi6yTSs+U4Vl
BYIYF4vT0uQRKnMeRBeOcirTLwm1qt5tDmwjwCxHInnFhi65c0fYeqjK4IBaEv1GoBIxfhJw1pEu
sY74qkOmb0bnqfVMLJLgYvh9kSSC3t069pswvXcDqJgH3Xp1U0lW6DsWiFixOQbGAoX6u/rKdItV
tal7rPgu9ksYGiGcHtagWE3tDqslzPInGmke2uj9rVPQg5cfiN5+1B75IFd5NT6B4ostl0WhtBKz
dKD4cFtqpgeP3qVHbhA1Qck1ixpi8JaOoNfdhaEtvfw2mFZ8UwMteybnV9lZFGNFvAd3ZRULrcTm
7Mlz2JUQ+tDTTodcAmF36KxZPfpibrHdNvPb4AbThjwxVrDT8drZES/k2pS0NxdwQAWBO8V6Oh2c
gXS7j/UmiIX0U9TfeRmW5hgKABGVfeWAIZuBkaG79kYzrG/2dJ4ujTZdtWY9U11bfpmwFwG9aFMr
FZdooDqNvbL89N9qNXE+Bwsl7yrJZCPF4i7qrBt/8SVOafE6+u234/+wFtzmt+d81TRoNyaLdmtD
yiDxXVOw+fUZAgBS7Dh7oEY9Le9xl8d4wljsy6lNOkNZ1PeVTqbl5io9dXcYO42rX+SwNmsYT2Xn
+eUtoKpLyEDF39G9J9liiPpLDXPKARQYzrncufEef6oUbP2cRrZ34xCoS9W3PFNIMVbBb36ZmQdE
7wqsZOYo8HHHziYd1/UluxWIzFQi1WpN5jwyawgapDD+7pnze+ut2G+8ATIOtbSIva0AUIAYap3K
sDKEPT7kDIYFbAhSszeVk95++6KeWjxe1Bn4jeufGivziRhVAXNorN2nc2bkU3PJTl7dprxgH4XM
prKdordc5Fj0QOwyIJ9fNoVn/JpSREK1EUySAZypHCRAmYckH9UhVOEGw0pipE//KhYSIe8f9zzX
Rkw22W+Ugau5nGNOZEOrREBmdxFtUxPBQeqFZvrAqjOuz/eZjOCcgrmGRa5E5oLlRE/joqPuDrqa
ds2m9998nyxW2eKiogT2jzvk7N8pfMU3/jQ4qI/rWjdEdjSqPlkg//ZLXZjcYPAs9A2bblZ3Kzf6
o1NencfqAKHD//Rvruu0PGwIAr2KOX8YVkXLzx2+77RoLUJ0tgrF58dAYVQJGVaJlOVPF/byFQh/
vGrg8FaVdpKkUoiJRAGkipaKodxVyiJVvmZa2lKmC3VcIA1f9a8WkZ3TrfLIiGvTU8fqc0WdpsEt
dGTgyGXEVK/XBqBAKF+dku6ikY8nFk0qokrtcZM9NFAqcwUNMvc4LE77ZbfsFP76ZKX7fq/VnPlC
dKRGsP6ZSTPcyve2hQ+uGm3qDlMVHJqA8KfVBLrZ/y6Tr9iGLbEr/HM9Nooz9RY7c+kzAmQhe4fG
bJjejNdVIjGVZkqHsW+TsGVQ43fXvLKk2YXaJjAihPGIItyQsrOClwb7K2oUKq/q+QB5YJr8cafq
B+ooGpi4JbFeXbl+bOxWFHG2ybW90ROwSHPeaPDHguAsabRmxxXpxr1MrDia2+9JrmaupjRvT1RO
j74v/hCjd/tKVjezygainofMXP5BAoMcCFEOnG1HF2z0ESLqRck/YSZxOoaOfqF3vMCKGZ3As0U9
tKzGNUZeNivebX2zY6H52z0vwEX695bpj5+gat5ccysDOueZe5zHCyrPrD2lLGrWZfUMSmpv3/d3
ZS9qS3VR+oD/DwOJ1Aa1He0fzXcwjPbPLAIqE+YFXDa8OPyxBQOPP5XAhM5GxM0/LfCG5rmXhgEm
DVVqcB/tVdBxnwP/YqLa5ScYeWivL/8yAPgJFvpziDCN5oMxE6Z79JleJFbtSX+z7WTXXJdJgtln
vgcy4wNHYWxGMm3LVJquUyTktXlbc86QCVjMZMWm5eKjy6nlbdkLmHAFC7ugOGeVNWw+DpXiz2Jx
dSgxpMXT2hE4gxt6R7ERPBjsumUW7xKVU341AAdFlR6miP7j7xZa5KQBIkORLBcXgpcN7l4/Q57J
y98NHeO0+XrzyDzke2Ky1QLUJlQki/wT8WIHAwOPTi5sIyjA7sijsv8f8Bdd89qSzqMZtzqUMdR9
EXssTTyKz+26RAfH/y6jO2quD/TK5pOY3VNN7UfXWNRHZ43b28HH9d5BqVlE7d/cAzUrA0YyfH7r
1Hhj2nSIKhluRWqb1SJ6Xjj6Ms6MmtQuJf9jzzX+ol/d8YvH3UVO89eti71Jojk6Ws7NbE2+CJan
JywkWnEC5BFXkBfLt+sNDWjMMSl3/jYRSlfvOGhBDHU+tVkm0IKj7bpO7z/mZLTBnLLwXX7AUAzq
RaUw7aPYOeviDQ5eeRhWHuTauku+QdEjWhcCQ7E/7Z6Gc3WMjuQyN+nn1RAZphK3Usl+YGrRfbfd
RG5Wapebd8BebvKicfRhJAXbCMSq/rZCiy4LhAGpVIl6BKsGRMm6J8z0PWqUSBdkVG9eMMMPvNKO
2Ap2AudVc5F0xuaAiNzt2E9lZSime2WfRscYBEJYwb+MPmahtrfwR62GbU9lZx8YomEr9nccxARd
B7FJF29mDH9eMvx7XB1SJJYfGYssY+OZ0oAEC3W6qTBILIyRN8Sm7Jf76pT43ayqYNqlGlnnOQT/
RNU/oxmOgRDhOiP/EYEvcVWvhyEobc247c/GxCa5Nu2rAuFiQNJ0upuuP7ZHs65A5MgO0TBl5foh
vRLZv2BBjotkxWV1dLflaeitjvaQWVnV6gdVfMd0CQgtHK09ZninpYKTbSmQMPGa5Vh7qsobcIZc
0Z1TrrsdtJ4UPvi8xwwJHLJbHe5yQl+12/vbWWzBdDyV7MkzWhynNP7oYyA0lfaL1SSx6cT6TfcR
HLp/kzrCArF6Q2SDIpJZZjdzWfrDz+WSUw+OzMglFk07TirDlsB+Bry45ip4+VCYselIysKVKqK3
I9ngvHsLUsOTpbdHsuuM2O4IBe0EJQPvMgHhLtHjc2sIcDc/AiEL7T1SK2DYD8jdCUsSrTWJeruN
sq6Wpl+Wts9HoPKwWnj1cjD3AWqaZWgDXxKPRFJjoXUPGEDR2Z6iJMRU1VjQpMxMBRhzMn+n3LOt
mLZXo8lrGSaHTnL1NMHS+mzyx+NVwstbH0LPU4uY92dzkgvNc69ccYn+Ne/0tIan+aqKFquu0WD4
CePiR95FgSNN8+WMs6RalfYn0ynftcYeXbIYce+Ssv9mTUmSQxFHuz77XmL+UaTJtXNolYk1tr+H
CWNKJ+JfzrtmK/5rjn2FOcNzYTJNe5FspUSiIIjPBEEPe0gbCxNOStrHUVLWc9dJXDevU9dSAv1T
ogwQcHxq62hU9/YqCzqLwNzOWVQv9QU9+H3lMImgvuJc0XQPP/8aepzQmJS79NKhloCi5fd9hvvl
KMBU3KWytitqjcMtgGDDjH1IkZdvzmz5jieUYf7uqjv+oC/NReNFhG+kCOxWIpnuR6zb0J5XCrtC
pSZdtqnh1/u8iX+hKRCESxKQygdljeYQGARj8Uzm5+M2G9HS52fiM8dus8jkDR+aoHw7yqYcZnE/
HGfE+xWbzgHvx2bm4/DPNmWGtQZ+HO7Kyuh/SpkwU4dMoPgKWZC6Si2uC2JWxlWV6MiFk8x/RxeM
ro2tti1NU4oebUm5gnlCinFgjWh9Mfr9zEFsijM2ARdQ3G9V1Ksl12uNSFVCQKre8K/D6+Rlm3WT
ltncaeGPKaOmYRqOvZJObgsnjZgzF43A0VRYccwFmFOz6sLV8YV0p9xRrLxoW3NH1nOthQXV5cCi
w5L+uZr0PkH7/5F2R9hizCiwbi/NyhCnBAfa3FY6fMlZUghMfIINakgzHsHmLakwuTtqlslZmihr
fSwLt+MIfq9UnCJfylfVcyeEhs8ceXuh6sl+xAYIiP3LRldjdu0afuGIREumulHfZ/w0oq/qY5S+
MkKnos6sC4Zr1RbmExxqYfDK84gmrQHjt8rWgEUWOk/8Ef04JGu72Ds3dY7t/oQel2OctOgvxK/u
8HQr7eF85CONYldHoB+ejbT0yJ6+nDYIbtoelV/7R2I9KRPaiRwZpfqKc5m+fPIo4WJaQjQm2WzV
XdWIcCUrk9b80qjASe1AEg6/05PKkBWBG25qum6Si8nqt6xEmvblcIZ9F4gWO7kt7Xo1n8S0L96d
QNNrmc9Y34M49kcj8cBwKb7NWccJu5i9g+aDIXKL1W4/Gx1I4mydI9aT5bqmJL9626zko3MbSFlV
LRTFWDgFZfs74C8eyenOc8ctSaMX0ZOMCGwVcRs0KQZfDTiUdVzPewNbhsgg+AwVMDIr25wB5C9G
4HAQeKbdfUgCOxrBlEyfcxmRfLiJKZBVGR/0UniWO42oHu0vjClBC9HMStCCD4RUydNhcGi+dhnK
MRQR/h/EeCPhEHMiTVfboeRjMXQbnSOBU+TVk59i6sIaaoGn+6NH9LG+hvyloksbHOld9x8y/fGl
f6ecMQKpkoTd5joJC/9Uoux6+kAu5aRwA2TJAc1KWMI42lLS7GShFGX/KxA95T1lp5mM+gRAcz9+
adxbPsTJeDW95HqF0fmsSsHC0bdP1JdDQcaELbGD4HkhiwQ16JuFikH0ROBvi0qqKCMlXGi/P20n
h14J2rgRCBQ04ecSuzHh3BoUI+TEmx3mtfILzJ1Z3OFNHcf8g5SpMwFT2rqj9rX3wBxJWJfgnqcb
Bivl2l4FirWl5vw0iXjLSZbLAQxCOMK1dxzrKqIsHkd2ZN9Opbyn1rbPVBnvh8Pv8DxrbxR5TZbm
/36+xUB/dtGQEcaHG9AfSoYA+YstxeJ+VZ8tzPW0xDMtWBelbABmGaxr8GmtKTJqdwqf5jpJEF48
T7soOOfP4y85IStX8owYxX4mIbwEf1icE52Hbv2Lf0YVoKAtTSHjQjlJHYPXqM4K6qJGb9h+lDAJ
OskT41u3FRbdzFXjhMzAK3lOKqa8eVS8R1GbF9CCno71f/T2A1u5hwDvRWP2+de6SYXzZGa6VA+h
Qn4CITeXGJucW6dVV4hYJEBWCokIqcSIlV0EmrOoDvUOvu9+khyGoAWEQDfqrc1WhxD3S5M/OrLx
2pYc7XmLJcXI2vGXXyobHfiRAFQaDTv6xApUw1vVjt9648s2QeUEkbk9Uarzv5F00YuMnO9Zgujl
xyRU1ZP0Kh1vzxyL5rin7L9BmCDkHUEvWMvodtyhBXzMZ8mkD0lBTzNmKTMUw0xQgAZiKRyBXBhK
RHfsV8m7CnXIdwMFfLP9Nd7yMbuXjoqXKeavjK6AZnpxPENGuwwjSf1Sq3GkJvH0Ed64PTZQ/Kxi
7IU/pbQfBZNwOK25KQWK3H9h1EwxLU6hP5bEYHC8CMZd67CtglrSWuQJawc1KthsfYFIs3Tncgex
BZiGwNEttZPTumWgnProIKp0VdDHoTcAOcg7H8vcpM9C/fAhkjDLcAotrHasTs9gvfp8fYKkAcoS
sAIK+Gh9m0nkN+tvo2w4Bk95Zbxl+CKUQC9t9eY9hYW02fMHoFyXNTXAtPJoHw2eIC5s2twBda0l
ybnPTkfD0578F2HSQQ5RUmYvsAZ8/btwJQW2aM+nLMRx3xoVOYBrVuSi1Nx/R4TqHErO019DICi4
Xdbj5Z0pSkJtAtRslK+Ig5omjz7wodNDWlxGGOKuLKt3KmLWsTZRHeXMF/U5mb/dgJc5CmvQFQag
bP1FYtvVmfNfYy6QD77jJQlXPTZc07yfaxYA1kPBgRYfnm+tgY/gxKJ5+bcqatVON0Kxq7rpYAVM
eP4qRIOn0pBGdL9bSkpv6842j3uc8jFJrMdGaPyaeC3NnyZ8tW+n7h33jGUmaEF8D8t5WgpYGsBJ
XNhzlskPWaturs2k8oChHz9sqjKVQQQyA0PegtbJ+Fcxbk1R8aYM+nrzy84SGvyVedFGw1t30ckP
L+9l42urPtBS9Gp3PkRvtLQR72SRbKSVYslDkPjAd7scswEt7bTc3wVtVPm5hkslG+4NpvBf0tMB
9MZFlWBQrryVSfnO6GMlNBvS+2CiUrLJdg6ipWZk8yXVi+yZdxn7+gof8mnSb15tIF09tuqSl5CV
qVmLtdjEgLDRYm3xauWVYatAKU5bHm8DykC/LaeLAuGg3022yqfdv8G7G2fRJzKKDJKrmISLip0Y
PSAwDRY9JEKfoPmooqdknkBNv1ZwaQL8oCTN9QgKG+riaT0TmlG+2lCozqvj2kgrycqcisLHetnT
xKHl13tf/oa4tcbva2iyWzd74fPUZTnxEtmfR/lpgHwLiczNqKfyrT/3X5HlLnQCYPYbPAiN9i6H
02bhdtzBjeBzGszA94huKUcO+WUWT1DN1/4fIvo5C/VTgBiYf2Ez+Z8BnxP7WtI4HDxLUDUSg2MA
u4ek3MIDcRPOmJ9/dGA47wtyqhcTtF8k00J1hlt1PuoNhZ7UAkYd2+KrLwdhUKJXMIuc+NMozaVR
+dXxY2j/ymA7AYiOlnl8Agtfd4L4r9TC01sPnC17hJpEeY13anE7l8m2LEM9HmCY8DFyqhRBcNOT
NByhwf4nweZjwZ3VUcpjr0aa02pHU7gq0rL1g44zOA7iohU5IaWH1myvk8k1vGGtTve49wSQwtB4
5os654RUAa5Jan5e7cI+p08emF3wIRwkGYcQImQ32TGMvJTnTfetFbuyJhEAspgcNxO6Ex1OJ3PL
cw1JzwjIjAID8nse2b7kkEmC6ZQl+RCGj1E3Zz2y+JqgUQYbYhqe6EkJZrw3GKkhKXora5vIPVS1
lQp5tvGkna5S2/tMk4VAzIwysiPRgJ6trJ/7VhuUy+0YZMwrF4Kzc4Ej86mvXnbt84fK0tl03zw3
qTDFDi8icwWYic6hi3+mG7sXSC5hTpG3J8V/79yf0OksTRRb/KpJOfBzV8Sd/B5B2ynFjif/3OwI
FPAPfPDOk7lsRtTyHCck68ts3YMPmo8Gmekgo/NMvavpa3qcB/G0p+onch81Wrp/rQ4C9kKjdjNR
OZ7DSSPSECyUbxdIW6ZXeVj3egCWorV369x8YmPB7yw0P5Sa+rdh35U79q+CsSz8/5yZGJYpCNFL
7G3kstEZ+vbXMJi/ozqYXQ5glLR/FW6L+oJCO458THCXJ/Mv9yIkzu1hSYXa8ogZo59DELoEvbd5
7dE/5f0scQnj1vALDsr+gPaYB8YG99rWr0+3wRtJl9Y9qDtPPBtc39NTzybt0a+iqOF813CzF2kM
PnA2MZ1LFq946eAoW3chCoZaLKGUPe0r+L2Q1MS8obqIwwa0Lc57OiIWJVvebZecJeNdu9LgCEdq
k2XZTk9HV27JANu3kYHQh9QwCmwatGhAkemq4ADt1DWfYrJIeDx6SIDH8kOS5wtxxuK4oBz7YRsX
BJDOq1sqV1xuY9VdEgIT8AHiZzX1NXnA08d7Hnr0qZN3D408VS4if7QILs/3mbgjZBH6zfp4nqEl
8mFCnuUDqfO8arFZ0A669A/V8R+XZNbjFpggv/IaNkBSJEPvVxLAfTnPqQitlOTnMZL8COp8/BOO
1vegWSmYWtiMHm0GldTCspL/TGnwjsshKsz11Ymjo34ssUjO1AvxMBN4Put0k3F6+seeIeSqyPAs
IrBmn947X8VfWy4kQqKFSTpTPNv1jAlw3meL27tdTts21zZkFIeVchE85UWryTeoE59HsxTJjXFM
XBJnmnxSxx9kd9r9lrUn8UhaPn4tC9gdehLSlgNi51qXcJV1VZrnrOw8mPOzQlV/12vxd+JRgpiT
h4uxjQ3bMuAHfYVBngHYcDGLg0yBESIRsgx+OvQo/gvLTjxumX0D5yFr5EKOF1N1LJ7mEDMwl9Vk
IjF+cllxpnvrRC4sKVkcr+muYz2lGed+sSttKt5MCTO+p0VYt8GPIuIlMwYOkWMXdYd+YgOoFFd4
cBCyfxFh5wf0ShTwjWHtjOG9C5vhBu+i0W2wKN0s5Da/zA6ESYAFBiYlgUvX0fucjdGNbnIZHFDP
4qoTVEt4Aks2P+C+RlPuAtnQ9M3wrrZf77o/WO3ihFkut7+zqxD4lufKXR1IZ8ellMOOUBMswZhE
a2vIhAwl5x5fuwooE4zdW9s14mfhuVX/vWZEUSFQ9WK0pRQNIdfCp+HoWZvCrN6oe8SxdGPjmH+K
ftSJgt1hAENEyF++J8qaP7/aUmEoumntKsAaP4PThmw0BRRukyJ+AzzoMN+RLTWhOXPHEOQIqJXh
//FIezsucVkV5njs6GEZ5gTh3l2TCDZ8GGZpsBy1CT/CAez810NrFzy64NjyunO2nU2533XJaR/U
W46RwkkS7fpyYFXGu1a/6DwNGAnGzvBg5om1mcJyn2TJvrrmPKCHQQUooh+sNDO4GAzLSfYUAJjP
GojbRwDv0jOBk5kyOBo4dWOrm+XfnbMQOqsBFEq/LJGnvOqiY1ztS5gBi72BdIeBKT1DTKMfqAEW
BzeDITB/FFfRcsKXFAtSydrsyuBzloAdoTVFqXPqdTk0rDuuFN5f88K3nPSMCFSAvG5kuSYcTIfO
XIGdZ5SNa43Ir8iB4cdZLdO9Zmqg2oCqw8Tf+WaylDKVXP2uRaeg+rjkxULLYvIHnpYFM5Nmm5s+
ZVRqnRzYu8BwvoETvsP+yBnUdfH0ANy/yyVkiPEv9ZD26+x78NH0ESWAgaRDQ8lyv1bK/zjXaSqc
n535BCPCCKc4Xkbl8KQ/orMLiJZ11vQHLKmsuB5O6AQJDO8L8zP/aXr/kCVYbyejhmOKY2Xmi2fN
c+4HmruHyCtBHMrCLLveyt1cgeA8fB3zvM3IOFp2l25Euhps932CTikk6SnTP+USaOzLJRcoHCGL
+kVvyK20bzI37bcQVqR8mzn0zuxjnVyTf8T+2ahbq66lx0a/bkU9kTpW8lp71qcHwQ8HEgtHCd9A
EGjElOzmo2k1UI3kk1GQY3hpETU5gjEqMTFLxZDN97y4rOdfM2G+byD70Ge1dDYSa14luKeeoHaN
tFNr3Zp0YNo96OznfYTYvjjunoXElu5uVlFHIFbt5HL+mx9gjBKvK9oni0D+EjyeqVSL4rmdE6wy
G1b5/He1G+nn3G4fvWvgOjar/B+oxqvJ9RItMVtdNZgF10buQHwL30MsPx3RKd91Q50n8gmvBNol
i5KtNMCUzphkGGMCOrxu1y6/LFnrmF4CLikNRCwYPbl/cCyigmUzT0capdgWjisWy/K6kbmSXeeO
BYhsD3QWFfgTug79VxpfAH+aYzmuKhBBwWIVn1Sbm85mfpXvN9ntPQ29YPi6Ap0GeTcMBM+zpPPI
geFqaV7Cieo5kOIdWJR6JMZc2O4g7ZXwHwuWmrQ1qL5Cs4H2FhBP8py13zkeMd1ePv1ggWhedFqf
EGUg3e3aOgwIgC/Sxgt2g1M6pf9z0DKWdWXzONOXv3hX/B9OSDTuo+L6xNB4a9hNkWb9BNZmfccl
t+apbbYai1xr3TFkjNmyAOIaUtpThaGKOAGDWvSGqUZdor2YXtt+VyHoosvghf2pZW3ICRS2x2Nq
0QZq0walMsDGrKjpIx+x5VSg9OJ97d5oCU2ABUmzEpyzJxmAWYZeNu/y+q/r/ux6ggR/rQF4r2RS
eI3SiFe7HKJWXctQrCCFBnK9mpUNa9iYPfVpwvAvQNrDjiLClBmHyMjXqphkdJ7pEGeBiHq0CbEr
NljA8SdrGwOTCE5DjOOtFdZWI7VC3EsEcxtl7/X5b8HW/3kOIOuYQvsBAKM2y16F3oI9/SOmbNGV
rp5Eca67y8jtPKJuU5+QhdvTqgYs67SwCEXZwAbYhEtG7/skdHdBjbBd713GYA8L+lT/d//vfKSH
u0/wMhuuEBTPCah/MXA32gg1S3xRyGKIUxNTBChWAhRwdCsxp4BvpIYenShcKun8Ju/nWGgWshUX
tkk7Mwu/RbVHqXpVN5+A81NevZYe7nfPrXMHcvYF0rQb497kLR034GFJS0tplYMSbhkbftzTJkPV
PrxsBTJ21h7XCXgki49zGg6RdcVheEiJn2A9HLPsYa8eLP6BE2lrI9WrrI10c4W6oKRyDSUM8z8q
s7x+P36+9NhrwU0gfk39Qe/pkaYyH/SVTOJw0AvPrNnowo39e9Wx+RoyoYa024zP364iatS27UDe
IsdGyqhs22fw7cCV4Tgdz8Wj/2Os5MLRKu7Uu2qo1hStywumw9u0WR2Psb4LI7bjMaLetRw+V/I6
eSWlWbxpW8nqVvxrfK6jxSQ7QXKELWri+jjH7OfmUCnCBFWQtDfUR2b65CBpdEEfYvnIQ9/yUSZS
zse/YhEHbdO3HcDWvtDrzZzRhMRQyywc616CLkgPTqL3T0OnqKw4Bo7syGrf0A/EY9MkjKhIUZZR
OYmUO+vxjSpLayW297dOi8UI41NGpRNJdUdgAl0gMdq+0gTcsefz6SV0A9UaGe4XwvJdTpaSUyML
nzSV67Bdzz2MeorRMQ/qO5rQ7hSTD6M0d2Gdd3WztmFLM+LB7GSlpKwyI8KItBojMUbUjuJ/ejgL
jZOcs9XmfVG7QcY496wa+WhzBK4u35+2QsUsIqY1PAtNwjsyIO/zgQyYFf3Fxomik0ifAQKCNOHd
V5DfHolL8ZycuFL6dF599BWXouH8XWmDZs7OMbPhgEpfomucr+Tj5ZCGuDHHSz/DtuL7+g2QeZHR
eBDr4a5mHZI6g18ur5YSvN67OHq8SnjbgPPu47A+igH4WOE/SYiPTQuIjSGvtifK7R+3GdulnF+8
dFynaG61zcM2YehvCiHLRW/LzqDTvp7XMgBqFI3usx0qt1PNOwAki6bUeNtxZqw16km9Jl56DWlB
gYrOANEPTgclMVTG+WyU/G3wze0+tYpoBnOvXmb3w5AhwPWL6l21sz58YYW7ISbS0yoobfSFpd0C
VNe0epfy6Q0uL+aYPmklbyqc3oPzOufUfcGZaH49NCZm9UrRNEuF6Wfx2ZHmwV3P0HwSXCK2RmhW
MyzDCKCfRCy4IpEuxyhkEbItTCXRZXSVvlxpoiWAxLR0VQUF713fiXZ2K62m82D+xBebx599DRLG
fMd8rQYNzr/yLA4XWo7t3+W1r2fFAoRNicRNPZzZSjrg+Qo2juIMrBtkuVgdt7OwRsH1TyZ9zEXw
EcLjYKFe3GN0ZGOo5NPiDLU2Vs4mu0ZxxW6EEZeXnfFytiHo0zphsH42EhpwHHG5QTS4/eZVw7kc
p4tzXLkJuj16XkuNdsflARNeVxZgHjx3U5zba143KP+KiF2yrxd5/iZZ889te/YJcmFPcH7BoEEW
uaDPZFQ7WmcPNVRSBlacQC+WdT9KVH3Gmug5RguxYmXe0EQA3O/ajkY+kUyFZlAOoiqNBgc6BlHo
QQeqwvqukBzTJYAKJONE7WPjwx8iUZ+ssdW/x9QF24RB3CCPy5+8vOhu13INB+HrA8cV+Vkftz2M
8j9ncntDHk0krrOf5c8rzGKWunlYkrmqJlDMRsoLcqXP/iBifV/y9dyoqCrG0vx3f3toGyvjbwda
A1FHG6vta71Xc9pTPuwgXF7/vBrgwMUFMP0ClgsIMxn8z1hY9rleg7Opj1XMDlkvyMcnlIuxbNam
44pq4eyVmjkopuomqcCobgJBPcdWshSqOXU8sdbRWkCx2S72IWouK0xc5CYcCvSFHAP8wLiIGhJl
iNml9I7xTYRNgm+xSfuUgbbe1O4DyAjba9EmskNlGkg7nPOl6bk19iZcu0qCsDfqL5uUYrDZ9lsy
/+h7G/XMTjuYQ6e6JGnsDfOSJX71jZV7IXL3YFTfyYLUcv5siJBzlBtgMgy6tB7c2jY6/XkR8QAi
Pg7mqj7OOnXVkS8DgotC7RRmLlljmSwYpiBpRI2nfc5Z9cTxs+JGhPSzBDxVTSfXplLKFWYfgX42
rY1MRqBRopDVVaNPCF/tbW0ZohxAKYdS8hbZZEgzwCPL4wnOuIwOonR1kFEOn/UhYJFQlIAXkwNi
k6/xu/kzBLc7fP3Hn6usEqdkCf/unsKnpVer9sbbl6HCZwDhjkGLZQ2qCgUxkDHc8QNiAoRx5Ds+
OLP1gGqHR+CwFCrIoF2WhV+7kTqp9vSFd0XneHVsZbJ4dwzyypkRhFJD/FR2fRD/6WxdFLsVLtSb
ZxNPuZaN5EgONS8wxvegCB3WhiJy1KONJrA4hMD7JU8gwHGNZ5a/mKzNMIBtLiNST0Y3JzVZvHqe
nNfvg/p1E/RHcn6AlZtbIFGz8E0QcWUCwxURqk+WaKiAnKwPHASnUV8ntgcAVRZoKVMXNKum3SNy
82HcOJR0QujIbawBVP66mr0TrsU96wy/4kmDMytDMrEZDNjbOcs2woh3KqPheegp36kzUtdsyTBW
qNR+5w6Gkp8dp+wSSfEWoADvMaTPpu+184KEpt/sVUiGHQ2U3dehMebAXhi3YWEY/kYWVOyTIKxA
W68kE8HpahbyREdU/CHILPhdijJEojTweJAGx9jfj5KkxPdsYL4SlpIStaGVAwa4FraFdJAdlm45
NzxFrL2/ZKZDmFdiroBWboFT7HihF+Rl8F896Zd8iCstNkVAvClVzh5Tu8X41/sHsrXpc/twzRJw
0PmgBUrdLPOYyDgCmYeAmHj4F6Z8l/bQYKMWqfS1vrdEUke7UhVdvK0s00bSbUJKJASYePez7BYI
pBNzljb8E7Y2Bnx5ZFi3JuKz76ULU1EsmXeC4K+B75H/sCIl0DRFWN2qH7LnU5u+pn2CD5/0NdFV
16Wx5BV/JNCsSv/sXGQGuunlZRUpVkpivB3ksmhUBdH5jCQv1CRHRE837D18sJIjlwd+wJvhgKgC
HDnVtVskFn5UnwrNiB45KlExixrlmJ+bigtiSmAZTA7aRoLRJFElaaEBWajRXDdvc1ieZQt6rSl2
Crrg8ggTEjv2tuQZIztV46Sl8WXF6epvHsf0/MTYOJqnA/MLTF2M/HjaMkSBD7R2ZI5ciGGTJa7a
kbaIjZvYtm1loUfDkRTlP7QiDOQrFPhfC39eX9RcjeDJPGuj2VmGV8MXKygcBEvOctvvGAuInIqV
tvGSC8kikqm+uhqVXI/EaJQiFLh9UhxdekmAuaMAQ7VMWXq3Rj6uBMR/ifKrhPLcJTsd/ih123V+
q7h5DoEVe1B1LCakN3BkOD2Xb7mh9nb2N3hLPiNYkZzXvEx3PP7Uw9b9ucgCo2R1iBEjMIX5dDQX
wvi6mPkSXHEVbKjpVrJJLOhgEwaHWD4pNzVc2MseqJRF9n5R6LGkHxyU7mZfb4VnSI3awH4mrYJ8
kFyqTzunH5/Fatjwhyp82a1XcBsVYc1iP6JnpovWiVFiOisenEuIhi5rDy4NN/zTdS1AjGPXA0Ue
xSVONH+Uc8itnh09gt5QAAO7r63Vm8OBvSS+2jXmEPUMRn45s8Dl2de2IuEpl06wTZ4kxJnSWLZP
X17IsNnDQikIOML12IS4jj5ex5L8l3gKVcOkp6vG5uB2QT72E1M2FlaTVjksHDk0SP0jzUVZwUiE
xb6GzopIfkHSmyW4CJY6uDhsY+s5Sy6LSRgrAy1/JT+Y+2QzklIrrHAwgo+2ESTgl0kgbsj4Dp5I
iyKSF8a8B5+grocDPwtQXz0M+zhodNjRY1+JLSpt2gxQJSpCMTc3JSp825aakQeTPV1hnjLmDg9L
DHMKScXl0pa9O00LWPmA3ovSSHoH+kOAQ5a9SMhj6eF91D1sL6Ichedj9XeDHI+qOc2ZgDixkWtm
p1Yb0D0tiHmYq3HOsQpb09wLzfJlXRQsTT+Oh+w5zolPNKjuB8OyeI6BdXo+/5qlYd9oRd4AK/qi
HO7A62abMa8TmEyzjqdvoUrL+Ie/KRGBwlFtiCXuPqj4fpkQz/0cpgO+qqNz7EJzggiVwy5SamPn
SaHH1810Y8OA7QPquvaB2ZVS26S+q7j+x+n6k2CSPxiafSMYT1gmfgV82jNeUO8w4XTfhKNafVnK
ntMUTBXCFMN0kuNREdpKLwgXUiAvIU474ccxlBu63ThsC4+xYyoR6f2w5LBIJDcu1dnVeKXb+oqA
w5OwdVN6tG8Q3Dy6zZVvVGObCNb5TAd8uZc0cqBEVr5N7+DNSvkQcNgwt5/5GsvmIyi9hxJnCYbA
4ZCjhlVtQSiw6Ld7P0NAEX6Xl9Xa8cE6Nosm7QLn3to2oDbNIRKBlkZ4N5+CGjhQnScyLKiRqxiE
Dgzqaf7GrLjJ5pw7BMyV2a9j2sw97YzWp682kXtwMMKHFVIxBpnrXAtLogcK33M3/aMKK/nveXWe
YzSsjsyZSr74wq+9cxQ3JWDX9j4ZoPX3e6+1vIbzUkO5aOkU9VYO+KozkZDWkv+UnmwFo95PpcRO
gdSzgleGCsASb+TcPYaM7qX235UIja6mmSYRbxbCm00YeO+491+RgZ3FedEqno85moB1c4NcfAcz
L33Oy6CSc9jhM6N1hqnKmZdr+IbHET98LxZBYNmxc7fvrtmfdCADwdmf7gT7azljm0PWwr984gIn
+dd35mfbS3XXN9DsP4ovgv5MXdOHcFH+ZjBz1vT701LgKzhN4akbfoKCT4ZdEMhBi4wBXEJBOHo8
YsOHJq1DjE0JAVSrG1nRSbeUIJahL9MQWDKhkgU/nQERpZ6fuiai57U/2z3mD/4TjSBtEf+Qt3xC
VkIVurGulUX85iwWZJMjP/lXPlTaUxV+tGaUmbUIOp4bNVNi3DidIwcu7JvB1KRS6Rw5YvZ33Dhx
IImPN2+x72LFR27pC7xVEfLXrrgcFvvyweY8LvY9HUIhwUSM5WnhnPnGwNXARhL16faDd8EIeH1F
TJQ8H3Qr9msj8+pV34AD6jM+vqGX5v6REtcJeZ576OF39yuxAziqkzaBywJrooF9XRZ4SFM7wrTW
eSxROQMf/yWh6iR6HU1eGguQuaJ7oOlnx/xtbShKIHc3B5hdUI0PcMGL1HoHSCorIB3wviDvsOsM
XLpeySvJG3qFEBbSM3OndeWjhBL8+crbitYCTw/fWOYmqt+7xmtYlQIctZCHFvt1tJKCYAUSqiiF
xe4GNeB2AL7DqUpF+86LdowF7yXUEYFAcRieBvIbFD0zB4SwYbEu8zkkHnkauJ3lOSZvvsIPLQms
n+xYvpUKP8IoWQ2J6gIKVEbo+PlWJbQeAqQFVFukpsXGQvsXQ2rwApVcCzLkHAPY5MDT04E/EieD
19QnWOg1QNwekmeoxyxdxJnzG2s7RVAcLHyLZrV7tSV6rEytzepTWzSnvEAWVNPfytXfhkMkBoWn
ph4r7WZaKKdKurwjVxkLax9fyFvneydPBZ733LmmEcopR6YDOZcsqHBmSRgws75vi6StOJ52qHnv
vRZrnAUZVZwWYi/7E+oTPh0oXTdVaF7LHxDA4yJDsQx19ZbUtFox/zi4Qr2qMtmvlDKuTEHVPqvx
sQuLYh4N0nNgfVrsL6Ck3BTj1rNiICj1yiu/i+LstMpFrDvMLnx0WVeYiLrluusG02fsx9MstiCb
R3fi+NL6LlMXQqur0HzBU0KksxHLdyNNoNMuXyVJPeG+4wuSXKxq+xsEgOKUn7SHWONRFzKRv68Q
yFtg/FuwStrqZPt3hTxUsWylxI5XnMQVZKFi7r8jehNOKQsBNyKn2XmokeVTCir3lR1g8CoR99WI
DMRHYNaPuWsEXCwHWO87MoU52A6XvkNbFxG8oIlBVJqRxXXf0CMkg+SzXwr2MfDp5kVaqXjSP5Z9
iIiRCtBOMbHZ8x/JbX34YTgVOQeAEHziwceK13e9Tbie741VoJvB2Qrupb+eH8GPKznldJmUu6hm
35/dytgGAA9BCURt9HrxsBbtnxlecLC+wVWwGLxPtSWpOQbyVVvmJlZ5CRHXJBrbxLABZbrTEPiE
6eU1ZPi9bolnDCvTK5VXl4tjXWVll7eahuDfYbflQ/5jk/6CocHSdFX046HGa8xH4y43VjaLhClH
M4qIhCupEwPot1Dvtd6Q5KppK6u4qEQ7espxtKumK4ADgk8r/WwZqEuHTJgcc4aFqEGYGyJAbjqB
gCkGZdmGn4RrPATtGwb5pnRYcQaxyCDqCTlj6KmZsLjCP4cZJlgksIxfu/ENePFYG0QU/cPRDZol
uVSc3OlS6UusPuQbdbB4caIJRRxK5JDhz2mlElhLvprm6lUsN5JnwhVtU1ClwLXQddst4coklubg
TyZID3ze8A0cf0DH5Zd4MN0sprhUHFdxyBT7bVI/Nj+c15xfjEpWfqspYm5R0yMmYUKc7JFXENtt
9xSYUGpG7Nk5rNczsa0CdgCWOm6nK2zblC6+NrbKPqrxq6AJXh+xHEbyP2CnPHrxZzO6XOS5+Nbt
BPKz4NTKXqE8+2PxgWUGMc//sjUXIRIY9BRVRmsITbkclBgtNcTbTLhObpcgG3b6iLe0RKq4gYiz
2tHRgQ5xex5rEYql5eHVo5FxPOw4UElfcaL3n0kAA/Kr133RG7UJ/0GLKM9wiHQdygxrrtFOuosJ
M04bHpVF05vtiLAbmyC1QgEWp6Xk5HkZlwTh1mycguPc4eDpqw8sLJHaYXMdj8l1/hq5PQXChapD
DalJbGGxRTetR8L+rqq/os5J9HW/8KBjPkE+hVZJWNuM5aZM8Lw26ay8iQVQ3srJP6VSC1c7g4z+
V12+Kj8SnI7OmsUJeStO8KsURzZV6woh+ZxXiUbGhUd/2bKtvk/kBA2f7fyZ3G402H/KzfOQlRou
q+zhn+Rvi1gwtVUTDDMPoz7ErIeSIs0pvdNiG8vkp4C00SvDWfcgR+6ZwYHvURA2wdGDaeZF0A9d
ytUbslFS6kawD059tUBqUkCXjNcVjvcZ5utDZp4i/w4iHyDMzAI8p3nWG8sDBRceN3hfF2gppKFT
yB6Q+7M8uqPbvgyZk2s+6PfIO+YfZ2/RMEs7QULtrTdnCktWvhN8XJr9bSxPG4s7fjgs00nRTStj
TdaOmMx/C/fh+kozhKx0yB+bzlJYfwQpgtoMw0M498Kj9cQaJuLHhTKtpoXr1tLGGL4OMG/oFn7s
uA2BsClsdmFL2p4T7iPE4IkqhTWUrpEb8Az9Wnb0hSjmpAwnkAd9BaoWlcCO9hXdIrT17W2/6ncQ
u3E2oHiUfWbV3Rcw7GiSTecGv68t6NOQY8JdBw/dzRUEjERIflZ6SHdb7WfvQmUm1/MFEw4qMZmq
UMBJFVxM65QSiAvbrTk8zq039loiaf8U32tHE73wcjyF6prKG0dyYPQ8WbFvrl9MK2LLEjV4HgTL
WqL4U8jmrxUKl0cLKnnpaVlKiYcd8eZ+2ktDVG6olcSkAX43JL8/EZNOZeywdMt3NTPfOEwtFtoG
2X2yTb67utS4wRyRECWDw4PHikHNRpgA0mHza41Hs6ne0o2Ll8pGBvK7kyxnzSoROcJlH4CgeNJI
OztL4ghY/sjyp+h915TDPmHv696R6fMGmXuiX0AuT+N2OC4Rs5Itc1WwfImyW6oFEMCzOr1OKCtG
FQjtYiSK9Z3nKIQX/dVt82hfTOqvqxck6zqfXlipZuz/19nKYRQJWuIQZ3y6NjzywBiyJw6jIjih
+WM3gEj/z9ZqajY7+xL8cjf6ooDokfYt/E8a/RZphodZ9KLCf12WAQT5ZTqUKFyHH2r6JOEq26EY
m2BVlWr9ZKYmPV8bQwWKP2ULqAxbHFW1NEwLeeiTtoM/7L9utSx1chAsBOXYFSifxcdH+6Q7GjOT
S14hxVjmHG85ZSXNo5J1iCZfQ6MrJK9znfDho12a8mDF6xiqWulY5vwVETeunOYtJE4+ETqrKHkA
XD+9FZquS+YKw46luTA1GTwphz7UUF5FKyHIpebBwD6Ad661Zw+cEWBMwGB7fyST3A9UEVLSPIRp
Z21epd5A01x8lu1npjHj97x6iiSoslxtozK2zN+ck41WTw30cGd7ab9x48L1N1rqJhXz39lJlFIq
lE8J55f0mX1o5kjergFqwux0epZWZtulzjl9SjNUmgG9OFy9VgiZIl1LaaoUJdwc6EVrTJPGq/Jd
TQCrqG1a87aS/sp8VL0gduZibSLiAEmQG64mISDSozZT14b9Nl3Fe3votEYlTPa9Zk7SUg+TOUGi
cYAtPFZNvNus37euu90sMXKfOgmSSXr0FOdA53tOjcUKTMbGC0eEio/cgmXuZDsCQcr6RJ4LsFUf
cpLnU5FF+eqBGZ7TanIyFtjyOODNCWgO+vOW/AGwUG1H3rodLOtjQwwX9iXx/oAzj29PWsGO3zPe
eIGlA6jJFgk2sHoKmxWfGsewmxrH2tp1KekY6x+bZxP41k4rmc29rScZRv9Vli6u0LqRWePETjcu
s7RFt503ugrF/XxV0QQN3K1ILbmYjhaK1dcbtHyhrcOkWfnHoos5SC7ZB1ftYv99qhwnhMm7YkW0
u9G0vrcMz7dmwcViXBDIEwiVscrf8hpUnaAXQJRK3a9mx4csgbMeUJ6FSTII1UbKmN1/9hSiFjyg
1O4vdjNwWHco7IeNvMtZTI+T+U4uqRwQh/0Bzt+hti0OA8EXZlUWMnY/wUCWZ6f20Dx8AiVaYRRE
AM/XO70OzpRt8+2kmdl9/zmcAQ59+Y04rvz5PlEVd8FfORmQjjYR92HhFCVcNWgXunhGpuLLXpz4
wrZ9RlzKJxN4Wy4JKq3qKoCIpVTM5VmcMFc5JCHlg4b4IPXgFgb3buUGTty9+fqgDup1klY23Ue+
K6sYHW32JNswf3l7OcDLxTyqWFB94DwBOgMrNZKz47oV+7e5P6KyX/tk0jU39ozBDy26h0IQzuUs
X/ofF7ndcSozdwPPHgUl5tGe/be8pQvcSn0Zjkm/KOE1Pys+j7gLvMxlegCCFBwHX0rGZDZjgC2y
G2EebDj4FjxLA02/SDeholpi9CsF2GwrlloiNror5VVp1xpSlpy1m/gEses/IamV8KXSO0SduSNZ
Ii82196sTNhcgpaQlCECCb4NBKrUE21tHi3L/p7yh9JmSGP8kSwmDPZttHLB/E7ubfBkZQikfKzi
oTDTT4/d4twNZ31Vs8GclM0LXyH5KKpvoJoJbCTeLxZAriWBQjLVK9zchJogZm+FyddtElu8fR79
ZshOC06ALgoX+g8zpe4QXam9L8phzIWQbCOgqNwrkmXTPaWMTI91JkAqd6KfbWvMh7qKJwSPk7BW
3LvQMjcGmEfJAfEHE0HnTxdGulW+5M5tM8RDB24xzQwG5ehPGGHsYl37q9+Yg1fyAJ1UbRu15gyb
W4XsbgckPPPTUaJYBgv5JPj7A7sTMEKi+V8xLBgE1+bZ6XRTiclX+jlRqJrCRNH5Hzl5X52PJ/mW
PIoUb4UaAUHEIE2DFRwdgTAsNDZkvsXzuYzmcKPy5LNRRZZjFRnS0eUcTM4zUR564zY/Z/6ZARg9
uRxJFFsbVGvoB03+hzUZOJaiVLO4Y2HYmqBx4RuCKyFTNXzJ3Vs2GvY2Xm7keMXIEuKIwJ6Q4gp4
JWjWfQ3twuaAmBUkshE5zNKi4X/GMHsWAgZB5DasWGScolVjQBomc/OfHeS3IirTbGHJsrJOtk8g
9px4F6ucxmnlUSoWYiZi1FizMq0a+Uyr8y20Zwjt3+3ZsTUwog9v9dc0KQWHpFlHHYHl5OlnxkAk
okZf2JmB3KhUIzPSc9J7gksdzy+31iQdYhVRKmoME7syYogJZwVaQzvsh/LFNPho1nsvEhx/til7
L0pO7uOFLBLYS1c6uTkbWEi1EoHp0Y6YFK+ibpCxPYlA2OSWLBAD4HnXUjAI+36/Ex/r4hebaRrU
Va6nDw2vCECEoVfJSbBsKF/G3PLXPKnj1SBv3X6iYcCaaqXzlJmCTy06Q61PsG+2W0D/GxNKapUx
gCpXc+SaRN6yX3YUCNyI/SEsrLpEfgXfJEaAOVxT4HMKXSB65CeQoo9scbDLjmk2LykTXC30dzXI
HzGeqirQm8mWz0VsYM7igOJW8ThAoo0bSAx6awHzvHOZ5f6UCoxyi8uwUoX1JGMDIlpN4IgQaUhF
TElaBm7JwqSgpmOf0nhAnst6+0Uj/i8/9WqFZiHLaYijXfeOlEW+2lQbO3Uz69vLcwDW9oUcIRFt
DXgPvUYK7htzONuz1pLq8YTqhD8m+OTI9Latxt0QSBzKVvjyF3UkLYa2s6Stzq42RmwuwMULk3jZ
t64tyGO/nwHJgLO5WA49i48L51EhzVud3IU/6xlMXOSEpfoysx7Xzkg9huIRs34b1hDOCBdGKSxl
xMwTU98nwsyVdMJBIWoC2x72SE43zfg5vUwizJ+M68aHqhg15/Uf7h4aDFAXRQX39eeBW7Wnc80v
8mQgNsqFrZxMlB5uStPdGFQzmOaDkcxKEOm3sqQ8heymPfw3XNVvZ9UGCFjwD6DVKpLcKPr1uPQq
YMzgTmHJEGHCJFiGvHz1NoodOoLumRL80UEigN0SayB15Z+qwYcekHl5z9f4q1v0VuoSp9z92THJ
Xnuw5+S0iQW2o/WfnElgkbDvJ0zB7mRPTTedb7psfNlwLSpgM6vwPHC4A7zIUFWh8y+EclAWGDgf
3au4w/aDY74rbFSCmBHYuWWPGYROVXQC3nIHCBO+wXPNVQRBiyWh0A8ZiAnkTEaKOve/fbnA2Vsl
NoV7wcDFnRbDFAd86L3ZOdZnUJ0lJ+QdseWCgV0+vxD/qxOuidkpPxjKmgndJPbUP/5rI5e6AOaL
o7KxkL1CcoGawhZMlx+GrJCZdgm07TGgq/+fcdAo25FWJij649d8UFQs9firKLg3oLLeRuPYlfJt
4+RFgwUcSYqUKc0xCe21Zdm9142w8kFf9kq7inJDgfxvM/8THdOENSVA5oImaxzQzeoo692cYApe
ejgbBaDrX9Kb3/Y161Xm91XXFEWjLcLPRVkLmDKo7vRsG3TXyhM/VNSmYTa8h2PEhN4xLuvJ2MsM
N+cTOMX0//z08SVTZh3gHts17tdvImYQ+qNJpVKFsy+czC6ER/Kt4Xl3rrqeLWciSRxt67SbIpMR
nFedO/zguaaCMG0g78jtfWRLuGKRz1i8B0N47DHUQ05z7fyzKd3Xu0dUaIWhxnq07+jiWPYcW30E
VU/kRBcYqnkNpVUUuhc15Obd3M7nnrBW9qE5FKrF8jfJ/HfxiMNMC8GiMZAV3OpbJZQW9WNk1b3a
GfHug/2Kd+66OoZ4OSRFtPaP8gsAZq5e6q85bhp3YiRaGjrVAGoAVs/Dn1TuZLjV3SaWEYa3qpJp
HYPq/uFEEEhLqP0NkWB/MyM31g2FdblWYhNnxoqo0Qyq5fEq0gj7/ddAEc73+HZV024stofM2SA9
KLXCAD2cX6dCIcoqYQebVD1GHEAlyGTYT9TsifogGxBsy2tgrcw9ugqAx/72qk92vmS3CoUQamGL
If/PDVvRx4F8UEeKVIbKUHSqFlsbqYCAkzna3V4cYWhEUSdLiW9icW4AaCr2mQmdudqTsSoR0ApM
jzMkvORZT8S1CXZRNpP/Wqu42xx/otRtiezlpZp2C7ZwgqObdTkdh37a02UkgO7AW6KkiYXtV90+
Mpn5khEau032yHBgG+R7sn6CwK/17bvVuCsvpohKwvgfs4OSkPeer5c99zh6vAeRPuZyMrA0JM7H
eZIUYS6uC+lW1241L9SerhU5Titct71A10YyU8HW2hv778zLXDLJdNybPpPNy0/acPk+dqY5nEho
YfXq4gbCTPhuRplmE0xpLoL+AjL+9az+SG++GlYY0YBU4zV2Y5BLVLqxg8VYHkgxD/7zuIF+Yrss
0CMPIUJOr86hZdBI4nnJWstwLa03AqL4/987AXbu2j65eAZ0TO1bWd3FA03GEkEYGwr2e6kGJ1e3
wQqALEpxYQbHQVP2sioJ+1yhNaTl9ZvDHeoyVFV5g3f6op8JhxKNztJ4gG1rpbk3WZoyvcYeH1bU
mCc51cPPwJU3F9Bq4tcMinEcgLsRdxcLXO6ciUk3clQ5AOcZ8TDYWuhqJ6utLN7Cc0cL2C6YqxIr
zMAETe0lle2IVR/+uQeyT5fb0zPz/KhsgD8VVoWXhlZrUdD6vEC/17bO7INy4s0BFBp4VElFWZ/m
d8GeJr9KtpN98oMhuGc2PQOwYi9cqgU3RGCHehIepnrH98zPEipt4igocbfc96+VptVe/Jcqo6CN
T1rOHF5VhnyLdOHzFK0u2KnncyfZsQG4gNoiPKEO0NCoPNdu5DmCVMoW7tDN2pbPTbVA2sl+sksN
w3P/YqYGHhfC+xhCOM+TsKOjxNjS6HKf+c5y+8XgUeQeuLRTQ3FRjm5n6nWH/HZAGYACpZpVuqdW
YtCGZLt3LgaT6hF6Uoc0uWwVLBF4Zd65zPSJWcnHqU6AVstBnKLkFTa/XZ8MlebmnTBSVR+EuAna
suRw5qBvCFznbhaMcAdEN2DegVLnftT4qt9W92YNQYMLa+Q02fFJurN3uELpsR4f11WGP1tJR8XT
taS0bgjDgNcuv3glSB8JxhJ2CcHmjmVP0kcEFnBPElRRBEl8ONm25KNknn7EvTYxJMgUVb/x/G7G
EnSMVc3jjVO3r5JMJe5LZGvtcR7YrAR/j1DS7DvoTJAvj+NeRHPheqdUwJFRqqXwk2GnfculXNa4
/JXM+xLX0dPZVVOXZZkPIu+1jnEo6xJkIMlCb1N2pnUs5zpDT3woM/Mm6PPjr4DruIjuXHOZkSlz
l7cfNFkHSRubFy69TX4qbbcfadHST5dDW7KqxlvH458z6YAfVSRiDsiLQstM7Pkd2URS/xVOECnf
LVZtqeS37FDGdzXvTlruWejRnOlKIK1e2nTIDJ9kX/Nrtxl5dY65XLho7sulabj0qiW8Pek0O4Rw
o9jusi4vj+SrPrHTS1thVXulz22r8yQjAR54gk2MACdAR1bqc4so9594ZqZufuWlUbdSvso9jI9T
Zjq7TKdW1ILALxfTtX90fyMeVmz+bbRkXFGgAIF85qAbOtey+tRyK8Bcie/n3k849esviBfEHQ/x
fROOOTTV+iSNyP4ONgOXFt4RHywHRNZ5oAuoGGIAyYLZdOTSq01qM0wazOIcn0Sdj4Vzb2BGbbUT
JDRuNyPW+NRuB8v5aNrHEBbWxdjQmSoppNCooKHmCxvm5gByq163AV6r02Az4IwRDru7A4320akW
miR+u9UQmv6SXPixvPt2CEk8cPjno0SwzBaO+XaJNo1B9z4M3kwc/KfhXBBzRKj1iS1v+lsmWzTN
pymOzw0oeNLZOFvUN9wtFn0AR5vYlutjDNj4iYPuth8Ms0O1Ek61Hs4z0KY6X6GnsQ5a8fUFIHtq
z3SpCfs3fjMh3lJ3BrjYhcRWbwtKpFnyzsG7VKVBXFVu0JS0k6Gc2raBZZ1WOfRJ1unSJ1kjIF/2
rYDWi1KwSDdr+KXaNfGBCHhCARIm7nJqz0sBnB4y0w1cbMu5Lnciry+B2jJcM+e/Fmvyk2IY6/Jq
jAzUrz2bJQP3IrKz/awUgC0QzRPw2PGyfzbGDpIAVXAfVJuBJInnwyBN2wVcm1Bc6yxFfedMaD30
ARzFoaLaSZlyV747HdfN5Xg3lGT1PNi7wTIXeEj2sPcTKTYASOXxvfrGWuabE5sofnh1pWhvwPvV
Lbb0gBHGbchxcr3qezDGnWaiCdGzYdQiCTftvVvC5ZVAB6NZz/v84IEvXIm+cPfPU5PCJwQKvFzV
uerfCEraXVgxe09BXrLNxrMu37eo1KdO5++dTxoPDvpu28RUXGai1o13q0dXltztomB1BGpebe8A
vnJZJIb2qbEFrglzYs/5mslZr4GrO7vFlWB7Y5jYylwwR48QYA5pdGBJZ3ylQOFWyTQ9cYtvKGoH
or1v3EV88o2J3c6nQLmHVXC1COl2DIoafMrxI1kH4VI7ReOCRLjV4JbtnH1Ac9cT/TU64xucF5Kz
zF0LZpHjiBRWeTgiDWFjUjnwtQjN26dve+CqFp9T8c+0I01QtaHTbtseELzmwVdgs7ogZwK2w5YI
88dtkuYDbIOYO3DXC/wlsmMo/1b/I2iMuSEngAJLGRDLj5oqZR1Vfd/6hjuNkhpt5Gbr8pVE8LHo
N7sewuq69MaYtGMk7MPXkjQ7VnAcDdREv2PXwMQcflPVYHep/GLcXq6d+OPXFKFoDdhtGEqCS0My
+EdGNMOoz6w1fIxdOfxRbsjnPqIFT9dVUjBDBzpi61nIKmLv1a/uJGrxCbSCcQt+HHEaWF9sxwOr
iltyqp5EWWp068aKJKGkfpCn1nuxQBydf4KBSFSBDRifUsLmX4V4R4T9Z8BeIwoA68b3LH1Tvhut
T13yYxgkYoq+CCXfQaB5HK0nshD6M1liZIDeje104ROHsBpOLVRuIRTyi5Aj/hHOiwcifkCUJzLX
hz+6zaj9p5QQbs/7SlJes57nMvGJbj3tOuOjh70hAYbKm+pIT1HWqJoG3Wvte5J9aoRJCZ/D4azd
IsKOHFVsIlSazwxXSa7hNUmjz/XQGtJX4w8wRpbIGBXZu1/RChGM9tOXCutoSX7JmqMY8zlONN9l
rj/FPqUOVurDwuG0+NuRAmSqEg9+3FwSwdGFCY/j55lvS+FcfpAvmKuFWnYvCtYMptW94gW9DHI0
lyv1Lr6clnF2WNhB34OnC1ITL6pNGk4lJoBYPJqWiYA62SG6lbZCjqihja98VqySPmzBBWpgk3pr
LkkTD3KWp5hWar61gZevZTFM2WcMCewxJWD54eRGZFV6RvU6qaJI8ODchVoPYXeo+8a/z3ZT/4Pr
Djt1H3FNdTj+hQcFIxj49fqf02goGmQTT9dLnZvVs+m3pbfzdHM2MdKJmV6jljuK4qR+RIVBPHA5
QR+JuE7NS2HSi/wDRmKoq1AsMrRBR+PCu4rob5tTikdSCW5y0RwG15i8k86J8/3HpE6p9hnQCNbo
YyQ9SySXRnwn4up5rnf2QxAk6febElOVOhN7G0xhYe6cqNHNPADeQmVxgMrii5t2lrwmsEhW05mE
jvy2D5SM+83D9bG3zEXo/VfzT/nW/ufVofP9Q0EChyaKMjo/fAa/5vAo78hH4gGdo/Rl0PV9fMFe
+GB8ivLzb6OkgAIrlGheTT0fZbwmxGquQZ79NXJ7cnaJkWN1zgQEBO0QpUccKJEEnkX4IIHGK6h3
p8hmSP/PrWkoDwZzfp2JKSplNhfP+8aIrQywuj2TEd9K0l1M+7zqwAme/ln44iDwlPtR4dBgXp3s
rhb68ml8ieefsGY0O3rE/2Jr1GY6kQP6Bz5vC92lEBg8QPgVFUwoKPdWVVbP6bFMTdvcLV7nF6m8
PG+ry4d/kOkyxKta+p6oAEmTv5hgN4adxVQr8XShUDrXPMHJFlIvXOil5C6EPWhqIMo06z30rSt+
WMKdSOim1+ZCAfVwcoOLfL9P6gueFXRJh080ppJLx+GYWNizofYGEoN99IwMW9r1PYsq8bTktaJd
Obl113sidud1pGUtxQQHuTL48guOPJPxvLMDpG0FQnPvNFb5VPg6Bk3XHbZFBVAfqQiQIy0+o/Vv
1fZepZT6Vt2BN7HRBwK0u5PCmbZqvEsZuq9ezNqh+xSeNUBZnks1y8Z6xJ+FVahZwS6I3uK/2wjN
seLqQNA77hROcdNT4+cHPW9WvA7pDvDt4YrF4+BxJacmHWMXC96hxVyDTp1yScVNjEXqYNqHkCtI
ae1ue8XTJ8gYgo5pDfSX4y6cmlCi9XAVSXF741EUMfRwxG1xY10tmWQeBRxcpx22yNmUUnThzQVm
gKswjE1gOAFaAeOB+z8ZLZJndH+woQBIqgS+gj898O001WPg5k0DenWsjxQi94dKD126R2wr6tou
ngX5tlpHAjlL0HLmWv0LCTiy3HfngetApQ4HrcfLB87ZRW4frOVb9aFSZvYm5J0nEVp3yTMhOXcm
wK9DWNk4KBsR0lLEGjIjqe9UmVU5MdV6OtLVxmd/7ijxXcxtR8FGrqqH5t/arU0+uqHeAxg3DLz2
fdk9/8ihZhZbjmXKDYXGdeWF3X9oE5DQM+6YFYOGJfk5tSp0N8RX/KzUyAdqJaALspfBlapRue3f
BRpVrnOVayE1FM39aoyzVY8rBjPMBK0nn3Vd+LV0kFd8q1O0zR5AcPKGbSkYnecCt18wQEl/FbZj
QEsTCstzNg0uL/vpj6+OVTHca0wYhtseUMnwm4hwZuKP6SblEy0MZRiBrhh7nzVhwPbuPmIrJE0A
2+cxW1DIawMzApg0g2IHnYbMAVp502aZ1M7kG3Q8R6LqpXkWj1iOYRI1duopSwDlLyfvAv0CRpMm
ZeLr1kczfKwHs0j7EM2EIOaf4aDe2oGeBU361KU+2rWTRZaNF/NtOXpfrk7428u7Ri5+bgvnOhrN
9iMQWQrHoYPZCddG2WYwJNoJluN5C3Z+7nQzACJ7l2kAVR1tKjfYqydL3F9x4PM7wzGB8yinpi4W
PKyF08rwAXtY3AgnziZm2cpb7PfpRQk9Hs1v6izYWrElC0HnHzcO3WRb8FyyatRh7jJ57GKN9aLJ
1s3VYTtOttndlXsaKYOe34j9RSBeSkt3GgFCVT7mTMf/LZHkCK7B2tAQnC+QKVjgrqu8/T6yh4F2
SbIw8RhqH+AEgh7CKlcijS5TQ3OQRg7P6uWNWuZj6CX4FDaQDz9ox1Nq/ucu4zK9Yk9i8Xp6IDYj
BFHwGxqJV+3Yo8LjwbDu0QHBOBjM3h1sFB2OYpBXNpNNx+NtT7YQWUNNRISDK5zPA24QjSi2hqzw
8r7Gom265XSrpP4QZdMpByhIeRiE65zbOhy9bI7r+E28LVJ5NltzmmjpOW808fpCyFq2IM700Wnz
7CWQMYzGYfxo4SBhTi7oBV6+yxnuo99I2FtlRmA1Lr8pulDvGj2gjshXdI+sqDi0TY/VoM/pGVwy
JgUHDBtudUaz5Hi0AueK3j5xoeSgrPb9ztzgcDirHhbdxQGq6N76/zjimJKaDL7Lnm7SILwiEFR6
MB1pQh8ffOcp0/u6U12AnjIuSWvMyntEMx3e987U9WOY+tSyMp0W0NdpH3Wtz3U/lDnCWRh0w4ON
nEL25EbNTBUM4cr/O8b3OuVhvkXQI6QZMS0HI/iBmLgWBe8Waj+Jrngnv1TGlCK7FQGx/TUSEUFR
cX1IekBSQLPTBMMH3vkDOXLGbSFe3QmDRD3JYR1EGilHTKh6NB2UiIdPe5nRXL88IXFDfw09Z3I3
5+hOGcTv2OTe2KQ5pp4SiUtOAsXndi7t7U2zsg3QSYXscw8Hh/1MZHvds+P6BFdYE7zmw2EQfZlS
Rc4jGwITXU2AZMBQMe8XnUXmcCXRtcNuTfCDXqsei3UlS16SHKFWEy+AoWBRvHWICeZQEy/BZoyA
zkm6EW6DmDAijQgIiFFqLhI9Lw/Ztqj+2Tm8N1gS238iQvb3jw0mQX8mqT5wF2e69PQIJBGxwKjJ
7A6pTrY2VlKYhfnmAhVSeQXYr2bDZzIx4jQ1hygtyT0jxP1AvD3ltsJ8FTchmSDquv63+fUPbd7t
03ddcnaf6ziMl1seiMrpT7Y8yX70IFTuwr1/2l8Lx8NvXPyWXjip8BzeBF1k+WWY80uhK5po2rtl
srdLBZER0RE+ky9t6KCbkh9NFyjnLNvS8+0CIQKGkjN2c2IB6FYKpgLDRxxFUcVZmLKLARJ/rxRS
2c5JRGWa9iCR4e/qChL97VCtbQfNtCb3mr2oeQn8y6LrclsQ4yd4I4Qv/RTRUXbZ97PwUTThXVOV
d4WVZvTmDLmQKPZJQ3BpfG7UnUj6xbgrFvV+i5k39psUVDz40omqJN/Ca8rBP3SvDuuDwZ1q1w12
IADjolhOfWY37SMYJ51WpP15HRR0PkIQYMhN7/BKGkNHXfSwPItU2KxSF53x4d65fFn23KK+kUTh
vsPp7/KUiRV4cpZf56Qmcc2M+4lMKVmbvLEkrqMKRS+UpsJNz3YpKwFrjkrzZnm/vXla4HTBA6a5
KV4M+NkCjQ4DWp5qF+pUWqTT0qjHrn6enZGhtS8DRMEVLs5YWCtgQRt+hCgznIyBA75w02J9Zpwm
tOn9ioWMRXrRlz+znZ/oSRfMoj/PZ6GZClJGZofWW6/PUnKuVOsmST2NXafabIhiHlpjorVrcRn8
ynjf6djKEjjB9y6WSeJSZce7VUqORm9F0ikMTs+19a8GOXBe7Z6pSUj/hH9bkSEXXmprmKEQRc73
9O+4htvxzeDQZqG+mOjp2mf21jUdDlUkxuPF4AGM3vka5oToWarqmWEPCArvyZF/SsHSOl1az51z
y6XSQWxfXF6k4C30SVN9oUQf5DYehal4ziBzKLo/yDhQfOR0Zp5dDHXahBry7LotQlU47nkkd5LO
dScTKGhGCih28nVC8gwErbD1YJMP9/SY2AmaVDpjuN4t9mNPx8dODVIa0TqvZHQLwJSizV7133B0
z/Gi3Sczg0pEgk7bzicUzMVHzBWesesxk+iro6rmpNB3yXiY6MDepBxonW8nlTM10jjlbZSmbkN8
ehDDPxt72T/76XIghd2/lrqKi61aFyc9YGfsICOLYR5lXjOd0W1plpjvKe5N9IqzwkgE9cOumqbr
qJHDUNmCltd4ePjDXtk812L7Ka1tlapzNiioGmU/h5eax73hjIrTrjfjwyAQubnxLe5sWuBw+gJl
yK11xq95S0LL8A4GB0q1AaIrwKasT+u4RvTRVzKEQi9TsCBuUvDlubC7mBaCU5g0AI31JDSdKyYk
5b95cMbnAqBC+okuLirhhJOsRFxUNCYrxGJrEtV423PgbLxI/Si+oCKgiC/usbiBc5h5aTdB5vpL
7bJNw+evTJNllmxL+Tq3lUEOMVBxHAkWrjwSs1iDOhEMmjPtpVGZptDWVzLrEfKYGsKUGcYWrxjo
nAlmwVJnReJVjewiwE6MDG+g4Y3KT1qk0TM4B+RczKHY3JAHl0baZQ7KJBcdUuD+gxB2g7Mmmq2r
KYp0uJ27vS8jUl/N2El47UJZofTrtFkxLfUNIbx68owtATeM5mysfVwXWz3RiJtTX/t803WtuErf
ZT8vVTPpi5bre9jKzQcZ/0aF69vWPrEdZVnZ/gYHdhVMHx2NwQKp3EE5nczXZjO0clpXVVt2x6yd
MFZSCNxwepg2LiQLVkkVEdiJup5eyfpYYwXOQhU+kuTrJI+DLPx682hk3BbaENftoI5oUmlNZqYg
Nhc9B81MmjZA76JjLKOvAPUGhNIR3jUaF0+scm3AzheJc/wXEubaMz2HGroAIPwQnAhJhS6dfKhG
mYLzzWJi0wjIjL3TrZPfJEXma+WnjuTUkQrmDee0eVI7cdxAGtVprykRnqYLUmQyyZdda4BsvgdB
dj65ElDiCSTtZCTwD/SfOB8lMeLwuwli8JCCkbbNiOC6UVv84xWtKDPINhjss9W4bs4MUjCokPtC
zd/y9babcVQQh7cRspTxggGq4+rQn4AssW9jPgdd22PCoDlxwsEhMDr1nxTRyYSQ5SOPUqCDBFtt
jbKVXaDu7Iranb7utmHYxFIzjlVnABhTYyD2noicjcwaA1Alik2NA6Ps3rrlHGE1b6QPuyqxthQz
oN7Cyce9T4KusTBsQ8oE3zb4+x8gyy61NAeVBlEZ/TP08+toWkNl5snEWXqCRbO/mCTg0406dpO4
sATpSTXjvK+hB8ySk/9hp9PUz7iSKz6yqlqlGECxBeSoekZJa+C0ZXffACOkry7rXxXIrx6mJ+9w
n1Qmo0QR/ZaeGwybicvkQDNKaQC+klCdEYadNUGWQ2czlqIVm7SlYwgEwkjGzzgNn6i+E79pXIis
DiibTp3tWCc2mzq4OCnFHC7IeDlOq98+9cW6mJOzg4jCrpFNAKPss8BWBtienmojT+cYReVbQO55
Vc/g1I+9DpCgs5VTUUXV2J/C/L7NeLEByBDy+XSQkUhX9j7IioLDOAHTdwV28p0QR1s8QGw22FpN
5UaISOKg59y0PkVhELcMWdlN+E3rLh6Rt66ByW4Jnnnj4m+hZ2CltyjfUOlc7j/XmTVydFW+4a74
ZMkzuxj4RhxiBCPHf4hBJ1zwl7QPYxw7qcqxEJAabXyjix2QaO/SeISCTcM1+N1vRByfE3c6551s
OsY+2/gzX36d4kBON7do5OsLMJ9Nv5uA/RJC8y6wJrymwPUA8a9Fn4VJFcsel4dEm5POiUYuNtQB
MnNNyyQcvOgZmwoAoEY0pMwyPVLwule1v2Is8xnFR2oYDwXVyu57EdRSPrz7wRkJuznSXznmtqGF
+Yk9ZQJl7eeok1ITHA7smwNgTNpESEGvj1nZ+N6GEexOE9wK/6a+KnNfZNICxhKBh0LsS0MCgodX
llfjlFpujwAp9QJ4T3eMp7KhR7z6sFAhcoOpq020k/8gg+9VIjn3/fBNXB1cRLktCjVl1mqV6jp7
qWQnbwhLEKc93/UdC53/0Fgk30yoxtdmLVgCc2rh0+FhriQ6ziaGn35rO1D+UbUBaF2107AAXcCW
LrnwRNDGXp+StYdj7G6Z3RLWrcP0KAYSUp+ThoDRZSH6MMh/SIhoJgymuAB8xhZboUgYkxjI/v4e
vys/+bDNDvFjsDN54VCwBI170B5UhJuKICUsQUlXTAw+l8wFjYCMTaaWsR2JKk0AmBLIetJZAzmi
MqxHBMDBaNW4AvVGTcN5UIn3KQJM1D3byrBiL/MrHu16n37oBAaWIAJxNtiImfBzHFAmSSfAUkCE
UUWB6kAa2Oz8SYg6t0EBkzSMdomtaRGipDyD4nMRSTvNqNoqdz8pqDievTx4lfchS9Vkmd0pTpnT
C3aezbk9IrrFuyVmaf6MEjNqlTXwaLerv5JFkPTBKxOF+jjiXos8p5ghDwHlQBwONfc0h3rYhkj0
ovOJdkCoHwUwidvg51OQr8STDjJ9n4moZZ8cCjTDv4I9hPvcrUP58kGDII6soz2AlJ99FhRyaX1x
NHLCpqd8JhtutuRJdEUtjDddR0ldsaxODta3sDxYzogbDDUS2HUUb534bDeBEygb8Fjzu6rmwuhL
2Q2LeJt3qP0hN1rr5MnUUXOtYG1WAy9mg4iFhgiECYQdk0wTA1WNVSpaunhbjqGIKlX12bqMpCvm
7yiLNvD+MQ6Xx1UipO1LUa5aAtZAIW/9pcTimCZ+HI0hBKLCf/i8ZrWi4H7r202amHnTnaFGURrs
JjdxwmvV2UlUMQto6sAoap0pxabIYkbeSEMv/jn4J3orEoXHVBlegvOoWHMrSJzM0jsR9ub3Sh8T
iM07iUDtK8Jgll0qDDmBioDmpXyy1oHgps2T38HFYldygC5Mr23UCShaBTsOnFcH8zYnU6h6Ghw/
oWI6R3qh90NuMJEcA4SUxGJr5lCleuLpyQZIIutO3T55fwTzvl4qvPsuqDJt3B0pUNIbGHSsTFYJ
yiA3dRwcV71CV9X9NNCDcPZ3YcjRZD3GVtBCIkFk7klJoTBx5t35vz4M9p2Fyc0WzDOW18ud3Zaw
Yq7mamSgYvV/L+i/pyjOs5qdmQic3vio+WRoNc72Mpgrt/ySxV9QSYMekBqfr67bJLIrcCNYwl6l
+ot6RhUkedAyOAdQfALwcWfzCSEBy1ImnJK3fEr5o2Twc1x1vMN3++8dIRMITiBO4RI67kAPUjKL
fTkW1h6qyJJCl6Jch9pQrRlfUgTaI9fYoFmrrk+H9b0K9e0bcG46S180u5IKUBNNC87rQ1WnUpZt
d93hcfoB0YFSYKVxUuS75d0wXUU3haV6/iZWRJ/e2G5NBrxlUu/SuWCFFo3DD9RSpm+g2D/f8Pbh
qFAmPQm1weYFbupKzx0pBL7VK9x/0cRDP6/bBTDsJc2vYBS7myAneWCP1bUCWaApegM8ly1UohR6
r5XJsRYbn/UZCAGaYUNH1omhESdw2Ai9ovydfNsDQUw/QZWJSM7AGfCgcVEy61EiD6gI3roPM75c
DfCoEZ6tje2M6SCe/MeQqrrc/K1gAqogNRLDq75Vw/CB3tjGYaCJTVL/7X5TQtzwpUMS6spFPKke
gKwKihejUckK2blnOnDJ7A9TPyc4Ob0I3QmPeISxjqNevb+IR3I/FUHFk0LzldVY/9F0WodBN6L0
qbe88MYlC0un1Nh8wamO5UrX6DTjrddTOqm7djSF+QM3+pCowVR1YyWQXPSvi2qPp10LhA2wQe70
CsKdrfrIPYsRuqyCUwMz6Ik3lSA4RcbRgJdGkHEYYEoPx/3YxjGWGHNixJZ5IDOX3v3CtqUz1m2W
5bOyn0BCfwK9niaJkWH5mnRbJKArrA3vF4WKp2uU8+0H2mfHd/WHQCSOXOhojYELak3tgg5DOPEP
rcVgtrLx7O9mPdVDGVjYAvb20nczJx3iGY1S66azG9KFFPo9krvEbDgrdpkhNHBxhr8sxdKob2jw
WqjeHMPl90jWPcurDck3eWCu6fWGcj98kW84On+IrX1+5S29QYVsC8BlfXGnhRX4VdKt/nOvbllq
WKlOTfe+48Ww4nox+C6EW2iF9lUWLkmbRudlNc7lo6PyMOiiAgrN1CnR1eA61/Oi9lCsLjtmjCsS
PVZsAHS90fn+Sxf6D8VtK8oph3PMPfKcuNxgN7F5ldnhAiL7STPqw3sSfwqwI4hJIXROteYU4XPO
Dqgs0yrTqXpJgQBgYVxJ+ugj6U2TZFMDELoDM1nT2WFbyR+91FPjYVzo4g+Maz+aYlH+B05yUUm/
qv7zIgnvW2M3fTWpQAjbntG1qXvbLNpONMKcTFE4VJ6ddCofZ2WjmWnH0bidrHlQJGBpPDi8gVj1
XwvGgkBb1d3proh+JW/3qNFDUw3HC9UC9Nabii0A672YCoVqu+g73JMqbxbGtdvdsTUZ0QaclmxU
GFOuxL+jBKpgh7VFdzIV04nDY63ISWkyBfqOcpWGTYJsYI181/JOSi+6A5ECIFrUzr3+enyyqjyW
WqV5W5OBSK2DrPTRd8fT+CWKvh0vs0N+17GDyQkkevGmwRkwue/faXullKf4dp8j7Ut5CJdnlDmQ
yMlXlCzg5K3QLOUVMcSPZW0gHoJ+Pz5RhpIl77delRsngohdJs+b8fPQDCLFqQb8xMTQUmTgRb07
bo07D5lgpWIY5Dw4c3a+OJRtOvZAdAwxmd9WRM3DxVFj242UjhFzjs/2oyGMeJuSanI4E3MS7kyl
xmio6VxZU7XJ0EDPVB+RJ3KZUGK1A6Z3JW9y9y8u2dejaj6TJTBvpbNq+p1ZpJu22KATERyAXADJ
lMaApJeZkeu24Gnmx4DNbkgQgNkfoecW2UpOEWFN43ftNlxkTjPwYMpCBMCfNRAE4AXJ9x71dy05
fXcWoL7oetm3SYpxeNTlYy7Pfn4iuLQ9G6kd+vFmhr5Ap4LxO6JWifJ/MkEpg+fwT+WEdIQR4Vlc
3cP1gi/CjCiSkWq4/VrrRkMfPROrChkVcWC6gnZNxOErzaQxYIUdfatUiCPLlwEaSXD/jRW0cQSM
CYFBueS253/FrOc8Z6dEZA2czf2+U8SABBQHKui650AB/79EjL7OXV4ttpdVXLoAuvV1Plv4YEhd
H5L+wgbjEOTySnJcf9AJIy7vHgHIuIn0ApwOu99CH1Nl69/3EDmK5eLAWPVhFUsfajaL2kJfhh0O
gFikRvnYsuwrGQR2ld4GNV8a2zI/uUp1xRAizjmHykfVpkjwp/JGkPXvbzlsecfNxs2eJC4Yugk+
kBUfsMbj8g8Jl1L3jlSRBuUyx71haaHleljHGnRksmSyIbM664+kNMTQeIc3CzfooOpc6vZG7bUk
K+3Uc27LGRZa8u1t3hl0v99rpy8dqhfdmD/sr4h4dAa1MbpUy+psDD3S3By++q5q1SCOuOhvry5h
L8MnLKVhbbjMZdyZHqDWaaVcRKLrw2B+zA0npNOjRngPECw+2sNjnohECgtllez6g0L3cNVaI0Tm
5v+4IwrfM5GlCO/md2aztp6mpeqjq7GyoA7v9othu/n2rqlrTh3MERpVS2pODb1zbPq2qWc+EIac
sd4fgG8v5cfsxY70BCQCkIPMxxoWaDZlXVtSss7QQ/OVznkqcwCPOOtfhQu2fI2UHeuHj5ccSNKG
2UTKy7tEoLmu78Su1y0WCcfZGj01DL4Q8r6pXne/JNlwYAjmtgl6HtAlEiqXsHftBWu5FWeL6HeK
PbY+AeQskFjiI89QQ2jzh8/glJxyu+/v9yCJF5PDO16eHdBhSkaA8FC7Bf924DvONh2B2BdDFCC2
V67bzCsyVlDFrdyySwlk5xSBAJyH4P/HbQnKdOgNDAFkxAwFrwNCemaEjz8Kzl0hdiXulT1Wgkh2
bVHmz3u6R50S2mevZdFBWqiqSganTYqiaUpYjoDGYsJsC8JjAla3I4yuwYrawc534Tg8YK9I1lOU
fOTfrN+1lrAf+g7gB0HQMJCexoWtj3NuRI22y+tixOzYxNEUhA2layd1o3HKcFDBeoGGwo1EDjBb
Y8/2l5Hv99IanS9hfTOFyDP3dyFc7xf71tE4yBiNARGi4TD0JhUxmKauHiBH0Wsdg+LcoZ0R5nHS
EiFeCh5rcTupdfG9Rvc/Yw5z2E7xMkoptiqMREq98Myu0bUUANMaTBzB1yZS7FHSlHdXRpL2b97l
Fc5xfocHUQ+A8GMEzics2Nzpz9pjegvmvBlZkFDwcubcrAqK6Kc4FBQIJIk4t/jNPuiK0YaVRKsb
sGlfxcR0QwbS5eSgRf3Wzq3GzYXmgZdMI6zy+xfbu64BPSL++dOORePudRnxiOFuCCS9JjFmL7R0
ku8OUe4sropIVx+lbLUSjr90KyAVg0ztbFfqSJ+rirjb18N4dbr8SDh39T1P+QB+QaAzfGGZ9J8F
LSWQpohHxf0jKgGWaxvdKjz3Rj9CUEgq+yusz36X0F0A3OtMnFUKxr92RYM8uPI7qu89N8/geWhc
4uKov+AduYRayEy34V58hdgy3+ay0Kj/hAO5aDmyXFyf715zJJLS9frbBN8YjkZohvtnWa1m6xHM
HMpCUZnyWPrV4anwR0tIHUCaQz+i+96vCxRx8oP8q2OmBZ9ZnvVeJXjaIiHyRoG6wUaX3FnDorxD
QrzO0J5QAiRxOdDBDH3BzD5/tl5+BjHQB6DSf3/iyEyOPiy3EYgNJD2cYsQEHktM8jQmh9knpCEL
6qA93NujbdD8Bvb2ue3Fe0ir41T5L6EPe0hpa8Z2wPtEHu+FgXrmYV1i64pkEhP5A8kG7LitVsBZ
tYVxtKl1PygNm61OF7wFKNTTAzpm4TPCvgFtfglg/TJ58WGEAUHJzz8d4qoMaTAoSWAUVKScKypQ
Shyl6xdBg8XrcKiUg0sCA+dqlbPqydhuUECVWF9li8gsmSOKDRsILiMGw3EeLZaRcyldPj5DepKm
YI5M18T9Y9CklkDTVDQLa4QVDPTYTzqNpNpHCSYJn90hbGu0vvBus+QfdF8fLORd5qLVXm+mbOmn
GUGJ4tMucOGQF2OTXyTshaoHilIFhTZ8IE919QyXItHc0j0NoJBvNcaOhoqWISXVQ/alFBe98eMq
9hw4ahFG/hMYMpXXsvuDzq11biZzgenjaeSpudlg2VJV+QsXBK58O3kZwClLtBn1hP7BW/obAM4S
GU6ikwguPQG/l+WrVqZirq/fbUVfK6HvncU3QjzekdT2qJLd6F1DBXIFsqLg6Y/ulXGGkWDpHSiP
ULp2EfWzuevmGhWO26JmwhEQIGpSGoOG5xT+ZniFsaB4QqzUDaYEShmURV14ws2cxOYSlP21XlhP
aPECEXE4afCd908YbwDVY43wr7wC/VPwHKwD4b1ic3M9OEU+w+4K4IzOS9WNge5dcH50n0pjhAGG
qY0AuZxOFgr6DDt1eKcA01rntrGiP8lt0l78396ENaIdzX4NqY3Eoi2T2DVH287GekcVqwfI+KZ2
iOXQCFmwjpIEPWwZrorI2r/o6v28pfgL9XwX47nzDnmdXAekD6KEO32/0A4dXZOmj14OMTwz+WP1
bVWrUQKu2j9C1F5XuYlkPVHWo4UEml3NwKFT20RGDAoLZVdtvG4qONguzwteZkLTFIzhlbuP414J
7P13eFl2227rH2uwg5ZdkmP+DPoFosoDscRbAdq4afb1ygncvVxddwAe2Fko8DEUzsF7/+T5+kWk
1cny/SEx4fHfL/oJWRPXJ2T/SCFGQzidNwKsjCTWDAsBJgFrolJe4kOnXFDCoIlab5C4Y/opxOrO
dWKSLaDXvonNRQZZq6fhXW816x8gQRhzfF12tkBq/Hs6YRHaPwDrm1Eh2Wem7nvvaIhqxRwtv5J5
Q/edeAeEUwSWAh3fXKrMf516JNVMVhZxaLqhxU7tu5iiPHCzjH0yrKFCCdYc8C5F8Di4KX1YMKRg
c+ZyW0z9HUuUz9rckS6J63bMjb66F77k4a2pme4P09+AcREjnLLcpJko3zszzDf6F0GztR+YdgjF
3G6MTcmjcS8xg0X5+4AVg1QAh647TN7tq9Acjg68or34A8V9QroLimYeCERwoAsod+g9cyqeFiwC
zzdRIBuoffPdUfceJ354DmlHnFZhl7W+sF8OXe3hoWf1tKCBEpqw05HQn7gjUBMjKZluwpt95931
t25vrOZ4HmU5byrA2Y6F71dIcP+5JDs44MDl1BaF0/U6vSfQMx0r89nwyoStZgsgmSEfKgunVmHG
iReKIHH8SwmhkKZ3HJuJTZ3jXiYhcTgoWqgwQhiMPExRHBao+sEBAr+8cul2rPMGu/JFHJA7y4PG
PYyPSY1KPlbksaM26EJwTJL3sAGhrOzG7QWcXcil2WfVvaSZYsygR02ihH90dW+fV7ycV4Fs5Ufv
z4Ka2444BsIyMJNeaZGY1KGxw4JdgXravFWp1bxPY56xx7tmPHBwI6pbvedhpACss/1MYF00Td9v
MessQJ0w/K3+Bv51/sE6f0LJQ2zrrADMJUYXFRgiPOz0BHx/kGAkIg/UoLGKUrdpPCzMgLQQgUjv
SKy0IlLF0y4bfvXIwrvMHSZ5NkBv1qmFBVbDHE3EumtWdRPne1uHP5xof4Z4/lGMtdV2cb2Sjic3
1RtFUj2ANMngDDVOWbwQkh6ehDOF6sgyYeolHOJ6yctmpvcq2BewX0q2nFKdFMtwObbhqKDelFde
u5rX3E/gYbITUOzc7axLB+Fbha33pibAq44l8m/g6YGB4KxmDbGKEyroD95vmf6HAMvWlUmLkyyx
OyRW4UkfJkPo9QRbL6ONlvdTyxGOvZ6G0PWLD7Aj8Be7rLLbCSjK/044BVUVOIiOPVZDrZ9diT4d
1ADGsdDaSzgQ9ZCOH1XR1RwiQyfiMnGKCVz5KMTA/dMvuCmcC/H68CJsUsCzzaFfydJ9m6G+oSPq
eMxqk9CS+Ch+lXe7cz+rbBOUqQtmjyZLcu8vGQB8kFbveNNFE/rnWQ2XRPFBQo+kRQ4xM0Qcb8/C
cFPxq9xZ7n9I93t6oJHdKdLz1v6gvTh6JyfFcPhk9ttjNFr3FkMAYLSlT5xAgAv0Mc046Ba/0gWW
ELa3ALqoXgbPswlJmMm7+CkoRIUYF9sQjlNbbBc7q9KyE5q/sRzz0xadl9DHS/hMX72Ssylsjvqk
qvU7aCN0zXqk10DlrrzY6yohdRB/YlSWn7pOy17Tpuaaj7TsdGf4Gl/1QOxTagdiLq7nWpiHpSNw
nj9l15mGAjZos68yTobSCSF61CHFDHY1kuzgtZKyIg1HXTt7mYvFRva7Q2EbB3MOp5g1TC6VmS5D
Ch/Ref1NacxXXH9/eKs1BN9Rk9hzneygK7plH387pgf+J8cy4oDoJlKyLn9LDTE68+q9+rklhnK7
GFickfTplocDIEZDKYd4QCdF1QO4rg4hLuFp7hLuBw8uXDrfVUzdNJOKkrUPvXKyh2UYn4X0BZGk
i6lM3H5xDbTvxKr7gsPSaLdKYVdaKWjaHc5sCmMbni4ZgrsY1w8e9F5IMsypcinMQBYleqMz6+St
34/UJTo3GJcamVLHxAZYWHICTA9b+2cln0o8bY+ZiDrjNjy0MlY4hYPWBHBVfl0vKW3INJ9TWJ5g
IxJNuT63rQJXvOEWmmwFGrALMey1LEAKQ6LcGQIWX9QDXa1qi073JBfWlhiHG3J99aFMxSHpBzye
dbA7zkEOSjEcM3fl5Z7rp84U69X5iOpqvwuFs0474yM+Lb0k5sUr26qGL3esQOFu5dDQBETnG7Dm
jvALCa6Elda/T9OKXW84/yZEj4YhiOLBD5dEJmCFmqsc3IpIwnnb7VK8mmn8vriqu29cVfNp+VXS
oZTO3b8l3Ddwr2YexU0nQGNrdGQv3twQHM+8xGdgvkvqdz2hEHAcLPyr1KrBr52KmYAUdkb/k4w4
MD6BrmCgvwrwUlItkv3qy5tRtAHfFFKp+L8c+fvBgfh1DvB7zQKcMgRQ4j5jYdptPSOxUDgdIDdc
CVyvFVU1UMf2Q2OnFxWgSZrhRRv+Ke9omCYGSMiWC7WdtPIq1IToyjl6uMwmFph+VUkRSNLhFYM8
XrK/y0XxLQSFJ2T3T3rBZN968nQK6HCdlw+F1smUfLd0dWz4ILQETy4gVSqKr/Z+J+RTBc1H5ezx
ILiovBP4q+/CYHGgXlCVabQHkkMeJTmmDI/ITS7RTQME0NaUsW08WONPPwmJe/ZXmuDMTuJPSiBd
21uC6vBSObUGUKIvhbZnA17v4ICqeJIgPrMqz3cBhy6Y7YpvhkOkHIcUxoQjJcVnuocWXPNToQM+
9h48tQ7/WxwU5AiNo4hjYl7r9WVee3FRHcXzFIcbYgPdghs1aMrYjaNnMRtXJx1qKqtUDdGHQuS4
Qb/Ym/TrMXLPCfAICw8E30oQ8bX4cAJ3h4FRvdXA2UUb7pEMIvzFxUkkc3fwEyWyeimhKiPeXJ7c
sOhZqO6TpSnXlh5oJpuHyWqUq3O3/U9c8OyzGJ3Dy2y0rAmtV87OwUuLNZWVy51NXR6ASx1nbKxj
C+RmOH82k33YAiAO8JIbTG9O6HS0FHSc2vZ1W9WNa1GHdSpiN6et7wS9SqgoVLEF+mbMSnSktDua
8rd0Rode04kcoKekkxXk2iMHFmM4RlvuNbWoLW5dNJyMRuPnbQKb+g2ZQ4V6RR9360X3KtSd/NE7
3wC14rBOcHae4NTPAoVjj5g4v+dhHs46QtgkOfCgRIiaghxkiU/+wMKdEjTXz1X65dlcvdt6prJR
V2V/ZQdSV2InnceDFzMQyo0NReyW4uCcXirYthCQsraduasEW4xwGYJnX50Cz++MY/JTVfc4ED+W
pR7XyMOfnHnXDS2iUHWEeistRVkkJ/DQa4bQXtPG3hL4QWb1UroH/G7jBaqN5yzaJTWcd27QZBZG
At6vnM0KQoM6cgRpGeFWiopLmIkA3wG4ZO462iwURIRRDiZVF1+kvjPNWZnqB3GhoRRVCNHD+X8V
+w9bo4TmSNgN5b9tUgLGR7Tivjq6q/rcjnF1t+esSQH1jFaGkrFox40t7LaNbR/l7E4jZuimzreM
bDyqAHLhXeQqvK1UDqdH6Os2wJNm5W2kPa3sOejVhTh8a/3v72hvmqhfaoEBKbDLQ7boE71BlLIa
eK2zEiSVJd++U3uF7aMT6iwK3g1uEn+CzmGdw/xOhHRNk1ex8bkQqZnzKUvZz8SxHemcWVg7zfb2
35DCUrZGJHMjDEFP2QkZAAkrlOjtmUYI9vGwZLf5SiTr0fs8Q1vqzHRsEXbZFmVq9hIqYQJG2/Tj
OaPVQNV2i1LbCfUEZ9Ibw2R7CXLDDIjarISB1NPwstR08hJYgZt4bWxtuAChI3Ym8PZN7t+YTZUh
ftXO05M6DTsp2LoJ6V5v0ZQoXPyj3EMbAHz6E9g5qAvVDTdJl0aNqq4m39Nx1IGEy5e0O9c6zAex
vIMJ+Eatp8Z3CE2xxMUIIuLIM/8pW5a3zupuiGKOHSWVi+e+ACQr3JiznUZ5aIheT6uYYi/YetFP
UBzm/HXQeWDa27AEBLw4twVcFNTJWguj3Ne1hQuEuj0rqEspuXgl6DIyqPCuw0hWS83QuBmUvX/U
tlV8eZSbCQNDISutRn+kb98F6IP6WXZRJav8ZeSTvqCih8QWX66TFvH5O5g/2oBeWMHiSFV26DEy
KwR3kYoWiSjXnZKffGsD4UCj65QzIqzqzkzrp5WXLVNNFPLdYF076NRrjBuFNNTrbLh4pOwR9XRr
+NRLBaQFwshWlkQTOHrFsXa1PmaOU59wzZy1LQtrc15RJmZ0RAG1X8AnH6X8Orxn8v7RnWObWl7r
oLLRcjX2ona8wGmCZ9cKrOe5Cu7mXWsA8M6vBv7zyg6h09p7eMHm0x1lktzS0f6fC3cTIdIbzsAI
E4l19OPxQUCcwvYB7wFXgnk74iqUS3EVnDDurIuL3jWwZweDvkSaaD7aOYe/q7GgWIAB+jNuwVmO
pV/W//I4r2Lovs8nUT1H13J5dB0QBXBEWYr6tRFAG03xvx8CHjc6jLzsLtsotNmJc0L5e4CH3tpp
60gvqiSprch9N/vtjZ/UPD6EPtHCUq1hDKMrWfpg6DnYGXCRPkVAg1ot/xnT9x8mf7oa6izhmYrc
8vVn/9gA0Tl4QkKwIK2ZezCPaytwmBnAvUxUTE0QjktHBRtsy6cVeOBP64ytutRWCNM0Vpe6P8qf
MhhXWEd3GmNEJ4aGAan+p8Ko0qDAcmnS/YEYJ//yHHRVubM/TWCJS8iWxFz+AdzrfOmoiQalFkFh
Cc3rw9aIcEdisoE4l49WZU3Qa9bdJEKJhsR7KmXuDqqBoz0MELEF1meQKGQHW/Qqy7gzAvZ5Brn5
b8fGStiGvb8jdfCcSULnTJ6w685Yt/09FOuFbeCzKH7DcdDN8G7a63dISvvLddQrKVPhVGtuntyb
deqmUBLx6RdZwv9zRSeXqp9DGx8S4YaBUWJkcVUuF6kWZoThXsFp4Pvk0bo5UC6d93euZaMoTO6s
lupJs5PkQYe+8ubOM5eOKyp7cxpSqrhxb+hw9IhOaA1WZIjKCDWCD5SHs9+gf1u0tSTrpvCj70Fv
5zH3zqGxnUvZGNgxLz+RZun/ad4zg/qoq7af3GFgzsPq8003dRGKhWSuidl1xqPX254ysg1KYplM
VS9SECt/dz/3lKShrtL9wDLJBXjuPkd72kVAGY8//pFyx1+ZhQmuRRvD0tp7tv+3W5Ci3T1ekX0T
9LF7oT32O1XuYSD4fGSw+Enqhm7PcSa8prtYm1ZtoRuWjtXECcHf0NxNE+u4jQD98x3UVtpGA7jH
AT+RojSanNzr+V1nYNCxncQbN1ElhdFLvV+CfbWtGTy17LM2h50vJ81uYzGOtjaY4CrcqIfP7fhl
70UV/Lm2ayyMyM1Vk5zSfhTlhUEd3UcDWhkBS8ivGb2TJEdq5gpTtJ9Gg9ZHfbYuA918M2HsYjEk
IdPD+bdicE2GLJPbAkfjZHnu1v/94SdNDMdkeBVmtvyl8HdWtfgip8fwrs1wfnS5vPsSe/xEazFH
uJNnlpvwHyrwasGIOw8AnMeHlqY4lqLCX+D37avXl11tEgxEUddjI6j1Qjht8dfhILnyuh1do35F
JNfAPXfuXs6nlslUilH9tnQJusLqzH34DanskejOovkw1ZTCAyDdWo4Hm7TqRmo77gYuBaV/bIrV
gDPsYfuoBdWAHEmkbblBgqL+a0GNaPSDlzM1N3HCbM3B9+3VpILfA0IQsbL7Ss728eBmOre4okW7
nZ4zh3edRscktdDZNQiu5NAL8zXEUAyn60rcYd1VR1pSot5yo+2t+J4qB2mbBL9EJLD/qixIVeS6
+Fw5kPvuXSMShO1DIWyaW6li8tr6VqioIenf6R7MM1mJz3krhepq6q+WLF27/qbeS/86cdb3AnKN
wZPHEb9t0EO8fXsLLGt69ohWaoqyHg0PIaZF9UEPin64JMqlck4URuQ3lzCGnbehVQPHABuAn3Mm
wefNv9euttfALV28hsWJqdcOmspG4Z1kHWHmFHMP+9PwGcSECjq3GDAhimvpt3BPPrr7zdUNkTuZ
rAG3g1D5OqRa6H1uVilwqDNSv1ToEvxRhUjuBT6+pNaiYiUO5QIcGWlKpZdbgFgEDrH6lcUA0ywe
jBktHEOUUe0yrmdAF9ch7CObIZ6zvyZt3HBC5o8qQbiW58XfGTnOa073wK2YsZYY+n1h/buUCxx/
SLh5bYd5HBv13zeR5kDW7a2gtxtB4tXtYOPTbv8KgkDNl6/VkS93TLIMsqWFQKjiHnH64Y23uU3j
TmDYCpoLGQFzECktvQvknfRQZIQxzb5oumV0JKkWemrKIEV5T0h/3GsWBoGm4onwasoNP4XgxgAl
AqdAamxQo6JGfw/JCF30EdNSlt9mb++ZvzKCa2pUEb484sioeoM5ZPiModWbqsGrQ+Al4a2mGNM7
gPjyYyprx9yF9a+01aeviKurMHnEmJ9jVTJTQyzzDgMY1k8RFBfjYQUL+6a7BK0Z4YsbWD+jQTPz
StIExNSjkI2iaBpWW9bnRHpT4EW4pB+Mxt4IWv+/juRPpZP64y4zst82ZOUvPgU1pdoUa+Qfw2Ha
4j+o1LADn+BND1Yc10W2xXg673jeHTMftr+YQnRAIaSmlHHM7hsnEVorYnl5z2dou4zlDpbhTrOS
MpNyOEql2CmCtLGo0Iy9gvg6JgmVJc4yOpSRd9lC1UNrA1t3a0ZvTP83Y1W6H2H28h+pBuGx/X+2
GtQ3d9wtDsA45CJJ2CM32i5x0U0ThcKf6naJOV4vZjE2feKXiYeSy4Gz1nm+aLLFm3THb5WPJYkm
pFGFl3rPKXJk4WkJn8kS0B25ON00P2j+B2luWjIuxuh+kLSYNpWE7DTDjvAw1JPcqjLzc9pWkEaj
wNydep/7YBMNrWuu8a91+H7h+qxhTt1rl8B9wUPDupw0MFptFHI/BzoB/fyd92PMwfQ8V76LU7o6
vneZ8r51emM7XPcMx9ui4FlKIiEZ3aa4a4v6IHXtfAEiIR3bL4BDr0spBE+MZN2UNfVrXLLe4oOn
4QZG8d/2rIYkFRRsmbsvLLBwV5skh/fys8KOU/YOM1LUAcBRcM3DyI2uuELEhLLpLi6qkzM7Zn8u
dsytVsxvIYRZ7cauZ5omAdtPtgGxkmmRqyUJPbOqgwKnGAjhKBLntFabHUdHqC2VPIzFTIYouXAW
IgwjGwohz+juxgKqimkLOTXkmQrcckFrDN/8czXAyYPKy2q7TmkaWIyou4ltW99gy+Uqd/XQcsDV
1DCJWNpVsxGlxFq2WfFWAtaHmVvlK704kWCTnNHodRXYmn/Q3ZtN7YS2eyfJz8/FicLOrcYxyVzi
9X/Mu4TjZAFxWsePqQE/TNeQsp410KLf46tl215pS7k+WaagDoU/cq90st/pMOlKr+el1LQoM0ll
mPnxGNw+ZkBBmcKOnRkoOJI7Oav+hjew5AF8osH/LT3tUPmEK/rDtGZXgSVvAXM1ij+C9DtRkXIz
RE6pLjBkECW1FGV0GbwfTZKJk0uNGId4E1iUZ+mI01p+EO5kleve1QWdoZCaeklGw/EpO1Bm+g0R
dqiIuH/dJExuyHLyRkXMzaLfCsUh1nml9bMBKgYvdQ0m1/XPXDtAMUQdI9C+pVwy84b/GYl+eDPF
EYeXvRQp9+hqkWJf/+lwxlfz9QZ6UcttXRI/navonV2OkJbVNLID/LNC6rbTHdTgZ1jHoA+X3l40
YumEKGyd7g1DsrrgcOPdmOOOX/1/TL3tgUq5iPl2oeMjRENz7/mEO5E04CrBwMwE8WXu9+bBcNZH
6AUwPZ8MN7lFuLeOmMhunMniWbmu7fvHgioAu1Hx7Xcam6tZYmjt2g12bJY4JbZ7Nbl7CnR2jPVh
X/t5ONlTGWpVzglH9Vl8rpYW78W+wAaehQBKLsaqXdnp09ANCNZe+NPZvU5/jF74w7HN1dlfdUcw
PMOWwsCtDzumtVgtsJYM7rE0cmCvden3mX9d65xJeXzPh+UaFXk3St1IaduYuoal+n0yPedORxce
szRqYNwyx8FeyQyAsx0sDNAy8eUsEyeHid+1Q4dEAah0Zl16/+iIPxMINatVPgwMBwxkxTe96snq
XU9dNN0wmgsSxGow0Zx8RIIg+5Iv1pp8HyBiDXDdw8cOOFOit4tRT9uXqJVDZ/xDLx6VH1Ij4ZIw
tnOpXB+p2xrUboD36R0OdzxFrAjXz3JxtQ+qMKy0vA+4eEsBPddaxjrVOwHqeHEk7jJqBDd5EqD5
bDxsUYUecEoj9igtPeZMPKL8hBs3Z3YxWJ6RjKA9NP48c0CBr6yijzd+WB5pk5FkyOCD2gChD5yd
xJ6fqc97+NaPSAbo+w9k7bdXBL/RK/efJAApz0tdL7Vf+JijFroSh3KdtZgFerPwmKQl5ME3M7kl
MtQKR7z04ZWOzOQtDPIgLdHHtYSR4gh88ZgnUBd34oasKDShu4VYZcLb/NebdYe+aetH9JC5PkJa
FIsiKHNnDVUXpoAFLCVkv0gfXrsITXs5P3ZYSf3pqVxcX8JCtj20ZpwaTnd3CaLzcC5hEvny4A1s
kqZfPBOGBL5oq6gbiSgyNs5sb6BN4urdh9u+CRuy4qOlHEpQBccBkV6N51bpsGtBJeZI7ll4wOJd
q01Ox/gJ7/VS+NS0CmeOlYPEr9V2zeIHK0FGHjzHtQ1ezGfQ+PnxNhnN7pEW69ME2bLzXePyqQBK
lN5+abnMXJDCkYb+bhGr1cC1Vj0FTl8m0/Qi+7QSWYNgD1DYm0Yk168VIgGjiDNFTkLwScvy4y3F
bBk2+o2TtzzAEdyqVZuf4iFtvWpKIuNsbax6+qFDDgwNA1bJ5KMjReV3r5Vm4IReiu+Fgb7MU/gn
OjJI/G/y0tftl9XhUMWl+S25l6u8Yp7EyyHN2X0liQ1R0U+8ueja0KaXui/lnyAo2LJLfomYGsbO
JjRS5cx4USGbfw4VxwoC6ZfjqzKYFZaYTCOztly+ECgQzQk8ObaHIgKnXUWNeagIn67KZNtXmaLr
ZuMlrOiBkty65ZH3+xotBjflJhFho1yGZr8m70PaiMkxhUS5HLqxShKMYhAdds5ugPdBr6908uKE
Nijrh6wj/xRi5VB+z3bU6c0ROCE2U21nFrNHUrXCXU88n12o2+QAzX7lt0gbwSHDPOrNPxJGCtQ2
+dstwrsB7DbjmocwsCw1SQVMXazoE+cdT8V8i614QqTiYBWzl3RHgfLm7MsFkJrFpNnjHytHlS0v
69dajL1z/LSHl5zzRLey7Z/hFvYFc7A+vQ6zmxD9tRZ1xNSTZEO5TvRvnwsul4nljfDcixfJdocO
NRPpuq0N5VgTDJjPYeZ+o/KwmeNTy3rghW0PD6yh1YCUhMMZDY55/iwErx1VLyLDJqc4vLYf00Nr
y4HjJSdCxsoQ2aBgp1kxYk0ZZUb6E/PskcSuVcfLZIHFuxgUi4zPSnDfs8X/DcIXTzMbA9v2MdfL
YIiplz5o48WCp5d4imrfNhn7sPdILLuuoJelo+xtxfHtgLU1ePKpTQtoOmUDAhSo0tRUlH+e/0RQ
3pAZpO3rtxEEy7gdcIvGkFngLQ9FDKr1SWpXGv0maUuEC6XypuEZbtheEyltd/NiREEkpdt/AhPx
R/dYcFf2rbZ/bpbnFEuIoOBGVHfhZ/2TD7kLqwuAyTeWKQRM/h7e37UqYyho0CqIC/wd2SUVSMQd
Y27GTFIJ/YqSG9Rwg0u7utNV4ZcruoY2eBpEDoJZJIO6dQtCA0QZ0+FT11u47C7Jn682InvPCqYN
PnQRJNrZwgPU/5AeXr4spXCAER0t3SXyWhJNDVJWUNUqlRHOXs1YnpUz6DnTStnCVQa8j/N0eT5s
r0KY4MwaQrWFVE2Aj1F2Jpn9iusaVUeH20wGmFgPeMAM6Am4+gXH3qW1mT90nNiVW290yRtAmZTA
Rkv9LCgnL8DkIwYGHTodBIJknKPPA10eRDATP8je6TItwd39tVOJytldFwybbGcxSdDR7ci7OJtd
rXr6tWG2yyqAxNKOmVFRn9H85FyGTTgxCn28CKZp/MPXF9/Cpgx2c1ZBwLxngUO2drYEWz8vqm4F
venNw3ShbSx+879gc77kt4o0raIpu1+GzCwj/wnBteMt6oP0GIooO+L08zx8Cb5VlpPe2CI+NEjt
e/WBS8Za/26AcobX5HCxbQBLLAYnX2H/wApHzMlRWBWeft1503CXjqQJsnxvKA2RjzYXP2rassh0
HZ0b5yKRYCLGwSM8vSpzQMCpi4BOG6qlP6Gl2dvoG9RiLd2AqY50YMMqGIFB25qjLWcXQMRGQVO/
Bf37friJzsTjwhvgbO2YeNi4edPy2F6EFO05lOk3J4S4fGsRGIoERdSDW7An+hxj5SxK3xG17pTM
xbW3I30ByutPRLef23ncQckOXtgaroP/ytrRh9wJXtaSeOzntOldvMgK4BSqIbeFWyE2OLwUXKuq
V8Xq+egpx99MObsDVJV2CAUCcj9+U25ZpJdQpAEu9fbsMzL9hnxuNB7PxOM6t5fkxvMtHsoT4BHv
ptMfZuzP+6824KeRV2cfmQhZlCfu1eGCbBzZhYmt9buWxe4mhSYea+LRCywlCYX+P/GnPxVeWkdE
tL4yBhyJUxQ1KO3ycQAqex4TcOjj7X8IZ6/0orEJVvIh3g8w4pZiDAJQKAdtV0Si/7pqqLKKlVvn
PybwXEiKiT/7u7H3itC4JrqIUdhQBFqGXcs9bMP9evCcE14rrMzFGGxpIBjaaUJlg2N5ELE8153I
iCGESYOKXuCv+mL4rz4EYI/UZuYKyZXrCwaZ4sB3gKsAS5MtgOGFjfZAa4WYYkeHILcPx1z9rF9o
gi4yyH4T3Z6HIeaKsxhfqZiDDwsxj8Fph8ffWIttHAOD15rCmh5Y8Y5/L8XChB4rpJymlhuNqBKT
OZ91BqMM1edgWPcSnRD+08aYJ++DvTPcVtiWqb4/weLiCUZNM7FV9MPuZUQ6YDpffGoB8Z/wMeu7
PpYrJRnfDYd6TuUG0T8An2uy5uyRd0oPL5/oVl7YKYkRSpEk86epO9IEEYCz8/bKD1hvSFmFTOZq
RnI/HyPpY0c5045X/HW1wRKC+zK3zykEHFBVGAlcFt1yftLpdgBaxzZazY3NfeznNJyHD4wAiea1
f02QERpvfnlHUWxGHjV+gsc9E1XRh7/snGB2lOqMoOoCTl9Mif/fbFBWxg8fu/RtuUUeUoSdnOrQ
i2pFIWObmNkjxVURAYNo6qOTGqKKLIxnpicyX4hhYKxXVZkOo6h51oknIEdRBF5oxFS8vUMBfguR
Fwjsts1NsPOOpE+3WakF+Ss5anp+gGRHImEZtc0hII6tJ27oKWP+CYgenfpbrHhHs34lve6xNHFi
Fx6sh94zkEUerKxWCbokHEMBVq1FLM/LsuYLjSGd401N1Z/+y4uPCyS9badVOYiBM4213Dl2nyl6
JPuQCCmUqzC/q45THQ+vmoUFtjD4uyIuVqJJ0KzWoKvql9KGuTgOipI6icIWDXgvXiupL4QLxLiI
Lq9pvqkWIguWPdDhpfBhwGySJxDpDIhE1MMpArG7g3y2/5LDCUMF6fcyQ9dqzttRa/QQMIJhJeTa
uTnJkZPkhAfdFl13Vx2Zm73Vf579PBQ7x6MEpseUb3fKdgPFMdg+WatQ+A4AwsHwUQYcLccF18Lr
dGvRKQ9wIcsiEJzpFPl5oGT4t1kdQr0v15AEUL1uyVsbKmKgrwDx2cjWWPfqAv+O+wmN7YdiazKW
FL/p/Wwy9EqQNXmq+M8L6Na+5SFKhIwxo6HbFk4ax2Ma7JzalTIh77RQaD4JP/p86IwDRc7DqNnr
7ccJYwd1TJONYDUKIET6WP2t7PNaV46gtPSFfr/DL/XuJcf36ZZTvDmmRGbzGfnPA8Msw/s7zNZg
4WIoLTeVkZ+VSd3RQhwhUQ/jG53b9/5qrzUlJr4PTlJLhyrLQSoEYxBLEM8O7ISzSVsGNIapcuTc
6lcipE9X+sgoLaHV3Oyol097H6o2h1GeDRtqIRl5OWW+lIjRk4kzhPQJRhahDs2x+h1iIwaghNPF
Tb6ONFN1SZHXlB0KEu/EfrScvI7KnN8rTuliy8jSCktNwdeYzCGI95Sl9mGi6m/RWH7BMRazPyl8
nlbj5Cx1OgAD8u2UCCW2ppWVGZHv70hY/lStATgveeWn1qt1Mm7Z8O6sMaF/1IDUn81ePGVlL1Gu
Xoaqmq+diJw6qPLpXNg9AA7WU7p8gCYYGM5VxNQRdutrohWtZzATHQx4gR0TwpR5KaDb+/dh31wi
M4JTUv0u4UUWA/BX7l0CUHsko2/3K9Z5wYE6MKQcPot9H1h0PXO/Oel4Kjto7AJZFNCYH6gK4PRN
UQa9a+6HXsaDxRnyTVxdkUF5JyjqjyQbvxveAtYrhz8kKf1xOGAde6yIutHjk1diiznigjPruuPF
NNTfFcwQskx0Zc1nD4tKUrlqM9E2M6fFsT5T3sKSIkAHB8xIMglwmz4UdcxOiGNwo0kRk7hNFCaC
vUxuaHZNeBC9OWO2PpsCypfVgIOF8eL1BYQVlHhWgc9s6FRgtmUiHfNQZ7Ewjz5OlwjDJCtVL8MH
d+dlilL5CJWQW3DxWIcr5bnZ9LZyWEmEt+8Ef4Y424/7QuyqlOj2UulDrcpCk6NWttb87YW5fb50
MHe5IHUJdoZ087V/Z5gwYlPgHQhPukzOHxlQFDs/ZaQzuY3i54fXIO1vP9SWZjVodbzopGxkAQTz
JDYmYYuyDSsPygb+mP7xOc+abYqiHVu2oMWmPRGG4mhnYO9Ddx2ayQUyrew13momw+9Fhq0ABuHb
Eg2kICONB1qXYgRWULoK1iguSW2Jqwlub4Zfmjsn4Fry7kbs8ADkgQ+OxHDXBpJnDVYISM/jTka9
kzC2dWkhZtv1HFCBFzO5pPTU/P2s/CqW5CBIttIcJnR1dN+7mg4nUHrlHfWxrtDtwB1OgPIfCgb3
ol2gjpRjzi+i+PltN9xa5ETnICoprC0eXkh8/A/5VvOY+xWRXuSMXDZ5ymC55Wy6eoJ5v8n0mRCC
hNDPjPdYSZAFoMiXRo8aM97OASnRf39iq00NhbXBbxb3psVtrWmFurUBqM4Yih8uqK1gI8FXFS/D
97uEqDtmoofJEbt+m7Jom6RoUc1JrqYWKGSiltt4HqmhXvO34KkK1h9bAzX57/yfezqJfeGw8Yqx
QaZwbcL1itsCNkxUy8Vkp8wgTTs61GXzhgA1aPdpFR21WcjJmoGb/qCZpTyj5UJXJqwIm627W9RJ
4uSMfqSvXmyWTVTm8EJ5DUFBLPBcINGOUWEkGkvzLZUuCluL0kzCK9dUdihP9XsJI1RR/Nwyrdf6
ob/F4eACrjTRVEQJrsfQ/4r6iVgWpRBTQDoogSMdZ1/QhT/E5zGf9gZEqOlujCokU5V28WyiOGyb
41/imHchfxe8FGJa8Hl5eusUoKdolf1FcfmJxdaVFqJhjypJFvQRn2ITjap2gWWVMc7OKromfZcr
ZPTkNA0Y+9MPsW6tRQRya8qrRJ2Fmt0erekezkeV6jLmpOBdMAb66aVNaQd78kwfYVL4C4n8md7J
3ck+xRXAkYRq7YF28V4h0Hpg0WhWtX4kCBhVuWtxXXSkICRSC0rqrF68HGddQ8fqHSgZU6634oWL
+6IL8SzFFjXuMd2Z503TO6T64QqlmHd5k9DIsD0haWT58KAZAG68vhDU6B7aq8niiL2gxxps/AAJ
jrR1VzoxYyXy21S6j4CJMj8Bdo9iBDw3YF/jwPr3wMCfa2c/FnapCRkEBMX/dilU8nLGX+ubQazL
QVcNgxoUCtkvnBX1kiSR9OYt/esnQpwpSEERlO7N6PuPPYLOXMdVr62jbb4bgaNisb+SQqiVTq7C
x8Pd+dWwAROaSoBLsbzVNKD+cTQVYBb869msdB2Z29K9JJ/6o8hrp2LUbti56FJSN4eXEjES+QC+
PR2Rrs/95HCy0iMp7JPbwerBIoSZL9iMO71M9q7LhAkpTxketSe0THiTWmmyjK9A0YTV5AEGMf0j
p1Klk1fWn/CYovLtHaQl16JIjZhWIYWY505iDwlU/MJ4sncUtBvo/rXF9DvEAH3XRU1VKCbzXSpp
ydz3/mqU/q5JR+6nG7V77MMW/7LO5fZPi/UFQJ6uvCTMQlcnE399fuehs8aEMtyH8kqlF2PNsExA
ocQ059vPDYF/0CWM/b7fBpB9n76igY9BHsWVyZmt2okoSnFlK1g5AWvlOaqMPGW2sLtbpk7T6crm
6ZPfZF1fRIWwNavc0FyIejPCl0isZVkRu0y+NxR/d4vN9hzbBD37zK46bnXD3tknao/XLVP3MAAQ
y0Kw+t3BPhYftEhMthRAaWkZqXVb4iZbHHa8X0K6D310u4N7AhKLnoRwSS4n6NfDARClE1d6R+0e
kJrgtIOrikPVsCRtNMp55ye3lnbdN4VjRtPslh/s3L+deTVozMivSdUYPKFuF0Vbcnc3SQxIgNrV
ACTVUsF2O+3Dq3D215eKSLtewI+0KQr+gosBqqprCJlxJhkM4+2R6MLVKLfELC9Y6bxJOznLFmVx
rldgp0E871ef2Ds9KIQt3t2l3nXCFDV+OBtM63F0eJOOK6qKQRySITGYIWyBER7IfYU1hOwwC6bI
wNQRax7k1tSLyQzxOrsDfIDZM0IkuUTUXFgR0qGfnzeHVjXT1OESqHIQdb3GTMmEh/wxwO/GLkHG
+XI5omzoB9Bb07SNblLS/Sew4aIzcqMJrdhwt1lZXmx3gPHx2pj+nItOAIPgAU5abcPU/WCrFj63
1uIU46wNHoqnKUdF/lPVe919CK2mHcL3ZOHnwrBjo5oagP4DqFwCaAz+rFkY7MCfiBfBGI2dmrIi
m9qnA4M5dXOw+W98sVkL02gDwJjWQS7ul7jvblLg/1NxrOyqqcBhLzUBA7ga3yFQjNlZSkCkDqzx
wT05MOSyPRKPf29Imo8Lvf1dHbfu8CzI4T1pqeqgzt83swD6CBfl1XPOHj6eMmjHsfzspx+IiZAQ
+tLTxtSEPX+iH9XSAg4M9F9bNcyo+z/Zwp43uH5tTpdvEOqxEsnvwYQCl59kDJ3lnFkWCr/HdzhZ
InObTd0hdoCZUzQiWN0H8kst6O/rPqoFyiqkx+4g7okK4KuG889OFeqTHYhp2VhpwrLEzc3z+Kez
Cmp4jGJ/lbR6D2C2/98MZFlHKRywodv7BjZQiP3visauIpLRIVyJcMaEaoKiqDOwloN0Pwd95NQ9
F7pxr4jSNhdtUHxqRWPFNYWZ1EQ2+MZhFd0+v/ux4pa8HQJ4NAYRdUn5gfs0FDQC4oluJOCrCO6s
hMLFt8xvBMiMPwBXZby8VsJjDN0ki9e8ZfQ2dm0aVPI0XH0LAt5GD33s9oyEcNtMmyvmhlFUGath
7OEuTptQXZ6kQtFFVo10IbzsQv/cHbXdIZe+LLs/rc+5A4hGL2eyHlRZjJ287x7Kjrj0f8qMKYO4
AUm33j24+Sq0b6woD5sOnmS0MEwy1fXCuOqy1fiMbRetnmyxW8kZW60jl05KPFrMVB9VhodywIsf
FKOKAlFjt28zFPYvn5YLzVtJP8ReqCkza/h2CZ2JX14mmf1yIzOnylLX23sptFQ4iHZ45E7cxoRQ
FwZ8NHit/EwJKr5TgEUxfeiMSxO9Wh2IeDacZjwg1mIkN34OxJejBJITy6AMM1Jq9IbtFYwIkFMH
CkJhk8mlr4WVJvD7gGCM3eRn92ptjHc3Ejspm7Ylx7eY1b8zicYsKUZvJ4XjccSTerY3Um13OATH
6+JTz4tNrx+YKO6qwnpk+S8vijoh1p3qTGtpIRQflY7+sru2Gw/hhnqn+GPbj6w+9fvRGH2V+3fa
Bx8sOeNydDguohVTA2/HOpkRwFHPFL+ZP0ozfLs1jddsqGpnSn0uTlezGJ8ZFPQ+frnaJK2opmXQ
hr8ToxY9OH2iJqVdiP27TCxosEBKgwGu/ajbETEBnWZrzVaFbfVVAGiFamt6PgKeNMUQrXabor8d
DrcmGsS20ncy0ksQubh6aiGUASCBkjyf2hBEKv637CyK8puNGt9RJe1Nhad7FFmkkeq+DBS9IdTF
cNSpvdwJYhA3oaed6+3P/ImJHtSNT7g2HoDlkfboIfM355pIiTCLkqP8DV3zprA7Je8etkWSBXLw
0TN57asV+76KObwBBMFaoNFOCXAYl/Vv+ouy/G4QDyJpL+H4iYatEVLyglBSK1CIRpGUFDfJLGbk
AmW/LwUr45vuiYhR4QdUof+r9uN/p9mo+oombWay1dS7EK2WrX5VvaCwT/T7dEKMsI/jYYgoN7W5
sDqMyQEJJp5ykq86vG/yOX9lQ0hLIzJWXfZ+YiGcWKLEgIpcG1JdPRh9SAuMBueQIw7lhWDDHaSm
gqXyIm6+c8pqKtg7olOR6Ov0OQ2bKQyPeaYQMkM+H8bxO/ulpfLwZurcOWq2U+ex58tkSmVRacye
CAs0P4ery34NTHVE7KVSCS7PP4KT/GfhBCjw+koedAud+eTowhqRnGlwH4ZzUm7CRxljVZcSEkT+
p85b/gCz2E2SIRPt1avjjZCu/hg2oZFtWjrADMVVjWryc47+a+ZaLjG3qIo1WuhgRVGKYxdpxn5N
sAW4iWfLwYEHSWC/cPcQeM+TgIqT7s0x0g/Q2F5dxwJtaR4sDAnfJCezagOCOAj4ihi/IUdytgp/
Fs/JR2COSpaHm0uSkR3DdGrwwU6kJU6yYEfsNtJ/PL29bUIKFgFj3wPd2ImJ9cmFZMXWIP/Kht4m
Y9s2yiAIGYb3sBe5krzqoDiknUG6y/Abkcy9zK77U2dn7yztKQ4S+C6k5XMPhiVvF5mJRrSxYwxU
qSd0QEvIiMMV6HI2dWpXgdJz7hLLK9DUW04y4U6dBlRXo2+j41LorskY9Qwk8BHShiuIo2aD1Xo7
6GtRvwXT1y1GMJDFivRdMe5n7N7CxEYRr+2Y17ZlhvhcfY0PMcUCimvZt+fnRYK3s1/94m3ymBGG
/blxZbYXwv/JHMiwQA8meDK293Jq/AcPhNG/PSg8ubYnjUZii+OcMSenNjummbYELKyfc6YDeX1T
S44thX1wfeXWmkxFbP+bzbdDJN0s69ZI8UgqHpSXzNFfMafM+y8WooyNxJXkSQBZOK/jZrlHVL+k
J6UxHXUEk5hSlDT6xnQrTcF2GtP6jisAVX8nrTInrK4O0q1cCd7miNWq6c/AkEt699R6jJ2lFd/d
pBO+yF/o23l4DzMxUZpubrAV3VcGLlEM2MZn6YqsxfGHlF/0HrETfxgDXWk57vIZmJD0PlJJ2IHB
p7LluHq6fD51uj10wBH6YMKcQxYdtBx72NXirzN1o0rU3FOCEacFmo3RBAjXYTWokUMkfcPoG6Uv
mQ3LU54PbuBhwC8Mkc/ATPU6z1Oof2oGkPv5sj3ZAdp8s3toE5lVeF24994Y25xaQl9TwxzoBlw+
2moGLzN9ekiWg6M5+XWEW3/LZnyMWl70Gz5VGMrS/E3WuUTfDW0DCNrQJgRHGHa21FRAcpJLv7PP
KVL0lY9hRG7xV+5SFnZDu0SnFN+fOZ6ZaxT8L7l2+W/eXMNM+ts2xk3YnBjtJ4MDtlN3JrrARHrv
AFi/QHPR9bmYzUoX/a23/FmlID6heaCKmsMrYfet/8Rsn8lSgWYdjRvp0KIHWsdXa3AYGEUt4e6h
Te/vUAeY7OH9eEvy13DJz+/85Vn7YJxjvfwGlshSyswlcIKo7OrVYDzylR/ldwCVUEc7q+sNouwS
WaC67O5VvcbCZGYBatU9OTjyqcCAhsNkdyBwtfBMwV5/ltlw1LbL6014E9MPzWnxVxwRVAVqeH1z
7Km5Ndbf6epK/X+IC5CFXb34DJoS0X0imvCjywdo5AsFO4g1r86boNU15acSqFeOwDk/c6YhHG0H
O/5vmwUG6i+iCG14YDINAMSLz6waPddaPaDj7X0L7UJ8LlSPBQsXlLAJ6Cr1o//PpuYIz0UqvOxu
oI2R305jWXQU8tfZ7ojmBTizHg+STznqgf/buWHjUIj4eC9OgrCQfzfGvjqzeUf9ypmeN0j35+KC
Y2FxlDHtHH9+jfE84dzizMHF/PQKSWcL42L+Apba5luje22J+lHHoF3rFmNEKuY57HGpKNwDaUZb
RtdC+A2zSVUFMUAGZIA2xFk+TRwIq/dobarBMFAg7i2jbpYrttvnCGZebVWE/U2vlEtKCaqXnIc7
fiEtrrI7i3n7XU2oi7muJrvSy/rYbYi4JUDzzwf2SjsV4iH6uPEgmp515MOrj4940Y500BEjVU61
zIY5q0KnWSbx5bQZJ2lmOwtIorW1bOtAW0W9RYgayD5LQOKubg8COKvZz7XxSQWsB5eYnjZT7bEe
BBZthe/XAfJO5XPtMlA5jZNcRBWDqRjOKxlEJ3atixRYsHvQdaUv5HXzK+/5CeKuI4qjNbiuF6gr
ULUju8V1s3epGrg7xYHcpYlL7HYmWm1WnGjASL2I/qireal5cS1aGgmMFT+l5ksgom+ujh1VYCe6
Z6SD7XW0+46/xbZLgtd8Nj7bO/YIjhie2vUc+//ygr3LzEDGHcXWgke7cRy7l7gDNzrxyhYcWXF1
JaoIWAn2vZDEG3MgromjVXA7Wq6YAmwr5dgJ6Su/ottWqffdpqB6IBCvl+zegjSyzoWK+pzCCEkE
xt/9cZdV1Pn6NvcYny4i3HuIUIANB2bExEhwpf7wovD5FCkPmhH6XXYWLTnjfc5+PRq+plWfv/rV
vRs4AhnXBrt2l3AB3APK0Gj0zmkkPRgF8OzyB9JsCRKLaUNhIJWTFv8DNJRy3GIPzJpBH/kIBKcP
AnN+RGVeEH/56DiLaXy49oUvut5aPcqreS4lcQZAN9GzutvmFmmAzPn6vTXrKl3+D59J9krCxWz1
OHq3Gb7RzZo7od8oCM6zTKo+ukD//55GDFTZ9ZJEhxL/W5LN2p/0Ubk3mJxkYfxmGTbpgdcPMccu
CtjndSzJznYWkQTZMnem8W2bf8D7RHK6tEPNd3pQ9xgaa0+EcL0au/jE5XAdJ2iYYws+gytmElRL
2jrWjdZJiGI8E/sTojJu8csX6GiaZnrlbR5XAhtOzMNi8BchuieDT72M0oHN3RGlIk8EmEp16024
sZuS1BbyT/91YMZ/7oisOWNioP8RGDG/tzW5EOJ8n93uVrAs3RMT4XboZB/Lc+AyWOx5yl/FzfSP
ZgmE+XMOVLyzKjVhuhNfTeTyrLnGz0m69+lskwWEdQJ+qdc2a8aISZIEfzlb2jp4ZK/4pJY/q/IB
F7Gs4tnCsIZ06mdH9HlnpQwALefp6qBeUbHBsqjPW4o6yshx1BeUhRizzH2B1LU9wmcWNn/cMWAi
TtEWOBLH5ALseoQDWAsyyp/bxS4Xv8h74p4KveYNrYzFWUz1eEaMaS7wCqVVhqlzGztqDahzFMD1
wO1qQpabQmhlrf8gkPssOzE8ir5lVhDDskKjmA/9bxncuvZ4xdnCUeVHwWQxAq+5B5Yi2Casm4RF
p/6+nNBGOnz6yYJCq8hY8fOHBA+utGtUeTCoqxsqPE9ZzICEzZDmg1IORE7dilg4YtB+2+Ly7M4y
4LKbMevJyCnAHsLg43B2A8MQDltjTYjPz7Z3JYZ768Dcd/Uob/ZulGkFhtVJmZZ3WF0qbuHZaEHs
qiKO872vTa/xYMtNcKzPkIQlLwgKup7XBdE24JJNwHNMqE65+0WGrsfFeVluiV8uyJv5lKK1s8LW
6LAZ5M8N2UDMFZhw6ZVfyTImFNbIYwdWI2MT4d3vfjavp64e4CqtxJvF+ue52kC9dkzOeSE++U2n
EgRyGkgoQ+jLtDl7PyMC7W3JzW7LVwwYdSm3kQc5ihgoTj7U44zdRG5S+G4F7rFETVTl64bti2vB
j5UXz350TUKOsYQSXU40ksJ0htcNLbth2Xe7ITetcv85rZzrgyjm47QBcbhRqzxN2cF3vGq/r6gy
8ld6/nmgCD8zy8qllgLNXwcDwq2CNkNqdZFBQcPxdh3+cuEKJrHmV5VxNY4knwdF5I6MVGmJlssk
ZCfa2Nc8FFvPyJQxz2nDuVS3e9fXdrVlEeizdcap+eaQxsnU0T5LTXjqNqnI1i3wq+/MMx+syMcK
DWgoCiaOySTq9qH6zE4rw9/fsrXa8rfERoxY8HsiV4GpLA7qmAmPY/9Q6KC8gLiAunymvk4EjGVC
CXDsAiZK4tLBrN7M0qx4Ngg1OXXcKqVTtImXjl2dKn0tCOg+vukOTpl7cFQXx7y5aEbvuiq2+FrM
eGmdjHjD5RD8QWvIr9PjneOkaMeWKCk1FJez3TZ7NevG/HE9+8+fDGmT5rK7HPuCjYW0G8lytKd/
E0Cb8eUO91YwbFvBGEEFpfA0hVnhNNOSziATEls7Kp8zoHZ0ZLx7226vLYxiUCfTvxfN3ppC1O4Z
luFuPwy82rICKUX6lV2z5pqjTjPr0VVyPxmTCHDf+ptqkgRj3czWv4cfFgAoObwSUpcAlxdE3OSO
4k5GTDQxjoXhqmAXoOshJnMrPjsP7jME1q76akRF/BIvq7l2bamoBOIa987Fe/5jf7pWbqkyullY
QZ49A1E/P6S+sYedG3Ka40AokuRpCWQ7gjJtKrq7M39S9XVuYfNTPC95N+xV5DTNfKgIUZ8MjZzg
/IDbm6KdlHNXcUbG8JhKzOgaucGBA3UUk722+M/zbQNQiDnWi919YwemPXt6yHEuLFpLIU0BFPKz
IogzwWWufYr/6JKIDnehAR4bgPYKbJ0rgJZTdkJ208X+/YNSbtZyb7OUh7YjX/FswLB3U666Kzuk
BuM5RE4aSuf6puBV2/p5GWQ2D4S9/jQh7vR8QD+/Kmb0NdncLqarno6/lQtqcduIzy5RNliLOB6K
gcN5QjedVfbqEPyksvvrK1Cn9INaN4AaWcz4INEvOXsz7P82nN2BFwUyTxqjFkRwU+FvNGs8W0FA
ipakId7qjiTeLE4knpdXksc2ugwt2Bcjfz4NLUtGsI0m7VVlTB4XlGs1WIrW4zqXG3elb8Ep8WF6
m/6RIHtz/ZtgrLxVFcXNQBu4ZPTMQnoZ4ovEZjCnYPen3yJAYLLEZSLNJtUxdErLGsgIwMi4er+7
NRWGACtB2vHqwf9q0SKD7YR4RHtU0HAzKFi0UOOMEPHOPOop6URqcDcHAXVEWzN+YG+PWEes21G9
MlRSjEr8+xFNag1qDfPK0Q6Pbb2w3r5rQ7EXMHZfJXghVzRzlJcd33wXsc5PyrPS0M0bJwCytR/F
dRwnFs6/x6YupFa/RQFURwpcA0QE4JOuNqlzOQRrRlp/E+3g++S5C5s6am+idNjDnvsOzf0jZjBg
iSUKrt0lfT9h48yHeSPq4u2HtNuI82WgtL5u2USImEYpTb0PdAANOu0XMdMb8NG7qgaMOvq0en9S
Xtj/QbIDAQHfbPaf4fc6SbC5pKIzweSRmZ7o65ITpvY2JFQvLo8VQ5nqR2aluVzZIhNsFXOIa2/S
8KgD3TeUWXm9rIQmsPbua6R/Wer8uCQrf3S94yZAfFlfEz1yfY6ksDSky+TEHNrlF5afR/r21PrL
Ecse3SXZaxXf/dxVv4/xC2MYWXuxo9GNYJk+YApcbRy2wKF7uTXgtFiWToSSdGeN72GBgQtU34gQ
akxM3JragtWA1O6y8eYIVbPC+cLI4diT61dXFh8kmyiZSsYKSHCGJY21UgX+74JZyGf5IoQ++mk/
ByxR5DbpriG2MuzbCcAljTRfooQWrgttZAlw8FVZGZNer5I09tRb7eNXgDcicz9Quwty/VEQ3sQR
i4ZJ7cXQfr3RsylOw5aSAK3elNTi1EAOj/rujNSJF0DjnLnVerpF7cTtSBJVO5voVtWrcFlWNMjV
aIusIxQ0dp+9cAjT79sXGkEe5dQIANEmcmAbCrcAQCA0tjjpE8AqnFF8cm3cyRnwWBqfGS+LgguC
rYUM5qiDLyVzdm1436V1mWT0cs63U6LJKzWguKK8HNIevA4hcSl10Hke+v+kSFX+EpgZXYQoK/a5
IVfZKUzQSkBtyTCb3g/klUrziDlGG43rQHzk61MrcyZpHpn+DPycoLXvz6ccJ3e1t/sUo4jMY7NS
y6IVjZQdRzvOn7EsD/YXXh6V67hlWA9F9kIZU8J+BSDd9bC9wMJ0a5mNZ5BFA9PXvAja7ij+NYRw
9BUyTrPTqX5aOJ5xHp69dy87UQ4FEeRXuGfv6rW+Lkq5HafedVgurKaWC0I9k7wv/S000mJD5mtJ
QCVm4Pgpon+NP13y4YW+eEPuoW7Olr2aWP7QEvv3G09cP/L2sbL4I3lRcQTkjC2SdYykgCLDXhTE
4Oj2ZYLL9MoIygzqpppKZttpefJvIXWwcBJM1CeR2XfoVA1J1LhqDnOIuHBUu+jCi8EDE9BjBJfX
tkDu0HjSCvMZDFY1jauuUUk9SZJfULAD76Kt2IebWxkYnEyyuglEvgEl1dAlcmPkEf9zkB7Gd6tK
gj6l4LI7VSZglIBRxnT0MyZgR2apPV2dSxYWBmsTdGngw/b1i5Mbky7Ab/SWYse8rseOnX/Pnp3H
zAZ+YGa9X6wPvk2C77EshUsjkVDGJn/sJ+TN6bwqcxpAVODPTINozGdAVHTY2YYSQoy8TsMlkCho
eWHOq35ukn2YGenndb4gMUCP/kMUpSUbGSa3Gb1mz7JiS/Pl1L9DrA/je5/DQwA73Lu23t5gufP3
Ug+NiHrgshcgbSDlhlTdczaKkWOa9U6pFnkltBpTx9JTxDaZDtLpmhVWeMGD+T7DfEz9OYzu0SiX
+NNleEB6x2Ti/3BT6wWD/VVFBDXPgsu9xXz5qAxdFsa5P08i2az8d6g+x9fS9ILzkDLZBQjE2PAE
QpUG5FYcpfnQ9t6WALB+nEYg1MYoBiRQo+ad0N58OXL7mFqNma5zm6y1SC/iwAIUk/i1OQs8ezyO
CQyOahNFJu/IJzbrvE5u4Wf5LX5GCkn5S1ZU4Kp7e8w0nGqiu2nsxnBnSqGdaZFIFY7GVx6jLkP5
ZqV16wVdXoqsWleRJAInlI0RaN6r+Y3ye+BV6mRS4nOrtDytP9U991nMBbIzNul2ZAxw070PoiqZ
5Wy5oHzhcmQmVUBJadLjLupDTxwCU6XC+lDZDpWALQb0y5UWXBZ92UcryF9qTKq37GV7TBy1CVg9
YFMwXUiIibWqsuU0nODI3cAqzU3X7esPuJU7xVvCs8RNuACoplT4DYghA1xP61n4vBcKkqOaNVHl
gOZKZhwtqYMAnKw7dM1OiFpi+mzHBLxXX5jT7XoQmWuozhPOwRPST4s+dy6s/WSkmGCgiTaRhfU9
Ksa38uJFHf6Wkfq3xb1G8fgQzMZ6m3r59ZL98KqyQnrngCg9NfjpdoWxSG3wGXHelOATiT2ENWpY
pU4uxVqiQtxyWMH2eIZrPUClbeEpK2bCyBR5Sa5dZlj4i3OVFjnQbHEH7j+sf6sV/26SjEY4Nh+c
MXlwIBkr/qDbuNMNvNCDFQTDxuq6NTMjxyi/u+jwrnkYnjx9bQQ1z20gKkGMlxoXTxN2NNtCVkTL
MS4bLS7XV2wXjApNjG6/ra+V+g0OncybaHDFGCrkrvBVvTXcJQfAAQS2xv85yDAWD6DHU8peHcuG
tbeDTrvUnRElSNDc2p5IU9I7aoU97QGqqJMzS8N9SegbkTWuhzpYtYqYELKHdCBvQzz+CKCOuT5+
jVmSjYcVJbmM/2i4efFqpgKjWKuJjO8B3a5OyYWVPu/H/4gBOBC81QJ1jZkWtlmRgekaIEA/xaHK
JRL9j02shCmITZ+CsZihzAgYBXeUALyEKA41o4gmWh9v/guRzCNLU/37aeEiePhY0ICgycJeXvVu
MU7wVZgqMXUd1fNCUNuETHIkxXMpopshobuhUvfykfb51pQDbMrjUUDpq+UpSzWF2yqZbC8yI4gD
VGjkEg3aKOBsM89p59yLNL2aARrc9dgxTV/uq6sap9LLaxMb8xPOecbWlVkKF1HRule7bBxXWhOr
cpLGVFV6XhSNE8VO3bTlnZKo4EApTRxK3Q3O8Ni+BUV0eH2N1hDDOpB7867kRQ6/KWwg7eCIs/Iy
rlOTibtnyCG4h9XwzMD+Gt9Dj9Ad9pRa+S54/1ZlNbp3ms3APmpaAT9ZAmss2YdsuHed/Yp8fNLM
hRPO/i+EC0pfJbLZBu+Dot8uOSaZfcdvYUJmh2jVw9amdhUlsHYQ1eV8KC4MOH+cbtjZT+khrjRa
yNxYKVV2JXT+ozhTQB8vBIwkhDHfNNZ0DNXvzkytRSDptlaZGSBoE3RWW4ylNDmwjOGK5Yz4iruO
ml1MAgkcNw+UA4iRvedp6hPUaggoK9JYS7TC+zGJ42cN0lAXeVezPw4xxeE8fE2wTKvUIqPuZpln
1+1jfoK28Cu+432iexgUgFs4J1JPNTN3gzMZ9f8WeoYnLrxsFfj+wwoTpsgQlpekSNx7B3GUL6Wd
yPi4kiAsJmZibGsvNvKE30G3LpIginGskcs0W2+oXeTb1URiQYZKFNODznHkVvSZPJvnlTl9YHoF
9O4cHIOazbSCrOPZ8BTv1s8qOlYcV4Oemb9jfb4wa+5qPQAeB6GJTs7sJE0F+0DR3iNOHqz8Jy+U
u0gjiExIlMSOTxHA72AIVHgJyP3GBwE//6g2t2H16n/0DYS/Of0rgPQAp+gVCpXd0aOhXNYBQ9uX
VlFE0ECl2JP9dsfL8xLykoOSuhHWXxvo7H1ZiYq/t6/1bgRrODh55uruKuwE5pPSVcewWiFlBPXo
6em5tqtPYVmYxQbW0uulEZCneTVpVsxvRtZucDINAPKQhgFR9JHfcJ7fFQKrB42uASzSrKWXIgz2
RJSSgr+T3/YE8giPucM/eq2c3SJf9t2gcrHSnyeraOWFUGzxB7YT44GIUMtd98JZNKPhR80pa4DK
tn7f+pJEQwj1GpcWLSa7pHhB2d4U1Nr4xzkN1xOY5Hqx1JJFftXw3Dfjk+fMhigo4qSVEAA9ZEWD
3CpKUBcWZto6TGWTyIpAPkDMLEACbB62HtqyNJYjbYlWPceaMxUFG0D/Tq3FgjHL2/qM4kM+a2hh
RP5qGzPJQ5S8rpkFwb2AHeYx71VQkZBcz5kftDVEXOMfpbYqQWw6cegjOpy0/lOkZDm4ahYnpk5C
6/4GxhZ4Cne2dWUwml6NtTOpa3cVxEdDcsO+Y3/xnwMfMXj7F8rjcb0V6gkelcqN5e6m/gtcgA7L
HyTcO6pThx16m0SIMhNr+IjaixCFN1GbRRLR6NXHYPJsjux84AqT1HHBuJpAnmwOju5PeIk6wM/7
0kvxVHBSc0TgglZCyFF4d+nrSJJdNApcVk6IGDj5McsIdNy1dGhU9HkO9mghbN3y60cGglrmKIM4
LFU86lmfIlqbDeB0GuekWxW2MDxOwe/njThzJ8byvZ6RMJRsbb15wQiMANtsEslHVculhHgpiDAA
SiR3TZIiYd4yC+qmDZkCjnKCYlPzq9ykOdQFgfwnH6goaykAEtmQDxze6cqKAiOM6tEAsy7XhefJ
sADsWHOkfe3bfMH5SVXpScaaZFWH6NHSD4V4U/NMA/9BE9eTsHWWccOIedyScdAS+dHGO5zYBy07
VjvFuW7KIe4FzQC+V52U4O0WHkmoKICGXaLD0blqHXe4ilgTRAoZGpbnN3NA/ImtA9mBhtPZmsDc
/JsYyl+wnB4B3Ss/zSfCOWnATUx+YXszJn6XGbz48i44p4tsv8COrgUsgrByxXf3Ud/46CnUKTw0
5t8p3JYX/R8CQnXm/F3W4xajvUOcTfeJ8J+VQ3KLy7MHTJdGU39sKuheXLRPb4wqEvQYwb5gTGwB
Q4I8bPT1NPSRe9LM8dWIfI3IP41WncpKxp0XlvzPqLCqDEoRL7nt1tz/d8DBJeg9wityz80DyYh8
J6v/BfzG4yTm5RTDc9ejjSPZJoGALMNvMo2NLhzLv2BsjQJCakHpEyv9sAKkOCRRYHOqmcvvuY1y
jUgpJH/2eOdJo+kyC+3KLQDB+VpIGn5ts9CwbY85t3hqck0VGO2Uen8Gki4ZhfVK8jGdhYoeaORu
E8vSt3zQozTmAaAJnm0uvXkSmTGMRjFKgfL7h6H4gt/8V94uliQmtt/71vctoIToPsFPffho1Cnc
PAEPulQJVTCCfQ8odRr0gGra4Bo5jsyuamOZJ6bvXtfI54aLsEjZL/kBLrAvxSQWTDNatXrApSp1
2cL7CmXP6wuAmrOhkSbGP03s+guSAiGw3Y/eYW4MHRWQ/OBvX1BXXo4qERx5v3kfw/dDuUHKmuS+
vuiiIgcTUWQS3oCm+ScbOPxOnek4ZyX7TY7gXXeOWlChU7ZESVersd2OqE+4X2uLBWM/iY4GOdcs
HD7T4sjGwNUw4BQER/BS4AO0E89KB2xWmMQ6lS9OG80je7ESRj8cK0SsKr4Y8mcYvRfOflgHw7EZ
lAVc/0wu1MVWZ+dTlxKr2bRfHe7ALdXlHUC5DmdFUp43S/txctBfdV4pooB78leu4UyBY0MXnZxZ
MrBY108YTX1Lkemz4VCsTIKFNXMtvAMdznrIHM2ECZTN06jPeuNRZLddyHv6K9DDct0ZdbnPMw2m
nZI9gja6UnNM4FeKKDfP3d5VEySEVuEy3/hinXudvA9K8L/4zTDMt6Tow/Iz3E9HUveM2MC3/nPC
uDtlXFM6BdjPgJ6NpTKPs5QyGTJFWlf28+WllHLyk78HHtrTeq8G9aO+9Os43CuUyDKbm5n+8bXz
VVXfXJS2F5JC1btaQqSHBuOiSTlWR7RP92z0Hd/ZuXVeqJ+azjMfeSXtPis/+4KYRRHYodURUei1
B5BfQjc2vPJP7jkzOuuWolw+KgrR8uFLJ1k6g5LkikNur+n+v28qFzU4hZOLvMGYAUNKWYbMFaZg
RCgKjiIwGBrL3mPrO3txtf4vMdGb3sb6cz+2RhVWsw2v7OHVAJztQO9V47c20CAL1MVUvxhyQa6j
+E1xT6jaSOUsuE95NlGBBq5WRUSdxk09XzWtUYCJqRXOZFw15CJiB8Xw2eAY4SNoai9qxUR7OWyE
v/4SvD6GQg9KxBY8SybFH2roy1j3sQDHKdhQEuLtsqiJ+toyqO0dnxLjlgRFwiknLWkzc9fXxMIC
k/KLkk6RiKcD2V7cn5bz4DG0j3w+aX8i59HQ/nFqRAYsaLGYdQsyF9a5UwYs9/EFkHjMY8ThdP9f
KKm9uigfp3V6dNNxwO1ZHoDRHsNJaufa9FFeiXMBqCQSTWJkSDUQDqqdEQR4m2QLaumpb3j/Sgel
BnP3tJugViRCZmRLj5GZREeAJskZBZorf52yL4xAoD2u+WWrTg1p+yq57E8ZscLYoc3b59rdJEXb
RlZch9bTgkoCGlt0cx0Pb55q60BfqgXp5lDZ8r6mVN0lL3fVn/ADdvX34JjcQh18U3hKDsPeMwwP
rcd39wJuR6Wi8zD+Wul9njjWrMan8+1XqNDT1FKl2lcR+Zmm9Hm8UOY4cpmfjoaqz8ccNOUnLpsn
wguqw8cB8+w15MX/fRJHP4ScqupzjzTWyOCdhGpYqEtC+WL0eOLYH87eZvcVySGFRBfVxBTFy7IG
f/rwXOmpWyiwvdvZ5FUh6gjzyqGA98+cEjkzdhYHqtZ6E9zBos8bXKADDkcZiQS9+YB9FETKENJI
rTln5qPYvYzhCpOzQF8JG0AkN7HkCEsbdOCKSPDN+lo15Gj3NTTpVdfbGSyM2LOkxg2DrhsHMXMs
fkMcMXCXct0BSy365Z3WXTDWa1dBR8QO1AuXR59cBpF62xpRppGrHwl/KujskAy8ZD/DgeBCfdCv
gGoUqOWViBRRHqYd6Z33DnisSH5xp8TEXeJzJmmFsKk1KQg73uUWxaL7WMk2RoemsHIxTDOFE6zR
K0cqEip/bWBYoNTlasmCvamqZTAKA2TXNJi2s57/oZIKMAHS2B3nE+rO8Dk6/rK1YKWuysdjGT78
H8Hs0SoltsQkEOEyhfE9I8rbYgmDMCwNZuVj+vHTuK5cCYHrNH8+AIMF7f0ONbuZntpUj41j6fK3
QVXfJi5h01lBSy+kUlJhVxvI+0NxVLbv+47J7THe9zz8zsUOoaf0asCCzd9fePD+9sBN0dhJ/1NN
SWKdlOqkA6fZHyk9HPTkd+FDROOL6QwYvhgjTuONhNQm26XnAxWefio7E6x9zyLvx8DBj95sbMcH
m+8qaaC7HmDXVU5VFu5xgq0m6T98jTzB4i7cC6YtnZTZEczXUCIGqu5UMGYm3KtPoNX2EQZ89lr1
FXjUzSuxF+aXgyONkmkIeQjZ/YzzLSZOh48VkMxmNzRcsSMchaI2PEYXu1DAdwHWbXSPl5Ze0Tgj
PVRO4dWmjhbm7PRxz6RfgcAtMgtKk0HzBFhpE6OjyjMTqXpBq3dGq43TyHoyTaqn6usq/rqX29yH
8rRFF5IOoQl5WoD95YHio4ZxgLFVKpJcPJ6B119ropm5r4+nQtcH5lzlg9d1JwV/r+Z2cGqbi/bh
77w8UnSYFkFjV20ktijEfO7AwwaFQPcBjx6ZQPu29gVPxfZi5ldGLXkkFhzk94lq36qZ9jAZ+rnk
uYMS5SYb0OS621rlJXXW6DdXTQX6MyoTK5HHAgOaQVaVdnw/gzzBwIi3nZ3LjXT090rae1BOMh1x
ybXVV1yETaXOgIwSw0odvHsw9mHitC7e4gunEls5dt9ODitlDYZHvDoAdfYrpuMGZv79bldE1hNF
ydA+i5LP9LA8xW/1VEAg+nnBlsS8nx3gqvvvoi1vEVpDFXi38tBvQUcc78WB+S2bim7y6sCYXe9g
njmde2rTKrlU+3O15SgVZticHTK6bqUxDP6C9fhC6NDzeABA3EOT1sOKGySIUaJvECmi2w61/nzM
CD0jJpN4XP6PFneJxX5xP3UGgjaUoiRUVxkX7jIs8E1Pp0xJ9X4Qra4eqvsIn4oOQUItmoZ+OLhX
3DLjnrm4uQoGTy2nC2ye+Rdnw9+o4Hp87xCmoOLFVdzbmszB4aul5xdXgqdPhI5mwUZzdNjCuTYQ
zP0DyhwW2JpmRXDkPUi6xs7nfIaX7ER1qWa11/J79VO/wLpYXJK/YsRO5ZreR6FDBmAyLUF5YcIR
vTNx3kxPxiHsMWWBXJqYonlFkpjNpu5Lzhc3jt0CFsoCgj6EEKAN0S0v3nPvNrqtb/2IKD2ery28
mviSCjBcIv6JD26I6m1EOS+7wsj0E0D+H5kiiWJKcTvEBtK4s3rVrNKg13CY6PFHB8WrU4DgalBF
PDFT6X+MtzDoy1eM1TU6r87aeU6PXXSNBVTE2F4tVc8vKEBwQ+LsJpHVJC2KOwCrDyqIWKgLFHjw
pqk/fXod2HBNUjXri8yXcqxJuCXfMCJV9eoZ3sV4+R2YYc8PkhnqNom79ULP6h66Tg8Spls8H3Vc
sGEaTgZh8JPONLFYbNELYGX4FrQr6/M3SRGpxavBSrI87ako3P+ouMdcQF6eknu8yqfn0KNbzQrw
6OV4FcjSQJ6vlcwcBaxP6VY2G2A8/fXTwuAuhgg4RxwENSIBfsmy0Qt2L4/0bTZevspLTL7ixJrv
lW4rEj/KglFlyDXYBG7JJM+/SsiDn+S4ExrJ90c0TWk69kfPMI3coOMY8rU/deLWjnKKvW9dpGMr
HjgYgP3Q2HDd8xqqMwpXqDfdVWTrpaD9gbatz7hikLH4CU2JBxzu0/6xSHr1cFyGHSV9R1qf14qr
znOusy1gNBa+GkA5JlQiFzF/oDr+5twXiwCJxb4NJEIAesUljQM3Laxoj756wWXSMnv7IPpp5I1D
Cf0r2pXWh6JaO2+/ql02RB84y9XJAp5z4W40YGAhF7UeiJj94rV3IYiTKR5fzCMKv3Rs0+lPRGui
XssCxCqRR+mlPt9x5H4/prM1aPvKcuFhLCxXVNv+yMzcX7g7iRFP96mv3feqIBQThoeyuV2dai8a
jI6TfSfqOC6h2NZUt6Vr5M/TrZC73LAEWPizdzP3amilAIdvaPKEuw7x2/6wNo54nm6KtXgaI15N
UFznO4R2UWHribn8Y+2eZO5C0/MZIQMj7eI7ywZdL1O2UTZmv/lL1YaubB54oKZjxYwdLdpG7y77
L0HQoeRT4Fr9UgMwIkTvQaAxMqY9AZR8ymauRg/jgt/sEDAEjmJBN1jjF81ImF7ZGivWPDuqzv/G
9RRNWqu9TQtWeIEe8cGeb3OglzQPk5mfcXnbrY+CPBRf6/9+nOsIXTjLymKmQdYzOkmVVJ5Moxjt
Zn4uxdo/Uo8bh4JW8oOPfYnDQR6P3Gu2HQ/LITcqMuAEUlJXanS+K365StfZq2Q4GOogZLTfdwPH
vP/eDtSMZlbp3T6XK9DXuDKpZa//Y+Xpwtsti3LdKUFhJ++XEQlDJaUOiR21I73A2I3BfanwJ3i2
km0ShPK5Kx7f8pMMJpNpanT2C46gUe0LGgjgFfWruRxRT/bT9+X3kprIY7LnE9NK3BJl8qBrtHUO
0KmKLipmUFU9R0fC9hZQ8848mLCPmZu6LQyn8Mw8raa9jbYoyewmQn60hT3if9HnrKb21yk5YLDP
HKYlHTAWNyocdQZJ4cKHfbKuzhH+XgeX6RnFM4RmoKvyClLJSITg8nDxvL214FmMzWngwD6Gwq+L
R6SoBhnIkQd5q2AH8vHUQ8241K/Tju9DR0qJN+grOaHeIDTetjOY0u+VkLQO4x3M2S/G5Uipa2ZS
QwXXTok+NpG2QfNRsTdoWYyZAs2yo1uOpgTWvZciZzBD3Jwbsm4onTk2bZngUUD3hjX3r6Q9SZ8F
8uwrLs1Kc116eJlu35UaExi3LuhOtmGLvieRUfTa5YzkjsnMohmdDgjFQ3j+P+ydS1NlIaxFARx8
x0Znl2ADdZ1JpAMzjnfOjetSsWEyG4G8x5tC796Z9wzSWpoMQA4eToNFDzszW6tShSKEHc5IIj5T
832DPDto0NvrCzhVSqIOvDcsPxiyBxbFNfjL5h9/nccG+7WIsey7AETBizM0FDY8i2jVfhsRqqQT
AQQmM3qk/+LCnSnDSv+UCuKG8IMzcLQxGzqek2TLzjZ+5geAyM2vjXg42aMHSdIKs++Gui3eXfp/
Wa8lOceI6dlY2SK1iO8W99fegcRWq/tQp88vFYuPvvZQLrZhTYbt2N9FVd9YQcWHXzsoZ1wTwfrH
9EZNWGcoMKfr4JIc5EwxsDU+kBGT7Sh2Rzq6U4pnhJd4ivsLcOIHYqf5PDXt1o1b0bjoVoyGcNhh
hOh9OxmbaiHA2b9xOiNxyGjRNyEJNHv6jQ6ALqe5Nf1G4fsKs1UbwVtzHTrx5HdXoFkfwDZCWO0q
nfW0CFWGmI/IqaAE7xk9XZv3XdrZm0fD6tca2dvtyZ4JZqEaBMqi7l8cuXRtkQn24AA0YpAzRy03
0LSypI+8kas3ruwivznON76hfyETPE/LSHo//YjpRMokzB2zyHOYfS0XVRCxwpFnHfK6tUvl8Azi
eJTevfFtTFCnlgiZF+Dq8RyCyu54fUZI3B3PVBowhKlP44vYRb1ICK7Hm9gTlUhh7zpmlhFNEeUq
2rqP0+kUE8apDg5xP3TzcZ6lXsiWPCIMMiQxsJJuPiiEp2kYixCvIQO/WR6EvuitCOxNoJrA63MR
6kN8HxtH6VeRGzE1uCCfH2MfbWePV5iB0mJik4+QE0QUWQiiaA2ERzrppVs1bHwajjfdVULditHZ
vqigyeoKeBmzx8zTC9Qd+JzECatZNOR5VDYYE5WFMFf+40f2KhQvx8UL6IbcMPS9g5Dp0SMor1SL
pcGxreBUfKQeFGdIffca85RgUiiRQYMNo3BwWNVkFp95Km8J85O5fHAJj3KaZS0cIjQJ9mJutx/u
3e0y04o0rsheIp63j39GNSgkF5klVbPD2Z9/qCmcIv1W0x0HL/f7c1Ez3JS5wZNAc6vwBCkUNTXo
i1VDEQzvSsMXqhILxtkshbODWvOclc0bFa8bQ6Y9ZYkFbPSX5+ma9f50y9Bf5yCv/vWrkZMTPBUd
VUhBBrFVYs6kLJcXOM2K6Dgv1xXt7c8AomGO2bcjQTXlrasOuhNfDl6J8ntRdZ8skiyUhhsDns7V
Ajz9EQpzCwzKn8o9vEgbyKC5Qaz8G2kSxLPCS4Lz0zEcQdxn24yKEQkcJ6sIq+9zYXYey4gGg09c
Rt40IAKyrPODWvW25sEQsusBATBO+6VmARgbquIcATU7kUyCDFoYqhkxanvYRibDnQDyMqHrhs5D
Rw11lw2VHqr6x2q3uuJj9ZJ5kpCvgbrGbFTTqdD5ebhoqvxWRY/ltFTUfYbu4fMk/0fNlrbQwm8q
/vQaf7C5GBfhPFSeOp7DB/Skrk0gSGndiKeDx58Q37hWDCxTgfno7iv/T0l5fzvddgSLxeIQx6l/
CTi4WI9SdA5z2cwiXD7vOTskr4Mt2hAny2DMBObRlPKq4dAFT63TyW6fIOUqzM/ke90OoyNvBQYl
dh+OepSSM/5UTok0dr8j+3+RlZm/ekesjfVxuGN3cXBW6ZigmrpM8wcOb3nv4/gmTAEEH8W9nBxR
1Vog82KQUtr4HJalMagJq5W9ytFsNlxKKZpP4NiUJeCh27g59RD/bg2UEERhPdzq0a2k6Zi7pQWn
l5s/uPX8t2dNa3JtErBpFusPEWgQfHyd7KEXKvOQvlPVA+LcMTbc8rJNpS+Qh9kdMaOqpiqct7f7
xl/gVnPa3pItEmqAOENw5meuRCPNJYBd2JroO2may4UNJA3ta1FPf0hslbHdMhhwB3niCgcEn8Di
DyEU9hhzMa/YYNxMKDsOL9W6LSkkx0mOCTAj02/8f0hXug1Bf+9jSBBvzIAVfksKS0RjH+yYbdQs
BJarAxuvAmuh7QtB6dLp8ZONkY1Hatkash6GjqQXom1TNgTzvUUIL9fGf/OsHOQXOQGtxWwB6w27
u3Wszpd+aLZIneungFozXwpS2p+8rQJafmFKJCJnaHjMJ1m1jZLvfnJIEPOuSe69+jjE86dNF7xk
Yo+UdwZjbBlECyypiOrrZLvDtCO+4bT3dXnaaN6Z4YP0r+J/UVxC/HxJ7an3ZRz3xGTX+U/x2PKC
3k5V1x/SJuozvHGMZJFF4TXO2HWvz2d8vkW2aqKFEVBl+5qJdhcfsTOA3IMzoRSr+CkOtm+FpkOy
k/6hVSDBRAZylNx5TRhpKNei9mYRVztIOUSbtDyOA488kzslt5cgNNC8fr4OErgwgxJSFfF24VSn
PByuHmSokSIJBRqoglyZZkDerP7V715KQ10NSI3sMdDKG489rQh5kFc5A0mnoWhgkfQ33nkfCnRw
GJiL65WdBZuVBAEM3nWTs6BQbFXdnwlYpa/8Of89VnMj/0PZjvhizM/h480sdjtQjb8i0fGU6r1L
/4iJ30TtJm2cy9xf4HkoTsN78LxOFox6hc4jKY7RCSZOwuQ5LyPRigFp+xmdg7laJIfrY2VNEjcW
2O8yNH7Q78mG4XZFnDrttpR0iAUQM42djeQAk919PSpgXf57JnfMGxgwnN4rvft6W6VLS8/fa99q
/Z8YSzPVhHqiUrFVcEeUCidrzFxfCKg7hI6LUq6EHyACIVm1fTlU5tNpiP6yr9PJSOPnfeNK/xQz
nA8snAvj69T5ELr6EbdSdPMtPmBYnLG7/rNpP/hwgENi0lrf3vI89rNvATc0lX2t4+rd/bjY+zmL
ecQB3c8put6qGD3Z8KXH64gxXtjN8O2dlaR4kUF8kztkcUkeMrYKyBnjqLU0Slny9TiYV1/Z+1Lr
Y9a7iTZt1dfxl62588Zn8T2VXwNNOKDAIGqhChXShd/dJ3PaQhOgw5o8yVjVWwi9ssi4ZeRmVxg7
uSW05zSY36OWuFBn8YuFFug95fxc+dxtOTBuO6jYGjojPRLbabwffu4OoLnAxHf3Qf1AWhAeldUD
RqMY6shSd9Pxy4d5HETekmyMGKKJvZoh2GdNP4VYFbu/WhZy2a9tvV3U41PXnS5Iubg4HJAvTBKY
DSV+/3XhRdzoa2lWD/f9Gy2FRVKuxfPzD2cNZs0unCdikN4DDckBTPiwS6uy2QlC/uGttDupjYk6
OCADuvrNtOb6ZFsVXwOyGO7Uk5bDDmimsshjbUw/p7usW8Q41x8qhEo8J0jMLNO1NpXPiIhdFugE
HJWJOxrtCWAq+bll5+lnyrir2479ZA6S2sAN6QWBMtxLPIgf1Vm4OSvD4aD4B7X04vg7zqfor5Dq
0ljRzXHxMSFbY7qmXatBJ38z4rmUqJv4PNsOZokIVb+xxZkhZqsdhnyuriA8DzSmhB/HLo2dYJoo
Vcb/PoTi4O6wtYgRq2XiiNbnyCNib6SkAR1+YBOjTJUR6EslZrU7uR9a/lS3F9LqXk3B5RmRRvvx
oK0BkVb4AX44UZEoAFwirLPwmTvL0cSKw5avBZ0BlZYlDG+7Obxwa9arYBJX/jFfSZ2O7aME8pII
sMUfoK8K/IlQJVTmP0cdZay0qiPi0Ox9wOPzyGNtNpyHPGhLxWNCWr13l60Xtv3MiEakmW0xE7bl
LfzKni73K9knZcfH+Z/i7eTe3H4zUoLq6EENl29CGUUoIq89n+eQASP9u8gDJQcvJiAvxlMQzRd9
1LkZILKx8YHQkQBD0Ju+aQzYYbA8K34BhxaogZsoy6qK1Lkj286oangWbqUYNAkyIve0qefdHe+g
dsjGfqs67hWR5CU2Lb4gPEtKoHnCFnQAwNSPSoC4RHe+Z2kfFLUCRl7Gl7DE9jcUSxWDtux1oqNF
w5TYFk5kniM8CGa+hZkaKUup1FxMUeQZ34WE3u3dI1idi66KuatBV2lkb71PE1nwgPyRh7npNOEj
nLsLA4KaI7fGyVwvp57VmOdVBChIlUI70G/4NhVjlu+kvuYhfud0tpvUbTFkb1RypHFeIkw/EfWb
Ain3uV54Sw0ksujcu+xZRbkCirsdnASYWpAhbaItIW36bhZ818W5CqzMlqlEawfKVTI8bQnpqBjA
SpFa0LL4BKj0ChN0YMLSGkkKqUc+eWDhslIalXd86LNXSkn1ATs2o8ExEsPiOxtt/f1AqA8ZlMGt
AgFUJvCULmRbrCnYMkWkbLsKgXsde7beb6fOZ5WPLPf/Fum4hiRTSgJLa2A3pchCPKBTTEMCLi4D
X71J8DRCbYBH0LItpuNy6Bvf7J9C+4BLcfSQosyri/eL1ek6eALPJih0LPGZRbaL1xrOg0pb+b93
1Ra9dmmJp6PzUQMbbduT9YdQ3+C6PI/11yCcuvV0whr9wZee4Khfk7cDfagfsGEzk+5iQamGqtkF
ogRmIeTHzXltcN/DJx5+2+r1mMYzmZMcwe2LgkmeixN9DklqlgIBTOEsxMLKD8mLmm43d9FFeZy6
K2XhJqnBHeFQXy4HOLL5K06P0++YN1N2yG7ubG6gOOcZ2q19LPB4SYpWLLlE/CvGxIA6nZVYpPIP
QF30Dgh6P/FNH/wVx5iwP0Y5dr9tF4KxKTCOEEOTCdrzJX6fTvgsFiQiej9keCA4ZazWoLDWzzGO
c6bBjUvWiR/nVx27Dz8ILlP8JKSvuvo/dYW+BTipvJ6n/NDRoXBXNRVuJW/lDVgXXFTiwLy9Vl8c
9+fAxgz8vYOt2MEIlni3RsCIcbKDFzVrAF6oSZxtk43oLopBsHlLnrvH2bB4xDn5UWXUKdgOlmRg
YD5/QhLTaGE1IIVYHSre2EyJ3QiRHb2GiEVBkoJq3pd2yqPT69LVu10mV3HedNcuondetKg3v6Py
3KZgpdWw9oc8y+r5K9FB8nXL9AaFslsJ1QeIRwhQ1w86nr6lW1/bIjIf+AcscGd/J03ugTBwvtST
xlVO103s50KC4Ek3icxgmA0DteOynqhaacjgv2eYEhaz7R2bBs8Xza4PHdJIVoJ+HrKyXsJ8qUBS
WSicQCo3UbPXDMgjlKsiYi4uQCFp5+/EGj0Z8zvWAm2FaBrsTPavHa8dYo7ll4gQNxCSPknvXXIW
R+lPBT8Oqsa68hHxuRyYcikM4MlUXamx/kaDezK9aT/+15XmYoLzzSsfl8dZapWtjQSF2CysRKZ4
cvk1/QMklI9TlKfVKnAiJQDYPo696PRZI1CyOWCqFS9/8TO0kitX6RCQFab2E66h4TCLABOVzTsR
EFH1+MI5kmiT3LmBLu+kX11hKH10B40veuvVPYnWcXlrN5/ELEsc0EfBF8jkU2Y7NgBbCH7Un4we
59ghoUjfvt99LQSfdP31QavjT6LLnYMJstEi1hoqpcqY/YDeG3aSzD6cDyuIFkYmiDmMESpYaa19
LTYMJ/ROMZu7WJcLa6n1ztSEIIct0IynKdC68NCCmohAXjKS67SeJXEsxxUHJB3HMJH9rD2hDmHE
IK13fGLwgWQZ5rXq/9gSMq93Xd85LQPIhoKmbYBIAqoJbzDZGfi2KSRe4ed2iH7yYAO5xcHWwC5N
yq9PhKH6oRiBTZ5q+2PSWaqPZAVXX3q/ic1ZrKWr6667uBdTNaFn9Xrd3oyve+bOJCt3se1eFzlD
HRdjSHd/vJZex/wvJPaXnP1bhbLv8w0yJsKN1AEfGvPETqbbaH5OP7iQ7mn4uOMHtsTfQPKKdTkF
25NEni4Y9RAerNKleH0Ep/TCavWk7wpRpUf5huoBYci2Qz1ZaA8WRJ3EoGeROC/j2rlENdaaRsE1
zODcwAM1MlHmuV37LrIaSI4pUah8ubH2nBVFKOxXZITyV/9SEOspmpVWzkkEnNZQFov82C+ycRnW
BdyTbhRZwlK07jq6vmj8MY9E7MynP9vr69dR9yAYlnUv1Ci2cPcXKpI97WbwVWNfnHRuVY2zy8x/
iSpGBpXFWtuZvdoftZ7VWSPKPiS1/eDFVCqU098BW/6mkuNcdcV8344lBycdbVUVE8RUs/4Fo4M6
JiC4MmzBv6LLwWqMByHM09V+9nVaFyHUx61mLtNkPRSm6uugUqBGi8LSgwJYT74RqrFN1UOdioDB
pRlZa14zNFedwCO/4LIMbwbHaY5Onf9Kb2wbu7ZVjyOYPKoJEB46e3DgTTC+zdpJKcNUG7GUrYiE
Nl2CXud8e8vIwe1Jxtfhi+kcCpWW5MRTrjQhMxpi6BM+QS9pPAcJ4YGqM1j+7HjPgZkAlJn0gCsJ
WwrT+o2ad5NwZcQpm1deDOEU0wQtjlt5A8vzCNCc8mu23u0UvL5SCm9FCvL7Ykv+MxE6sWK1xTGr
ox2oz58/PI57C8ObwKgx8x9w26DnwVzZhFdszX8yf7o9sjBITm4M1XH0u/fyJ+3Z81a97hZpUhYt
ErE4Pu8nsHn3k4y1C6/7scZVSWag0R1fUNzSnjqFk0wQ542H8167hoVBPuHFF81sBuHuTFjyV4Yo
jJm6R0KJM+B204FowDeZ+68JsiuH970j0z83Cn3d+lsszUSc6Dti73EkeEOLxF8UEJODCSxRYcxV
18tUZlubXptk+me3yg+kkdc6Q5qFjJXvZ5ouFNKK3s3RKrQTh5CcLUomcGgAvxGJAw9M98WcrSdI
pagqTAiiEIqPfzdFeDQYNVi9atU2MA9KZZy+l2UD7krDekHRMKMC+t4lU/2v3/IWN4CbIUBrUxln
glmof3poSZJuf3hE6/sKYJstCpkl1rZD8RzqNiyTb/GyNtHuuEKHRGYqmU5rnOUMurDurhI1tYYc
J9XbscdiPCrHjOQmZqa/7G3hQslwO+r3x0pYdbAyUhTaCjNriarE93b4GkhdWuHXdpWSc+nE0OUy
oDPOVlYs51Ax71uqEcDhLiZPUjqL4CieTBRt5C9Vz4y69elNrmI+BmXw+CFoLmfh/Rj+js6ufFYr
ju5R3s89Iss2UU3fEE4MG5sYwKomTC5M4aJDj+nzU921/IxcIBN3gtE3M1CbLNpl1gZ8LCBcuWWO
NPNkcvauZhMnAg8Y4mZi8yTv4/0Zd6Ao1VvL2ttfy913eVjotHSlYNYzood+OYddAR1zPW9X11p5
PsuGUVrwSB+iP+GjqmyrcL/mNAV0sXUXiFGu01RZV6pjoZw68A+KSnCYh1nibEQykukwOmwvs14q
IZ0/8swifUEzJVQNcg3W7fiSzJm8aUrpflitk08wFl//o61lSZhVHlY37QrOcGT5aYwyAPyrEV79
+XU2C2Txt5Dcp9abMddPq7ksGLNVTT4KHwGtZxcQJEUzM1jzSB6X5vKZ7yo4A87T6h72tmTtnYGq
ToKC+AsC/wDzEPZAcL2LGvawOHXwex5SNrb4NlHq9/xE4rOaS7MJ34QBYMj6ankVWphv+rmNlODT
JoE34VQdVygKDYYNzwptNKVE0WRhJxQxNDkjjNx+zU0E7bZvfTVagpyI4WkwLXskRXIg/EaWYbLv
frOd8pi9bhtaWeGtkS4cpBJqvLU2j6Ad+L5WtHLDKY/C1kNnX6PqL8ri8sbMfEGGhM8K95Ts9VqM
WZ66ai+ky3PMwhdJUyFWEMnRBfLp2K7T1tjQz8z838E9maUzKVrgz1WqlM2Frwj8jZNbxxy7CwyE
PaidHk/5XrWyWqigb0DUhAjbvUKIodaWuO+VlmO9SerE6i5I627D4tLfCzhK9a3ABjaeBzHcSy13
6YkCYLMJbYMAAINvFOs6eLPIaUOGKq88uUlPIFeQYwZOAp3AaUaMdbFVdihlBu+wjAiBWyocyDFM
sHy0679lHJF/75bjk5z9wZF6Oy49W6MZtxW4BTJdpzo4+9Ih5Xw4BRxCH3OIHlVQTpnhEV9LsLyC
HI3AX0Y8ufXO9XtowaFQAkxlP31bqBIoewFMK1nVKYcZyJ/RA7wRdVSaOO0kZ6pxB6yBGgR/lrLJ
6pBLNYQH2s5P+07XHSFkqgbYwnJrcPixJOdOQ+cFYxCXVo/bEV7gc8IXPn45clFvanraaFjUY9Ir
npicmdZJLlx7PD3Ya4LxFWlb18gAEmfT+rod3lLAmC64eEQzzm/ouXomg6MZneMMwo7QjUVTw8nz
230S71C9gqaCybLz9MX17L0rLFdGkHh7oRT8kUwIGJ3QAuS3o/GATLK7ewIIGjFLFxeZ7dStSkQu
Qd50koDQ4vq8Pq3IXkd8Gd9kJDSpIZjClXIukkPw+aroelzvV/6tww6BFrIwuzO3jqy3SuntENeo
IyZZ9op/BxKjAOTDI1eyomB/3eiflj8IA5Sq57GrT4nJSSCNKIhmlDmC6Eqvg40XdAZRllyr1COP
SiRwRVkpc/fsT5rQsX8mwu+m9mICGt+4GEykwo/Dnm6/lCNM6It81tiG88TuG7+xwpTo3vAgryGo
yhOeb+8/BVC0Gjp4fA2TV4Kn1uEr0h97dCwo2b6XAyYy+wD++AqpLtFSQrJlDczjJr2/hQK8tW27
kYkg8HzfReMezEkzML/IWnWv8X6gzAhSNGWXoFQDBYaRfpU5bse9f+JZekLv5fLmY40ajGTmJJCd
Q8FqFwV3Ugz4b47aq+F+dn+B63nNkZpd2pMpoFvnwfLZ/jCthiUbFW4rS6O7+mSoSpHlOArbFkZz
kOhlt6Fn/E7t7lOaCbJxtH71O+wTuAwJ4+ph7Q/ZympwpH4zKAr9vM4E/BaZCkFJCZH+b/pI9W6I
P4hJ3pMMCteSTYEAAEwracusmoV9z755H9vkg8K+G5ebOp1M55Cv+ZbQ9LaFt3WyHlUsvIQxua23
/UyTDSNJOd8kzZofBt3Xr+uTDcSxmPHAVnchEnqAteyrrksZtPMcB/XUd+0JFtyEaJBVNcKX2jMU
yrTELb7He53ZkG+XRH/rtAwaF1G/7TP/PuUst78LDZR+lvqN7tTAlJQmqi0qjBLk25QCThgB1f0t
ybwwogcO/MDTSxygXXd1T0Q3qz+9Be+bCM407c+2RZ32wu++QzI71EA2A1p02C/BIJhLq5qbgryf
CPuWmD75u8666idT29wfFmBhZzmVtEov4MeIgZkm6ECvr3C4eBD0jHaxdY6MlmFQ3iODUWk3al9f
gHxenNMTrsWd1s4xByopNA2iIOAuEZvxZ/mpdK+VIWoDHsUz0MR/AQM1qbGnVi/WgUDB95vnNinV
u+FYECilARXJ0zprIhdIe8R2czSYhF2lNQqTtusULGQhtVMq7bGQEpvvgd7mTGSoT7v3Q21d/Xc4
iXYzr7rwyxyfn6qLDdjmUIasS5wvDchv8fx+IOItcvI8XkkirY6EOVm5sSeIy9+kbMm7oIy9cxd0
gAOVv8tCp2CIatCO3QQESx3G4RCfBuJ7T2JUJ935umwsukuSgPiGjve+iGepShQoICnQwA3CQosi
Q2j4PYwNU61kamrTr6zbb1O1RMvh4aL37ClfvDQ+ER9KmeFxmUSlu/atunRaDk2Jz6fXzC/hy8TF
C+wc/danWqV8W7fqdOWU9oCAWuM7KGfl/sZiLTCT+3iAu9hx0OCGEnY+BI7r+NOMXZdEJ0g2oYLB
3bQU4Zdz5sarbjcel1gUorSc5Qz/zjv1/2gfLKiBO1sHYTox+9Yu2CMzR4JeX+6ZApzDrLPX1Zh7
746fdBqYpdZyHbheZy5zWsVnLeQilAbgi64d9q4flu+DQwCGbBiy6u7Sjs5pZmnuPOk5FbsuUKna
DifmoBiR8wtSCuGxF+Ep3Jx3PmQKwjseIS+zM9Jnm7c35PLoV48i/jKwyacKk7Ac7cA4OdxB8Qtz
ZtNpUtA8keTKF7zK00AX3fFP5S2tnCi4vmxeQ3T1n3GlQQn6VETluGmBZZ/kSFz47UA/mCwlvJOg
/+xBcL+GTfK8PUo/dXYgbIYNINrPgzX2HuBiD0OxN3B9VQXkLDi/XBbZK5cCIx8ik1r14texW4/L
xmIiK7TYfRMUC5uQBOkZ8/GPkSNgwMAjdHvBOxxsmnXH11x741wwIPDzmtWy2a6IYyw2yudrf2kl
YLeG4hFkrlBw3ZYPBWA8fChvClB928ynX57I1oTqNTuMj0wzeBXGT399cJJwUPahdXKxxQRUy4h+
9RKmjKVY7u8f82xGu4YockHZleEP5+oOpMNwemHPHWVdG0KLj8hQsmou6FDDYJe0LXu3f6XT/AmJ
4tfhgz1Sneeulea2ueCZcCF1c3zjVLUMv7JN8MwPxQlWssepZ1WLrIpIcQx18H/I6mTcQ0XUKrox
S48T0EG5p8cy/RLc737E8iJF0OyBoMzG3cedTRRQwnMSbPtHaTu30XTYLg4ClWYjzLVsyePFGs72
fLbqIr/Cw2LMgXKoqNW/X3zmujV9uYOAIMxZkKl/Qoyicf+UjSWgEOAIwttR5CUYKK3tTf2RcsVB
CJxBk7nMz7gXq1SeAfi9wg4zK+3/vy/f4MxnLVNk6kI3z/pj3uVQyHPOXw9ijGS7pYEs102WqlJ+
cNdf/bjIoCKpyDZgD1VKiQ9wz7ptjCwAJkhxuxDMRgFz1omYnaSt1xA0Kar6Jf+5Z/gI6gMg41LS
FlMoWjjvWpetmdDL0Xs3dUVnCiB6NpX/z9j/hfpAvv6fX/8K36gtvzptOtKOgmx/O9KzPDGNJU8j
lPp78Ji9v01pAQ3cFawCBXqB5nphAth7xTOx4XtySA7pYbmk24pcN2cF02RzXAqHE3f1DZxX5jAp
LtE/mGt7IP0bcOxCGBqBxlrqO19sJxCOyA/ZqZgXz29G6o5C+ubIsAw/VQqa5V/NuwMB4tH1t1ZG
GK8drjmZc9xoAMuTuRLbFDSge8jVmb/Tw1NCEnh/f9UeXr5xvRSi+wZbF093gtTBvd/uhyFEJ0t5
+nHIx6nvu++kRU4Cx/1/Nzqat3zAcQh5WHeNSMyt5sX6O2surQG3FKjC0wqyOhx0kifoDn2Hrdcj
Q4bBAQ7ybR0C0gi5G3q1Lku8h4+Hxeb39rS3LeS7CVfya18gKKNuVuDZYf1C9b3uTWtaATFp7/K2
iLmu29iDKn9oE0gSA/khznLt65YwcgcjhYE5Ik60P2Sl9CLBdR/Yoalj4UrhgEl3e9agAF6EVFzf
LPQPwLE0XC+zck6G14jFhunI/5nswNNlnZH3B8Pt9vsUJNoVAy32XtZ+pIBva4JcTEe/EuHQPpAW
5s7mmHa+gNyOH4/mCTsveKLIsT0SIBT7ipzBKnLHpsRISiC6JSFuw1jUWLBLyFEmN48ezXSfOFCP
SmG8oHNB8LNzhRr7bIa4ebW/pr4us2tUw2SNg2jhexUVNHP5G6LMB+4DnVzWd4YuZ5YRVxJZY0Dj
rp1zNMNZR6NHlfOxpAOf+9tDI/liY7GbgXLC6ExhOEqeZ45K3X8OagyiSrK9R2qRVOiJjwLe+k93
zy0kZUXte4ckKTQhRyMK6S370ZpFRQ5Pu9FoPp4aacxxw0Zpbb0ZkV5RkmwJfLNS+TjFhI2xd4XE
9/pxs470WGMvQDmExiLtIhhsCtZiGyz/sCvB1ezMKpK7ilT1NZIqmj45vabPBflvVLhJQMrwT6k5
0TMS62ourFe5n/B7WzHBObKFrMgA37RKwox/64xsiK7n8MAYwb7VRCCSywY7lVYe0R3elxTdUfk/
8nu8Tv+oPZfG9m0La6H6ba4uMX9kvx1SbNpzBa5GgdQGr2eOLGaMGKwG2aNTcvN13AeZosQ35DUf
lwU1m2bpfF0NQjPYRqW/Or3imi1p/iYhD4EpRVNAuRXEw9GSKcJ3o9GVAyUXYxyFGNibjxe4b7l0
6NSQ365k7rfozOFpNpN3o+q0U3+p3WwdYvnhTmAhhPY0ZUrOyA6ne4MA5efG+Y2KFA1yQpgXIxiW
/J2bmdncArLx0dqyMWDZ8rq8wQUwzcECrNKbWDx4vxTBW0AbqOZN2vpZL+trUSBjcOH4Pp6uhIh/
pzfw4cxFiFurl6sajQrVL42vP6j09feBjiU5SewIdVHfgOyQwy+r7KBzmI5ULPcEjGRA6OitGWK8
nX4i6stzmOSmZrH1kfiRIPDPRKHVTzrDjImTQiXqKeW1aDwksKUsDAw3rWTi+1NZRAolNw3OgWUC
Fi9DiDPSm++mRLJyCofIZNCVofbChGQktFrco9gZ510A1HID7i71bCY6O95y9E6KPlJhQY82f1y2
KLlIee9TQzONrraURVcq2csWQVGzR5QlfHFhW15hayoQ9p25GpVJAayED702iKOhGPqC4wk29XdR
Koj/iagg2kiXFOagQOmwSNYW1ngvXQEQRdckw6QIfz0CeiW65Jzhc12J42X4pBC+BxGk8yDI6x8d
FHl/LIMV9/IpIoL8pXLQK8ugnrBkoKnXOcpOI8qeG/i9hvAkD4ZxTzwb6DoB/QALZuJboBoW0Tf4
bQW9CHLeRWhnvuz3pOWfe76IUOw9e0OFgCoxiyxRlKD8Eb7kRiDEAI8mXtWx4tX3TdvftzRBejhC
uLAvH6DKS8qbX84xNsOMRaDFSiPyxrRA/PV8RdZguJT+kPO7OBn0f2WNKYBfJ7pvA3AfalV1/etm
O61SlBxxmOd9Ky6Pu2rfVTbC/WO41Xx4WJNy7rOUQKJfEt7lVZRbQ4nG8+1psjaRUeEmWBTCE/to
4TaCKL90E5jPdg8+1QNX7EsCgYDPIxx+M7ZNiaNiMeKJHAEt2X8XyThpkOkl6/qEZuDV/fwvv9QE
TVvfGChmZ1H0WSuTLukuHm+8wVCNOqQjMbliKIrbcTXby3DuYcV1+peSVfOczPVjOQ8bsLLsQ5Eo
iYTCdApZeiEmYrdKWsBsfPXpG1paBhcHdzbKuzTVNEDGQ1RqtFnHKZ3oCs9OxFWwSomvgRfLKKiS
aGVUO7XzJm4fKkB2WnfgbKMXbtvdG25HSq1W6fed/H7xYVQJT1KrA5R1csR/e+8tN8Dm6+iak2dv
ad1naITyL8cyYHFj+N2f69RLY72AQZo0fAdnKB4Zp7y6efj++Tx/RZ4q6dMP7QkOAPma2hAfiVcM
q0dMGSl8GDLiXEwidgfWeIk7wp5dHr7+gQNPW9mzDSj9WJQv/VIXM5hEG74pF3RynJfOvvn1i2S+
uPtrYYM2YHLvsjOzPbUZB19/11s+/3lG/drs8JCVp02jwXOMBqWZwX7kXHaz+6/0H0LNa8xij3Sf
5uLJ+oaItKUwxz2IM/tRi1K4y739zTPNZFGRsioNV44m5Kio/s7uQ6CLefvN+19rLKlmMjAucSYP
4HiF8JvSMNFG+XjWkMlNQ0q3oTgOHZlkLPCLAukIaFbbsc19kqNWmzKyP4o3aGFMHHeEDHPB3KcQ
kMSQ95wdHr9Lclwwe74JoyENe9Oaol2fn5MrMjIO61iw7saQYt4akG7W6o120ww2An3YxiD7xtfd
VpZSd4kuzLg5wt3ohaWxkWXqR1LExwM/+/ryLc0okmWNpdFVL31VG5pgtGn+dSozBIgehvwvNakF
fP1TgtHWXytArKmGhpc2cii8uU/k7eAZ/jdxQD0AnsxmlH1EJky9lsVFQMuGHnOFIm2szAGsrq1a
5tHoq06pJCbthHpQjd4Iwdvs8+hH5m+1hhJoH+ln5rCb+BizGfM3LCqTAup6d6mF5ACPRSDCQG6Z
idp6zrOOvxhLKvOb0ynGV+YNZ6ymlYcwb+SReSuaxYOe9ypi8lPig9DHgIuJ5yezUMgx1b2ZNXfr
xEEKL28p702lYk5A41YtffYaBZjJb5VetvTe8UBcxeFCPPeDFCVgck1v0Y3RTX+1Gbdz2XGkJEjh
fQn0VxQ/sUhGnZa86+Kn1IDCsHmOKHv9VWDjteeKJdMrK6Mf2NDB4O4n3EvYqlB0BVk1kfyT+pHa
UfbMiRJxToQ1835G9meVALsSc9V6mWCIpuF689ZZv8YQhhMC+wtAExHsV2uzj0f9xVutOZzg4NEZ
7uJAgo0M7tmLgz8XbDu73cD07os+bkC74CQF3hP3xlVfnPS+s01iDNDCeqV1N1kbR9+Zv1WkoKpC
qIx4wAGs6LlYL0JnT8sB5xASfVGb8EcDWZaWdDDPvIGSVjxGcPgerjtrqPt1wik8rFeHR/nkZSIF
7J3cZcHjRLOcMz/YCojeHIFCS3vSj5uw2doQK/VnYO2sr67m3ZkcLtllOBum1Wk4Q3M65+/9SKGF
+v6qWioGh7nwdzrn8I5n52o+AwBb0kdvt2GRI/B+hcDngOSbY9jfOx+kCFpQPFbm+oDRjC7Okh9M
uZQf3ZpmRMdSZW6J/3UqjK/DCylXbu4TwYWr+Sn4I2fn4fwz7hzPWAGZROQeBwlo71nS5FOg/kLo
fCagaRe7bxky+ogkN7MEcpB2ZkitIVnNy21c0aEjLnh4LYaTM++BFsDdkgxTkQ0d8/7a1eraWkbf
GjjlWYElZbtYC+HQ2lv4gYd5vg3a31DZKL7edx2YOWSkjwEpd78zWYTVAsNHwisDHuQABh6ZuFO8
i7sj26P/WUQhYN+342WpYXd7PDsBTYPexaLtGsAMKGD0FxEldHVAN+bpzv8aruJTwcvP7Fq1TkAK
ZMVncnU6WPflvv93C9jk8j1Yv/qLfE977Bl6JjqpncY5Q5fjxEnB7w2srfJB0zLEZOK4v3R1t4dQ
sPhsy7+1zMPohO1QVVSKK0n7maaU3+TRZu/rVA2VoI8w1Bg1nV4jjjbCWvr72IHTQ7OJNfH6iWO5
Dd6hlSnrCwcqAgOfRCdDv4WbXWfZ4gqFLjg8vIQ6I0CX8BsMHWeYUl4xX1mBt8T8vwSX+8NRqtTG
mTIoOrCwECCeVyUGLZr+Ec2dwJDcSrAlqi0E/lnK/o2YalzLSVvyy8i1h86Bi8C0Y/JMqW0ucWsY
4uyz9agASamRYhkZRu25qJxSz8t0Mt0rE33HDgvvu9JjJZM8PRv/ancdPEL41WVDVIy8ScGL6/Qp
8a+52N498teqZTVpxrDF1fteviG0C6qg+Lyc2i0sQH0ch4re+CHyaIDhM/0sPJJitZlwAe42KLrz
q7dxrz8eaAQAoaLtZswr2dIm146L3Wg+6vDqeHe/Sk8qRfw4YoVTqy5hFXXe3+PH5+uKUA7ePHIn
ZXjIQqh+AGaQZdDt9B99lqsX9uFyuv0SRo1h9Ch6NiIGGv/dzZrhjmgI6jdyIDHFJ+I7Xq+WMfff
j3IAKcFG+G6WfYo6FhJ8iLLVWq0XPN11vYbEjoJSUSdSX+kITc2Fin7wSZccfYUXhdEIJkNlnfLb
E2URqFFMooz16xcMNZ8JKIHhYYWQinUKeWzE+a/hc3wDCkJhlmT8V1hkicDyL97s7N664nntDCau
Ga4DjGamq3ilYqiv/tkzKjHQcs9lK7L3UocXUi2K89/9IF8CdVgUq541KfzBlsc0S7OmSEXX8Z3s
8tLyVVBHIDCQAk77eLWFaxyh5ob554Ehq7bl+D4UBjihxlsYa6MYWsGoVp47oHEqG647mIlIlsu2
+GBmEdj7PhtpcnT8+kVE0MJmQfOzBUQ+4G7tEhP+J226P5q1BNg6qhfAj1YB0fkBbNtBseRMJlLA
wDeIwGw4GuKA0QyC/+L3b2/E0mlUVPX0nfvWZIipSx1MK8RVxPg14KC49O0bzNpaz13vbF3pGXxu
uNzqlmDeIv0yAHlxMngJyDWxnRlEtT1dwTNZobMdBRI/1b6a3P4+pwCC8US/IzWIQ9BbDlVZzc14
WYnCEMLva9neL8JM3VV0CTP5+buPHXf0xis/H5p5Lm5mu6eayFThQYLxgOFP3SBb2bzMYvIXgTxg
jEGvhV9AKU1RnCsTBPDCAT8/rZkDN0F1KWELNax3QTzDERbzxoHhUdFr1XTrxWZBK+chGeN5+QJC
8eF18gabdBh8R/DYBt3bnqTg60gCgWNu8Rv1eQB3s6dyG93m4EP77HMEmhgGHL2pgSb6TIBhXXZI
Wg+mtdBqDZ10TkQby80Dn+G0wGYwU8bgh+1J+kJ6D0FUnq9EJ7mgTxiz7VNWkZdgwMJYkVhanTSv
hVQcHVE9k4jz53/TLXinnXPZnXm4MmHrdMbFfAPOkgY3UGGLcvEHFn68Y9D5GLhmHIBi+cUhsjCe
Q8Adr3vTIPGkeyb4JEY1IXa1cLgRxoEXq/LdwgEGHgM50O8JnlaPVC1sU6VDNLCHcFi4MTerimhI
Gr2bnywUBNOnoJtK1hV4hl/faLBiUtt6kdTA5oMx+FSa2CMJyOZEMCAjTrHahGaj60uCgavZnkiT
hhGB7oZZoaxEizTGCPhOi/hFwvzb4JjGzgOAsiBI4SpS0tZFzVhC1OFs3dVwFNZ/V8VlycbA7npS
fBrHFYi4VtF6WMTZkewSnGNDGaG6bESKHVGrUrOzKCalsQz4nbMwlCJ6Nwt5/Vj8P4VLs+nh4qmj
cuh5anytP8KlqLht4aEUf6aKTn+LqxKvMy+IyOjZ7ogdi0YIM91L00XjSugvVSjXrV3zylewiiBx
xv3yP6FoA5g3VOiKgbvmT3/DGytmjfFPnaLDCKcKxSgec1TGlL527xV4QykgRzrRLZkam0SCxvjI
oAj9SiLkBc1gDb79Sos0P+oBkL3w32nkyXPjzsA0/BIZao0YUMsJQWBUM3BsiYYMWttUcw05ICY6
unAmhOQXdTGOJVs60aEdeIXgHD5rRuqVxxdXmzfKAMGsh5mMmcY1D3i7AHQif5oZDbPSn6iYmy+2
r4EXBBj+Jk7MAVmKqnTm7PCl4yhVuNsFAFNhkOJWLCzs+mA24Ie/dxvswhGiyGIyW4Y9ZXt8io8t
O1gifJLQ/wHVaOTMChfRmrJ7nLveL79A/wd81IroivplriEbJL22M9zA2DVAUahwzgrM8vOMpkOs
8Y6qUHUna66lck1RLjo9MK0Dybv9NK+5lQ0xK4nNV25eyKm7e56mIdWX0I2de0PXewxTJQp6Ih7W
piSLG82BexP3jrKY5JeYrJqkHWnyUO+esenw1Ue+Ebn9cjAWbVVbZP3kZiGo2eW2ex2n1RL1l04D
8IPiO21YiUUSHwc7QEJHAB3UN+unOGNsU1F/C8LhHIHM3aCNqxFkQ4Rzc1whqq02/7o/MlY4wQdE
GC/6aDlI+ldDSOzAt/1JEjm6yoWX9ZQGsxNPNBGNq3xASNnL3V1i53ZDB8inSgSdFskTdZ1PHC0N
OJAhsQiz5wb93ItX9hLGoTiRecqP5T3nM1y2wLQ/c6KxB/VfLB+9qgf0YLx9DGT2yqPR006+SwVA
vfnp8WXZ4yP12vRmEn1NR6kBHw+dRs85ZVIgpLUw7GpO8V5TIE68EdU7no11Y/eLky6+9L4pjDoR
WQxiNsCzPUXiT1NswyP1wwYEkR8tVe89bwmjiHIWnkTdDbXSWS1cctDHiixE+nG6jiTTIro4w830
Eizy8qfIL79I50RJKSrUoyWMwMoDc8ZnWqOC5DficO+VfqJ0T3QXHUQnpbzwBgZJh6vNeHpAQhSV
oBaPjmUZ3FZK+VD451dUAUGVHokhY7ghrSmI28QZgq2qsFWvGpGkO3VBkPME61G5x59Oimp0wlFH
X1eomD6GEBUdNEF229TvLydX6hwiqdghcYtDGOvoMUxp+59WkdcPyKEDIpi09wk2I0gvXFFvbW2L
a1wchq5n93X+bQt0r/g4NdPLKVl1LDGEmCm/RP92y1vSsB0pb1UfFYh2YKAhDOrRxRB6DPpzIpJc
/tpaelgVDdsA7j9JOk2BJ09G1GW0hKb8oIXUk1ErXLyhfBu+7CaNbnNhr/eb5ilFMl0f98dekM/Y
XmXOgUKYgI4OJug5czHF0zmQeCuOt/RDdfv5g2KqxetZRC02348KH5tk+2HTwM4AI8UDk6t0ndRT
s9WQdUKsYQ0Ww+w5gLc+fDpu3oSL07VrMEJXFELZm7F6GBxYIAj5LC2iBwPI4+91fyCq4nEye9mA
iG05wj35kSEIkadVlTjNzcW+oaQ+p2j8rVGWRLLh0sCR/yzkoA0Z7ia2UE1piQVrPkeElwpHp7cL
zUyQBzNfyodt+bVib4UsCcGFWIVD+Mu8yQf3Cg8dtBGt02147CqeL072saMMejX3tj3u2MYWLXzs
liTJxaTyUqaTIZ5Y97F2L7QuaLevKUAsWDXvrzTHpwodqvRjxikLa6NP/vihJaT03ieL1QzJyWGM
oHG7m+jSJUYDoNa46esEpbrOelWeQzXU4wNkGmOr6uexaWTUJWXh6hbRxFOlQgkhhred7UrS4CS2
0jsnwLlwrMnQ0C1w6HZCzydLFfenp5ObUsKDd0/jZgQ9pV0HJ17wvnNFxJsMaG30kEvZl5pfHi36
bhRqOm7oMZh5fQfwBmlbovyobMsGdr9cwXmBZGsvr0y6K9WNWf9ZdFgQMJ4D6F8S8uOq923gatoi
cwMtN1PKm8cdjv9OwFLH1oo6U8uAhxK9vW+FxSmY6ZF6SqctccC5WylfjYV+Q26W8isVkygzCRNi
mbQuZ7FnYw/NyYzxOMJLWd7PKzrhB/8oTfMoGV2WLsgRIKhDuvSmuHCmsUScxF3sIHAjjwKQkeuQ
KSy4Eq1NuGuoDAZJxasEyx1Mh5jFWo82HMs6AyRonG18oIXus0yt1UwD5izzE2VpYVfOVz+dHBlR
BpYC1F8uj86/6CtaLWKvGYEMABEEnmf5CGAPhhYyXUPXbqcQxBSb6Bf3noyWOgWN1u3hjIsMHDm+
37YxEA0RJO3jIAC/qPTb32PH6zVFDYUZEcWZnlv6sJeZcuuv/h+80S/3jD/YcJf0ugr3MLleHUC0
hB1H86jMEFk34v1Qz0P3C+piIs7kTY772wHxEHbdMxfDmalkF8R/0XWlKKhIbyQMHN8l42vGtnHy
KojGsKM7R/auConT+Ti3QbdvLhjfRssngNP43DIBgM8IdBBBN6LA5ZuIx+UhOa9/CxmQiLi6zi1V
haXeN7JquO/JysVP8/xoq/sU/AY8Zlzy2/DoVPsiGLjxka2eBjgMRKlxk3UzoDd24wKkqHor/rkn
b3TUMFly9qr4nb9OfXnuLQBOIthSXm5VvDvTqTaDngA7OlZQy7+tSmY7uCvxudnq+XsILTY5OckT
xsty4xyssYt1jzTq8qLfI0lcyc78uRHaHnfOd59+ojezDdAmkC02x8W0m6U+GfIaq9jm44gPaFDn
3/E9AmxdvR+YaorIP9c7adIfRs0vNNeTj4W5821SwtIRp6ocnA2C33lhB0TFKFze2hwzV8fDPANL
SJsTKma5IbCosHUN4v4GApRtBnpAAqDGivcxUp9WzJVTYEqt0P3y6FGeO5Fppq95rWQQ2EC4PwfR
BZ2sckthWEzazwWrJyGs448T41BXNwMJcDyIQYElJsD/Qkpu79YjIiyKl2LIruyaoJSvLbeaCRdH
5kovB/S6RhePQ99zqGMdmL/C+E5EnelFvMDTvP4RFRhothPvHQJ+ekIjYH4Deqid9yNbdCs5Leo3
Z2jdF/xSEwSytMT6qdODCX/7YeCPeXSSIWhkUPx6gA6Jq8LJ6c2EdhSuZdIlaW+9Ay/Xl5+wmvMF
3nuQslnqRFaPrESPWoF5xhny/Wx0OcY1tEb5Yrwa0CpWPJLJxxIrIxENsWqxw4pVPmwRKBLJXd4k
q6wmGy/J3WGt4JqpX/1WLP6OAEtYMv5kAUKEVUwh/W1ULZkboFVH4DZ81B27qq7hsUsLx5uoJLGy
wkFwn3oTkdHMzSSPUUVi0a1ADnUAz0bnbQDzCY4lxKJV3aeVE4+DqQi3HVpZhXfzAq5ZIv3+R7di
OAe+HEiYrPfnnReKtzLtj8LAQFHUaZQGIhNpyLpqFPqpoN1XSGws9X7oPfwA3pzFzcl6JU6wi6Zz
N9qYqXYz+dx3w+49Xla4i5DVr8sl2Tu/Tm9giP0xshOpo2yK0w8/vZRV/TV3j0EqZMPhmBKcOotb
TJ39D1DtAaaLRmIy5WAB7zNbXn0gqGLrA961gecd3Mv14dnp7gwxozyWWPwu074+GPQtxzAlCEJm
F7XloOxiWqYzO3uYRnl3+Bf84+D6PR+PzE4l8FFA9wYv7guBfRnheegbeYCeA/T46ZyjqT2CZLfP
PTofB5OsKRvllgebhSWKdvF/3EhVnvVd2huOhaL93VhshARhHvcV4bnR2NfHKzu8Sb2X/4Ujy3m4
0PkAAbevjRQy9S37BVDmtxTdh4/Vx6QB3xRMsdWJ8SeMWg9ZupdH9vXstjtA0PK71SiqU8ASmyOG
jAkOCAOybbDGff4EXRVNG72fz5dsVZ0dyOUs3dVFWvi/VgBvkK0ggNWQj53ERRYVF0rlcoVlclph
zPNGWdXc7JAzoWTb2zMtK6TnSNMJVQnWkaL9mJsHg2E3wPF5b0qNxDMNYQJD3aahpu/SXghZGBd4
8Gw8MgRmtDFuPQn5VpWbhOw2vboSpi31roQA1vnlmzJFpyAAvrV7QG1IYPjOiOs0tBs2nFFZ3Hhj
I/UTpy53gwoWXnNbXb0vmjmOj0sd7+Zl0cZ5T+KLJbF5q04Z4vhRNqajyHgYT2v0cBjuQTMsxmux
krqSYv70YrVfRL2IGtyH+GrGSqwNwo96KcFbDfRhucqNNUzpL6jkbJQHWi8mCwHiatYOqiqrddnn
4kiYgI2piqsp+cPXGIu6omvLgmmtYuv5WPfnNm7QM2qK3/2qbJ+P62BdzfOtA/cJIr2Ru0aNK3b/
2ax8Z4xALchtqdwHS0kkutFQw2wIYN2KhVTYL+0FmfdVrf3EQ6CPXZwoaqaA63hCpo+urZe2gE52
BaWYR32Nb07hLFfprRbvttx8yzXsBmd7pNsW53GbjJ3K9m7xuMVhi1W9AcmMq423qthCQqQjJj94
0F4+noO2G8DYUbjnkn74P9PXmFr7nyjbQb6UZY57kuYrB/XNALeQV3csDjeIhgiA9g01tgzzQM9P
BoKjapFgo/ogwbPfViMMqcVxBOIRXWfh4kRcnK7Xo3Bw6lN072PEZ4T6KSJZua6WZJazjK3NmFDI
vvDlsU9izN+I8YYv5U+vgd8bjO2mP+SnJLOHdyXGD8+5J+8AvEXDAyJtPmGu9hmw2CdmqWbcLJAW
wlhB8mrXgdK3PJsO0AHN39o2t6ZDGBESArLbyLlk5hfyOlCgNZmgWzuA38q9onQPicnNornyDYdS
JoP0qILdq+wIxhllt8c0WdLYkH/rOxE6FYjNqbfeHClrmCB4i84OPatahlIBfZqvaBX91JQzh79T
ahQ/7FfA8JkNmgEbykEwxOFp2TigIk8Lzol4fh6tBwI4iXnsfqG9anE2MJ7ihRR51KAPfWFmcxB/
BmpSQxYuUt71W/XaCPs9jQdKAXzZRD7UM33BJHh8nFevzf8EfA+bYdcdomD0/HTHopYXN3+rosWs
Ub5efEBtuuUXFCkFP76o3JL7tT/tMULMLdxWgonG2m5Yz/JLfMXbc2ZofOBH6mDyerHe3u3qKPSa
DH4+S2RiOeJpt0qnsFOqV7evaAidz6Hdi/kWeCY409BGvbXX6+WFBe9PmRpYsWDOrYCsf9gTX05S
Ir6kS/3SBaGJRiu3pFxoxmkX6+cN9KccyxQoB6jwDHJYlBP9oVvFTppDkmE5SCvKbYLEs412Hzo3
3kK0KN2Ol9UAWgXDAiX09XUIILcTyAka5y70bLpj/5Eiw79JuiDxB8UVOgFmaVYq3lb8CkbABQFB
o9kTMsMYVR2HlklWEdRECC2+agOmmFj0FxOTf+OFpJHj0Lp96Sxt310ZXA2GX13Mz5vncRVZtWjH
JpVjNDLQvTVvmNOn3Ds2DPRQZ+KRj0yC5wkwSD3PxN16+wXP9ZixxUUxsiilmOe2vE7z+1Gwxg+t
8RpXwf80zBsoZUuZSJToKKSJES/LHDSwcj+Xom2V5Cplj8o57k8ke7G5Zd+YEgRmZ4kpIYA7F4SL
85KTmchSbRgYXDzT4y4/HJYWdTXWC6Hu09m+9xJGdBFZ2BcaBOo/b1XkH2dhmbOm0H3EeCy58NZJ
F8xehFGwf9f/3+GksXNOlqQoEFQn/AWbiyitKTBHYXNLKB8F2HOH1AwW/uAdxFzpTYjoKmVaedy0
qeaiQZBT8unhv+m2RlIjlmtJApjVFhK8fDgxVq+gdMM3VBqwKel6nPZLP5ku+PJt7voAydmXYuW+
tprSgdNgASAk0VeCN3sQCpRoZgcDqURFy4jshTOuDE6+0ZLegSxChP2tAz+TlBW2iJGlWeTWK1Rt
PRB20AzAGdX2Lmniwhi7DRPdM9Qf3lV3Q8qnFcknsZl2sH0SbFla2NKJjN8Uc7PoOiUcn/KDmdyr
hIfGnYAkbySXSh7mR+LSVmQktGigPMcBX5n+lQSURVftzm3p3IhugdmK/BQZTjpb/4zlGClYEFhy
lK6d5ZVoUqA/yYhrUE6YhwPOQNEFONJw92iuQesoLzV8CNyQLRgDwlWctVYHAH/UPkKqft7i4l81
avzgMlZ9heZfdiIXoyk33LR6FFjirgcVu4ToLhwNDKXOJ+lTQk5SaGy5Cd1OOVlNC1rfSah+e/uO
yxowxpsSbpUjzqRLsab+FxyR48j8v1sbs5wNGI575V+l2aIBaWP+nGuvxnuDsWWj4BiAviTdRtNq
v/ExoELR3Z5xAq+wBGgt2/WQ1zZLt0vHFP/hW3lHDYFmda2wVPbdnbq7R5KkRYpbrTllC9RrgrRp
tbnw8QhH4G0TaKkQEwfaFP4EhU4UlDr+azdekagUhQedvS7x8lbISBkIOrG6TF2v9wYHqPvvyvzb
UMWXLNYgCSeJy5KSzdjnlGyoHT7/WX8VABOczNfkr6TtwwW/IsPfJR8ifCmD39rHw2RaWD00t6bZ
l9xTfjg7DOfp3ncGrqB53azhDbhuOHLF2SDHT/kt5ZMOKDR34ok0fWjxGXPtBVliEgXLrfBPGRur
jMfUrOX8gzZGyPPI9lYV+jxe6OCK0iFWSiEaIzm4C2KlbeB9ttJWHdNLPERi/CYyd+6IMAkJ7+mr
tgI8ThLEsyBpALUY/NxKEcYIOGilbyuqfKCs2DrcAewOybJD707/DKB+pqWKpjCcyVbkpAqeifQN
L0yT+nW1pTh3Al1w872ZTylO1lDH/Kz22TQvZ5su2e63l7KxG1EzyFsxre9tIj3nD7mRbcXkrHVd
ZwG7USF/iBQqKnN/9rWXK6XcxWPO3/WmuSZ4IhKLOITKHdgWTMcWvrgy8U0bgKt0URTJ3A8glj0J
rGU3WA4oNJWWcqBbmxofa8zpepb7aysR5Wj0H+aJ2xS4g9Zv4ajAiPH3a/fpBGWwrVB91+Yx7V3O
zlB9tG2ncaGWB30JHnwPaTyEfaaXDUYuZFZCIEz4mh4XmBJsMORARVVy4EkxcsAO2L5YhAKJEsow
nqUHWWkv4q19sXOeW6DgVJI5hXuNdFG2wwu/Me4sodyg/OirJS6PxrcK1MHoDink1ZUGi5Axdm/J
4rp19PBTzm3064igMkwfLryMXgGv/X3uA+7t5+GC8L98P2iJQvjR3nlglsj4NUQCizpVikRQt7ad
lmOgxn78G9UvH2YBTiHlYfQhFMI2IdZknz5hRk+YikQOunrvh3zBYCgkdnpIN3FIGztEACPBTLdN
NBvna7Sb6pELCRUk/yC06cUybPasSc7GQX07icaNW9EFTXuUhMhR85z/egHtWuPIHBjo794sAWcV
t/0kmFke/KWe02uGnbFTrlbTE/YxFZivpyN46D7XrbZL8Q2ZSAeu9u7jCvKR2NXU/i2HGQ15vPkM
HLvCaKjUraD2AjrX5KAn4nUoPKmRfToufFucx1rN+23Z5qI+sNwA9ieXLPn0f074KYpZAHdMr/0N
n90FToBWOQVZiP3o3+vHJjx74/6CptcVhd90gQ1RYN2A5EZ1BTv/rfQK2/1br03FJYWfhRJ3HJjQ
3cg07SJNl11Ej52YZ95kwW57zuKYO5olzU8bTzIl/+OdolxauTxQmZn6rRDvIda3n7Murq8Yc2PE
5piyS05k0YaCWMpKjEIBtqnJxvVDsfcjoYEDboOf1df2U3WgGF6uvZqPbb9ONsrGGRKd3ejCz/ar
mCJEuNu8G6ldUven565DkryUk25WGZTfs3yD696Am0z0jCbE32iXU6XBcBI21qIupGrHySECjC4n
szZTlJE36m4pDaa70+8A4oBISBOKgteZgraSK+lnWbbJ8DWlm1OmdRVP0oivAMn3Q3jqp6l7QiRE
nFkIA4tPKp3UlowAym6K06HDLVNjH/ffi4gHEG5EOH3vn/nvKff/virhE10MHW7SVwcx0ZIZIJop
Ylqe0NePCLuS848/bpX6RpJBHvHSr1Q6zEzcvGLDMf5rXAKmQGEOxvWjzZAqkbqqxYiAl/cScygo
L2wYQmN6fof/qAkm6fRH8lHWgNwKz4pThBHhkMPwjsAAWrES68yPtZZfH5E1bYBbWJL56W/948HD
NGcFYhlh0onVdIey0Laz8yiS21fog7dFsfLMpKX0WLnCMlbmraqhDAc7gPx2RORlzesnWuZjutt1
9lgLl41LquSW8rqZz6SW9aDl0IcNyujULl+uZ5pPY8wyRB7rlAJ0KDXeBMvA2e9SGAc47nIFJAG8
WJSlwIjga8sS48OcIyYHq5BL1WtYRn3CfySnVP9Oe9lfI/rM+xIHqc5HYFJ7H7bZY0jaykkza3KA
XxA85xq7tviJcbxROUB7Gxw0jP1Rs7ojOeGxn0jYk8BQidKWa5fBfKVFO2mLyJ00GsRKSjvF43St
smQSTUgTNe+ac7F3rZud1uWdT7XK3p3qzGUs1eCdsvSjAtuV2kwPPuFJukwokuOe/ExLd+QHlK8p
vLopA2mF8sm6MzSqCotmoVt/oVzLze6lIytMJEoZ/2r+6w+w0v02XZqqseYjFtAodAXwGuGfTQkH
MyKnM73nAcJCZcLPNYlOo2nNLTicKW1ZBzv8L6Rq5iJz1N8tHXe7B/wiD7d8FpKzlHxp5sXrBHse
VJHhK13r8xeudWdRNEhu/Mh1LiSgqU0zGRM9Gqqt5KRFdZaiQlQn/eI3VVpTDESPscPOn95loH67
bIjKoAC0wxqEgfxOrVq2wjP8D3waIDxJLIt+tphF0MYh6W3quZ/ICEMa8XjEsfP+QjGNA50y6CL4
AWIz1DOdJjVaaFGGX9sMda4yA3jqmsp/Iny8BafwwAmFlv51QyEhcKrKq6GiSTQntxctlR5qo5cH
S89jJn9ncqFUJJpBRRAz384VyofeJqnpqFyRyKAKYIpAbjSodvoWArXiPumsMwxlj4NjvEFhxv/e
wjr6XbQgWYBE456zr11Fg1kl4o7aIHEehU9P3pHcgLTkfpPMBZ4ccxa2dOchLP01COyHD3nnSOFz
QN/vsdtIKkWczj6DQFI9kZ5kXzk6V3c33td6s8DlsCi//way3m0G2wIp28S+ZBTiyMvz7jNjtUC0
jjwdb5x3CtEcX8o8rkq+5f5EmyKe8GMtc7bnKRKYRYXs/it0wvfd7m2i9kRxD4Tca1DeTLPagUqd
vm4Zf4oQNI6ikCVSkB8txTIi01ZeL6s+nyjWNGxGEH1kFBeIP3prW679aF9kXNvdGt/C7Ay92uMF
CRVv0gCS7sXiUhU+XzkCeMI7A2atCiJqzwK2GHytMdU9KnJjPreYd51x6MDI7tWTXGPToVqQWIx3
sXRhSe9T7GIXk36KNDXTHDTvAs7irMMHKuxT9vHjbx5i4T89cbFQoauYbdEKsuJJvyok66p/3ukY
h/GCyQ8q2/ix6P7SAZWT54qt25KfU96a8ScqzNVMsT46TBaOUpP97OXGDgPO4ZSL02P/sRjnu/Lq
TYMgQg9i/5YX8tYdrmxCP/GAFptsYXohHTVsT/ygWWGbVVOSfoOniu5N3bhxc86kLdiOO41qjqyA
65VH4LEW5t+wkXQhvUw6pI5IyUgDatgJYU1nYVfij4VPJmGNdcajbdmTRRpj+gJiU2Y/7hNJ9APG
PRiRyaHI2LycbrFbjRNiwNshI5wtl45R82CMH7QyBl2PLNxF+8vbixeSiJKo82kPiS+QLXQPJ4s5
AU8Qs1NvERs7JKNEN9w8Iba9LbIT1tfiQJijOlQ1uZZ/mmoFYSyI4cVyF1JtPqcyV2frjgGzor59
RTbUcDVr8L3lYbI0deDobFbK3cSb08Y2+1iqoVmwhdHMg4+M7d62GJ1IZQfnjXBpN+rNj/WBgLrH
OTZALX8/EIYRgtJ6kQxd1lCiC3InEk4nkvJ2G8IQ+uA5bopIyQ1vtxqNV7NRFDej8CnzbnESCbA+
yiYb0kefa7/VZyecwCr4ieHrhhonMZSJcXYrqzZDtQwEtVV7BM70vITwBp4Ywk1G5VBhhou2YWQa
O8+BgMCi3PECoQU7d/u4u+s7krGWMgkNorIEeFgb3qy+F8vklgYBv8JMYYEgpTZxROuHRmEW9vBU
Wx6VapW6KO8ST8OsxXw0gL4JRJZeIvjDs9okDslodpVsmpBEg6L24f2jZrxyaTKcr34/yCmmjy66
+6fT3RL0SMvrNSsIqb+8GDOahjTD3yI1hhlgT2YeiSm9WKsjmrhzdPfARBmtcHcUmAH4/uCDVsex
1bna2JX1ZbOz4iP3ILyFfb05jdHvbAdbOnfRUCgQf/4Gj/IrFo5HD/IQgbZdM9HZmkffNd5+1Jhx
G0APOr7GX+mgQmHO2nW8Re++0zA9t1scmxx7XFSSXnyxmGqbpQYlJxf/004j967zvYQadQtymaq5
KcRbEorH6QwoHuQzqeircP3KsYB1sLy+PkJ6PiwsfGHHxlK6vd8KxbPnsZs9h9WVVNBX9MytQo6P
SvpiUY4naQt2IwcPiuFc1TmmKHuIwEKIAyOmbPZRmKJEJyZ0c2zRK46nQ+jfa8Rfh4Cjq6aRGOdG
wmcPIA1HkfLKmd6qVnqqBzttWceAerAsqsHSOPo1SDE+3JTwHhYA8nkfEkK7aXCLkOnVGtMH2IC2
2bjaAb6dbkLRbGMtF55S7FO5YlbBlnFLylsZj74ZxHChYYrbA0wbf09fEUUYLBkv1TvaSo7dXpDd
LGCaY+r0zPk3EDIf2SABK+wgHHAVAHIgB/dJ0nUYBPJ1zzhGXvX4/Q0suig9fsZt3brs8UejuNaG
lv38Fl//j0DWq7MiXpilYj6mvoB6TJx01fo0K0Sm5HGMPMsHCF580CdTShD6plWx3xHQgswV+mqC
v3ksQaime7mXXVx0tsWU0Bb5b00bXQBLrpwqF6J4Vtk/Yke/Zq/hjFdwOP4Rw07N/5nuJXd9UbI8
w6xkiFrWuVUi/YK27a7uY9pCCzW+wCj2rcU4yUnyWwUWGbYYC1iK4h5GxiJeDIXHM29AAx2X/tDy
+xUe1wNck5KK3a01XoMGTjU7dNtOrXJPBH7+nSvnm5l8F/QFdFfEjFlYKyCONTZuRdNf41dETLc1
nqItWtBVg9mmSMJKQ+lIDJ8q32Lo2QlezB4RcTI3gBobVOXEkzG/mosoGOjS+DD7l9eSq7gpkvZH
jD9/esew3g+oXGr1RBeaHBfwu7mlfwlWS7zRwhyrD4rp6KJ2o7MM8rTiFxsIk4aJu6WUDHAukWaM
8FyOHB2eoUVvnlhFJ8OIBdfev/VMn3/x+AB/RrCuSGdrXsp9ZaHmuiLy6Atqrf5Gw1pCURGKO+/7
BjoagTn0JiDDoV6l1avHAFweqiFes5fbecWIg+NAxfdD+cl718TgQporSibSq/gAwHqjryA5Y/JD
EzTdEkX+5zO/4LXi7D12/8oYmJzD6unsr798Gnz5+NHxXrc+8APxJ9csk//r6iGlAKb/Jdvl7ZR8
f/ApDbCy5CmKazcBHRXJ41oWxrkRXGzm/0qsFt+thsmUhBlDQN7+cI6dpofwGXqzFnBuflgKRCQE
/mGwNmrgEdm9beP3BeMT2iVaPu1unlPEpnml2YsErJ9M7nPhs+IunNmARyvYgoehEK0FLHPR76kf
jDElr+JEEAeIqUOlqe0ZEvHXMATgEJw7smIj10z7drUzTosxB6OKSTyKGlDSWxrOna/mv7O0VmrS
QmPt/g6KVCoLycMMQ/T0NyGt5Lug7EvvHBpTSqDT8gTOssQwz946L2VX0ZDvwDqCoPt5o1duQKrO
QeM441Q4VAakQXPlLJA9Rw1K3qXm9qPjpWTSKQTvqFBZZG+A/ANyYEv3POJnhqHaJEsuJDGz4fP8
N+LVtyw31c+lJB5KoiI90mdbewkMdROAQQEfdi8E/f+rRLG1c6bP7iFPMFq8bZEKYHAV3ikibbtK
9orttoOaIx7kcOVo5cnCGyA3VJhGctwnhl/t/vhR5Ldr+eO04Apx01YwvlIAPPYiF8xBvmv6Tst1
7quhk+DI+tm9hmcjPR/KM+I8thgNAwhk1Yh0NUVviEVPudcXBA3SaVdRMUCa+BSy5gqODFR/1wuY
jSesWbKlD00/JmpNOymGTn6BHfXAcMB3DLmzUu+Onasque6+9BY2dCAl3ZnC1O49EQu7ZQ/WOfGU
Wj9JBNJ1XQa+XrOoBBMPFEN/JQ/ok6NCCdb5uttWNOZFg914ZZVxDzW8a0KyBkFt370j778cltep
GcuhfS8PsggdETOz2db3j3IkTQXxSqAVDiDh+zF3sGNIKur0Lc0YSBO7cLSQUAFaompYob8wh7O1
VI6CX1YCuBK3EO3NowInis2Ff2QahfL7aO+/jKlNgkUvTVw6GeZftKz4ZDShNGYkRT/2D+SB3r7u
0NGAH5W2ufDxxuqVzzVuBlx7uc8wHbPEyRUSBO1K0aHnK8OGwEuMbazJ6fvxL+O9L2TSm4/8wUZX
bl9QWnpczY3MpDSP5hF73k7TgfBzntLckIAuwjvQpmce+FHtiNS3BXWI5q6Y+GyF96bowweAZst+
qbSJM3PcZn7fuCXIBoCRnOHrWlqmFVz6LPFs/vbNqmwegz+Oc5nMAJxiqfiVF6OttxkasJYf/Din
pEaHBvWZ5iXHkiknq8lpIlm3HRlp1Tvpa64dVxrqI9yvY6+mbJMdh4PlbW/zrEd4esGspLHOoNZH
ebloQwfePQ0GcPAn69MabqyFmkbluTyn3Rt4M7dWmBo3ROXTLXcC0CjCmhkqlCIryzuJLEGAQj+G
1U+iRLwSJlmANv146wAEbHpGAsfMQwnwIY3UNvk0kqFUEFNPZKaFP3mWgTtZFVVXi6ekJsZYiGDQ
UJAWu9UwrPETzcfKPD2gkZUewY0YGKy6kK76L0eAd0g5505dsW9JgclivLF/lOMtv5iKkoiToqbi
p8zeTGSNhNkXDjF/OxB9pVK2/0tlmt5IipNciYrAvlPv+BKioJEGEF2XwkC2QVOY7KoRfuhbr2zF
R9q7hBxVvlYkjITRMqBTh1drWvz2CLJEgAVDc1aT0FbdkNOza0jKtjY1m1HmhM7IfvMO8DNayzGN
GFOEuF66fX+d9ddenUA/NYWuIHnp9oOMRBAAWIhEEREruib4Uji5+5RS8P3MmjR8ZE6Bd047M27U
2ET8QIULnl6q2SWoamlBqQei3WSgGLtqEoIaa7F36NbbGNhiCJns1oWR3IP4TPIN0Bj995NRNM0j
sMbVDrXt6ToJnzYR73A2ctyPnrSbcEfG+anbH94nJYCvkRikd+ba8J/XJ9EZr8aRppzaPFT5R0q9
aLs04fGWTc2ICNPWky1o4Jj5bjEwQNzfVrx+eB7eOtCiHAl6wpWRAH0EZgK9DtCeqqUmePy3qBLL
+KDlTG1SHOpdrVY2dQpc4qg5KO2cyEn+H7gQGzAjpcZeSZFvz0pdmd+IhSEX/k/WE6ACABO8mzUq
uWfXGLO+83QrPlt+y11+wFVHqvisiRDauL9zdYtAu6dBUBgXmJeY2PCy89uLYEv5GqALhZt1HWr7
cD85puRaUBcBFfo3IwtFk0A9j/gT664cLoGQh4Rge1PgXTNMIdRoqDvzm2aV5b2Ns7RLx8+0tJKs
TLB1j9gP9hQxOf/koaFpJp68iuh02jjvf+GM14JVJLEj8Yr1tnbQjafZTQzIfA4lw7GFCUg2oGSX
fgeqkD/eG21yEXAZQGFx/sLoLT48wweK5n/wWhHSWZfLuENr3Enl+066Od24vpB0SOtoafjY57wl
SDt0JbzpKNg0atyZKK0ZKTG3YTo4qUVSsT7SLFyTYKuk0p9fmi6VpuWNW45aYF7Dg2zih60q4I2X
g27CsxTgmRFMD7mlWJ8tWlvqmpjJ2KTm0kE4p5dl0pfRitbJkpAboeysGky9f9SKu9toCYnd7WlG
Xyx0KpmmPL2GtvTC1Hpt/vILgb7DkBfYhtWrSYCp9TQYRS0HD7GDoxw3Bu6xtSII8OwAbjeimpjx
zROhk4mZm7ISMbYWQ/ZoZDQ67u0ck2sAKFDtBqTXm0dP9F1i/Z8pz5eeI5/H4o/bLZhsxM7N5HLz
rGn1pJvFOCVTIJ6Z6PzPn/+h3I6gL4GiPY0COjVtkE8Kacv95VVADBMjOEbxsq/A29cwBgfuxV1E
jnxBQq2J1C4zHg8qvVsL+lyXOcA9LPkkrCvLFwsdv1WCA7IixBkmGLZg10fBgEBmUrGlNzSyLcJB
1eec83P3PAb06Jaep+fvKSLJ5QKGo6o3E8qR1xr1+QNYA1bwlUxid89JXf2A3k+ixXBsfLn+1kxx
miQXZOhxLSqwxYOlwzki8JhCQ1Qb6YziMxeW3KoCnNdDA1ZjlhNf597xE2hSqAAVC9aSD7X/esrm
D/o0YfS472YPbhDudY1F2DqDfcDLe9RuJ4EeQDYO5cGhkOPJzV2UmcMfDn6Y+Y2nyzBsl+W34WmR
FTFUxCqcFTq0G1f84349ryQgQl/ciLVpGFwNOdtBa0VUAZvo/NaSiOTcVnq4uFXZ1g4I1y10H+jr
EglPfrgZQ0KR5nOOsNrcI28bAZO0z/hqmYsXrGAajvruXNCR7k1b17YaPE4ZrhdTgcqUBQN7UJMQ
gO8sJM9A2cJcRM4dsFvoZ6YW7PFPMsyf8QKcC5/xH3TZgSDUmAaz58K8aYmRP5ajqT+l9QNtpLXz
HDOK7HukbX/fm8KnJExBc7rAshUyWqDOUrr3A1DzgvhjY9VnHh35p9/P1FBpdvHHjOKilCjma4eN
GnUnsOlbGQqlSXMvCqD0fro4MpwsNr2CI7tzRyMaKfeYYlMcc2WESJnCeMdjejUTv1qC8Dgq12x2
K6rm600keL0Q3ZLPyL5EzBE0w8LYTD+oS2HnrUfuOdJyBOWO+++SeK3CL6o1bThdQu1iMqAg6Pjh
4jVyLtD4zFUbKUvt+aY58TmLj/q14KWNoe+4WPUctV4ezblmWD8PAY3PtcchSPmOp3nXt2LSmtON
i0E+KQ3r97S3CDHljUHYMD17e/C52CHkkTXPgyHV/wULFsT9ct+ig9wMz8FdRkPODwXyuvfvqFM+
ew6PEYKaIEiAwKsUBZquEaGgjvyVpTnZgWGwmgK+niwJ7bz7IQ/4Uk+M1wUfTtmta8Pwnpg7V9Ao
C9PJzpEUNwsRj5/75O+ud6icwBr4rO3Gwdsl6dnn9SJaXZKGOqx7kr/q4/27akkPKydRvsVfzPux
k/R0ka698jyiXg/XFObl3tPh9Mh4lMMmuUs8TDpYtCTGRFDLDD/3JpoETkEDVxY2dtLfYTAJWySq
JJp2h5Yn0u3+5JJO5hv5fJbQwqckRu3BsTiqnro0ToLX5YMI6zHM6B6UkYZFFXkT9rrH1sCBppQq
TA46ksVBNz8YgrUfF0qQiQGZtRJ4qBAXHgwW5i9dReGGxUl0J//7XFsETsidxL4+FgilYVfDQz0L
memQPtrpmmDROOvGvbGVvik8DYuFnHDoczf4xkH+o8HgFvPcld9X2i7bxdmGXqfvgCxvwe4xC24n
iP/wwt0Lp4eEVg5lPml9AWdBt5uTh4AVQ1kuzeR2o4CDFDj3pDgCT4uMMk7M1g6iJRBusLs4YsA7
FMheV1AG+9TDAKoJz1DJde/CsSSqb6aDpYeVYY32PL52yzgAvZMnttJO7U9AARNU0WxrbY02q/r6
zUZJqjjigz533XKEyL9tP0DXeI0vGxJzmGNVlx4KA86k93LvtC3Ts29bLlLOW+mwhLOE8ua4lsZt
C+io8oCT1nBgQI2ob9CuM8HxtPcAgMCg54AXGbW/zc01fjtU1j42QRIYXIxL1K4j2NkThEa7Wniy
E7lcpXE7UNGSprGVoEQUUh7O3JRQx3KMgJacB5/tZlfesHzu8JZOrEIJr8eKEzKZRZ+T428kq26B
n0iL6PmOvPLl/VxGNzCvpOtPaPYT+DA8kTJbsk56Nb7X900MbQlmx7E2vWXz+U+8wHSLY5cHhvc8
2ZoBOA50TXxz1TFe8o/0tG3D4gkD85Ne7l/txys8b1z/OoSpApus/fcj4YrQpi5WO2BrLGW5NgED
6awMEp1TXsVeD79D86TUSne2QSomcD2PcaRHqrc5U70DFvs4TxQFjZYJrRPzJBnY9IpXVMDiV4aL
QhxGpqBV57KNXTvimcfk3V9LtPv/cEfboDahRyJv6im/8N71VPy4uG1liomlxu15nIuF3ouJ53bz
z6nbDhHQuwWB0AcABPmBSs1sg0oVbbzgrOI6xy17yJEob6ZaKMXzQqKgnaQPfDNa6GtCc16mkGUY
Qx2GlrbpnsPq11m7ZSKrCfsn2wTg1Iys3EfcvMJn4S8zrPIqptXlEHLbGbyOqRiFD8pGDlSPHd4f
KKEDclC1qbMN0E9RxvgF3dD6+J0Hxu7MFbp8lapfpr9yQaly/KB4DYjJ0V7Yx67KPa61oIkNWY/G
w2q4d6JU0XkvEEQTCmoEITrVPyakparkib8LP5Fa09Yvaae44ykOXdRC+SPCQSdabvsNQCwVDAtO
Yxxs+/H3R708IFlvsqzRxiO4CW65OFVzastg3Lo6b50+MEt0Ql1iW1g+cMB+Sa08JmL2qifWFYn3
Y8T4MM5xDkNGYeOCh3r9dPiTfgXe7UsJ89P1LG3Kvajk44rgaagOQD23v+QB1BuaEKWDc+bBO+fw
BQhUyru0pKIlSdapgnOc830QAYF+rY5XpNZ68+lv7RRtHzeBB2BZhPp+8ZAzvvz5ITZoXLEFgOF3
Wnrt0yGmjVkEUWpN62ghA0TR2qj8iQUqnmoRGUhMxOfniIS9WHs//HyoPFYNzC/JpbZqEsSFw3qp
9XlwkGVyygORa0Zxb3M+H7KZ2STjgTQo0M9jCDKKdquLi5J1RdhcBGzy1K/TRkPqTbeNKLAE190F
S7oV6hh5HxAMcfMB4f7BvG/bzIvjPvM93RKVb9CzPFi8b6NjwF2uKd13s/G4R5bJ9eKE3Bucl2Ms
esKIJJ4fq4pLs9qBFLRRKEBvk9czupED2CldOYgTcUBlaDpqRlvOUT4m5YUTp2b8ywx34YmmxycS
xtwJ0ULZm64W3LdtQR1/Wu/zgZWCZJh3kDa4ITSMjXhZojIubuoeCa5dU1fVLDBUXFgY0rOwCuMM
A+8hCpdeKEzacBpwotGcmIanNS+UMusXL4q4bvFmxpmUosl81/S6YcdZP+uK5JLeLqkLXIYU+kNE
3GJGxKXcYB8UD9XzCqLAkr9wgIPUjpeiv8kgiZr8sUJaYgF2FtFr7h0PBr9tUEiaylgUoMUnoejb
8aaEWOW8xU2QEd0KROnbW0Ty5PlW9P2Rcl1JZsSKaCaH8Xl8Ki1VOSmKjWEcZqfSbbAnx9yKm9Q5
2Z9AWwIu5VSfm8SeBQKi5W8BOhbYAQ9kEDrMbNiI5rhnbmMANSXcvNa5tYJEW+fSvBO+HDZn6BbI
ptzDVidIrwIOogE4FQqS9rK467ftRiiOsXX1ah0hTjB0rCWtokOB9RWlKj2RqytXGJtRSzilR7AW
8+96lBJyPJajSOaERuKudTTB2p9qq392Tkyoy8Vxc/rxOBGv5SmSfZPIGfkBf9o0cKhPFL3xDpql
H6W6kLbMfyOVbk3rEdbQ6yrkTqA3bTBMiSVriP5zbqCPaHkmSEdSZADtVY+7OZoJQBSSYipByfmv
3ZiA2VekWPeJeYJM1/D7jrTkaUPh1jDXoG3N90z8xce+n1uyGh78zujqYgGaUhi34ECK1PNdoQdk
4gLztxSjdm370Ms9pim08raj2XHq+Nlx2fQrZ6Qy3nxR+fErvnHomJ4uGC/ZVXL5Xcs7XH5SGZna
LVAz/TNUcAwicyTvz4KzFNvptGuj3hFMN1LfSBZPFeXyukE6mgLKqdZTVRmRAB2S2tIswCdsISjm
nsN3rGVm0iuR6fm0IxgFs7a0yyI5Wn8qNuVWYqlXeCkMBBJTpQTwsc98qMNlcH7EnarNSVBX5d0N
OKiD5tA3uL8JaS5QLxYCar49YPaV8VRSEsWDbhmggCpmN9oua6jw5ynxZCaCpEPTJ5RFjz4gKIA2
IwK9CbuAbDc7sHStU3HtFLKLZig/V8pKJqJ8g3I4ZvYtBEUph6gY2cUih2oKoKRhYdfB55hqLC9r
leg2NpBC/DHmDswJ8y6nHDj/g6Ch0PK9YB/ahZAABWy3nj1J32dChSVZ2dqLQYUt0NiKjKFWNcCA
uV80eJehpIWBHtGSaQp5MGMcuj5T6O2iX7kdAehYO5EuX6YNPy0V+rB6KLU7UxE4eNJSIi24NqWM
r1xVp/2tM3B/s2EiDSOf2LI7qTkerf9Ikisw8kQ5/KwkAmr83i/K3I8FzIpWenR059XtfiOzYgYI
Xsal8txUFK6YXywz1HEflt0L3xbiZ2hhSEDfG9WhsV155k4SovqfZhr+G4vPXFGi4vTZVrhkUuOC
8FxnMeL4+QowELxIbIjkgw6EwbYepGOOpvOATOs+sKL5kMfy1or8C0CKMi1ef7gMLizQMJ+23a9l
JLKrNWQkOGhYL2t2byerHck9uV/etIyI14hIpNcfPi9EgpxCO5h0gUQJfIf4F7hV54HnjWmnvDbj
v/IRM9esG4SB/CaI60W96haq5NRDGev7wxKZol+WTOK/OHuYIkvEYVPsrBDg30XSNRZLG97ghr35
jP6FTSC+VoIdEMuGulNOrFETPZiXMj6bjQgrg3cTVifm6jDPwtUFziDAlovcEDLnf/YGCSU6Omz4
l3uwA8G17tV72iQl8JjJH8N8FgXdt8X6gBk2RtrUOASuc0XvBZrgK3zJdP3BI+nGE5B5NZZM4ve0
C9oZLLJBpRmm2FusKFvQETWsoyKRIDzTR6z+EBIfo4bp+AxDASAtMx7dGzOL3N6Ayjn21jc9p3Ou
hSqAQiu1lgJLFw9b3ZO8UAXAn4JByT3Xm70dxAgUM6DAyJVQSDOjZpU6lJbOn+qKFvDSLViQGDjj
DPil2Vxuo7iO7PpuhXvni2QgcfYzcYQc8Wh5OlSILrD8ttQcebVq+6c/sjaGjT4WMYJdZPeEqv0W
FUrhQcVDGMUNJfU+OZe1P+8S8ZbBMQDM25tu4CWo0/a7rotsJYYHOqaBi217Rg6Vs6R0jpT3qLKs
4QGIdmknzuUuus5J7KaOaCsgFvd7868w5qxgM4W8eOKa99EBOcOHJ+ixEzARKFKNoxYvVyWzyLmo
OHEv4NE64VbO4znYf66pTCpMYNLTgv2Cs60WVSwBksdTRtJzIub4Hi99bMVSu1Vvv7BI9QbDx4Jt
K0o3SJydXLxKFylksqWVvGylK7T8ct4OgTY1JoQsQoQ7HD0ZuJRcC4W7cYV+sXf89HrMy478vNZ4
I7U1W1zDi3PcVb6ZkTbtoB26L14UNKSyzPb8ek0w4HR15KUj/kUmw86sfYvx83a6y0iXUUrBSQsp
JrBx7IjK9aGYzOr8pecfMvECjDLVFNYBZiRYtBq2YUDmvwI2AUNmEgD3rWfa46vA8IEQDrJQbC/5
QcMN97ydjO0PhBB/lHcaWoAXToH+b092vc91HpWXzrQKj6e587bid/SXhvGLEfOt8j9oKVsH66gD
gSqDLS6S8bjKOskvfdGDb3nxPe/21RyFcoVk9ej1GfhII/H1G/nGihGjBZbW9VSSffiADPPpsnCq
2ZZ76uXel0exFSj7304R0etkV6Y89die6f9UJLfsWKyKme2WRZzryTlEypaior1SME0pXkfSuB25
akLLESFcivafQpQmsoDzkt4AlmTdBjVhhvqtZ4v+mjMRE6pN3zv36ClJj6jvAkH6mUf2BOhoauDL
fK0QzeO4/CApStT06kIdV1CBl0UjXWsfw16TSbXbuMS7N6AN97VkZhenFw9dG76NzebHhTQ5dZdE
DZDFcMI2/4ApkMuS6cuFHLvPbIKVuA2D7E52mKq0jml3iz9b2zqzS5H73sqv9hPnQulq9iiZPzDI
nHFLUXsBoG7aMicUC5K0QKFeMd7BP812ZOilQ9hnGFiuPKP+qCktCZvlMmDjmz5APkwOCKSDMh+i
IOKDN1/s1V9eK6UezGhfiaZeiUTGVCdnGJTXFTMTC1wjgodqU3sQ327Xxd0cf0AoROdBbu+oOUYl
Ywu/urioJ2EYFI/rv3AJF7mALDdOT4lKBmp3UGmZUz6geRgAtySsUhdl5YAwXg/Sl/Fye7sSikEd
JnJ5OTFvi5fDKXopFfD9IYi6l1UT9hMDwYu7KnMf8sSsR4WrLCr/Qh5Y2+WzB/EO5MlTPJ46H+sy
x8g8uQKJvEjlqoR8gKvfx281BBo1wHEObABwg1dmUSNztnqpI4kXvXORz+KbLt+R5tKXGDkPBhxN
RI2NOasKkTSQn7AKpJHQmIdQy7tOzVvpMtYiXpkAJJ6YT8+bE+HF9jQMBXWWXBl3wMAsDqbsXWN4
2iQsvufhu9SAttDNrzWQjGlFHRrv4TzzrWPQ6RSxZZ+pabzZUp/JmMCTlDfU3WKwGUMQPAek0v4N
+rCTxv5jea51nNZ4kWUK2iDM1F4vXOUbcObQUCsp+ipAYS21MiqUfixhkyHtUCZA61JV2gStbJ8Y
jgcdFWxUoTuBZUdJWyLqn0zG8ZOViCx+Z+/Ktf//nN61EW12yuXAr/Ky87rf9+rE9IYHOeTqrQPM
qSSSdy4vlIHDhm3oPluY3kGZbKqROXOcnKBVXNAYBxsDSxDnzOtNPEwqAP5xBxZ2Vwz4J4mhcNxE
XUadFj7qEdcL9mb/UvKRWo4Ur4n1OkaBGQXPg2NXZhttLcWXe4Qhzho+oYASEMQVQK9dKDj3tUHq
YhbKmWYtQCLpQsXDXUkAsHekR2CjvNkvQAQ1x9XrpLZLqZMFE5rsST4FL8+YHf5ws6ITjrNlxdDp
OuQMh4pK4V5dXnc0zo+ut+mg1Gw/F72ra4flHkpgAnj2q9NR1+ZQJvlfevV276nx1dOK5vggHsQk
8EfveO/DJeW88yxIOYH81NaXiuof4yrDIHuIaYJF22epTD4eZ23qMkKwtsndBM9HirSAD3poCXiT
O/RVBf76BnUQMttD5MkT1Vo7iizqlylGBCdXY3Lt0yoq4hVGSlGYD/6G7AvEqeE6rcPe8c+1mmOK
DGtDXsk4u8ISK7GeiiGCfa7d+IS9LV/mYLrHcU1f8AayUXh5zUQCe4zJ78gA3qzRCb/aTmd534cQ
kNksfgnpvLuTcgMnMSzk6Z+aMpi9l3MX2du3E6862O0aQq3OnoX84PgwtstbAFRgmOf3KYEWJxEe
XMS5xmu7/uGbKHYH/57xWAMr1RjXmVryde/o4/8Np2EDIR+JWO2IGHKeWY573UNBALEo3y3J8Oud
fp+98qUfSi33jpKj+ttr6LYDfLvwHoDd3PssbMy3W5MhrfdOZ0R3ZAnGuZd4dL3XN4MUOVYtlIkr
IgHO8UpspX4UTREjYF8TLr3Kzvf4owaiVh4WOWrTkuFqq+9ZVrYH9o5dl6liOiun3Ypwrtt8fTOl
TYNz4LIOKTyUqSI67SvjmZwwVraQAlafhKsUirueSl4GPcExsVw8uEcoou1OByN+0mCMTNE72JdA
HKj8CuG+/tyyFBzOpuy1VmjFhvSafBPHe/8m1rmFy029GlisAybwdMa9dFy9vo2iFY6sKQakfhEm
DAO1AJA02R/toDG5MGVoepE5Kg9FoIelhYrvOY246ET0LdBKdE6rbsx7BbTxYQuwoGXw/7zO1Znu
nyyKS42cEZkpXkP07QbWHkh6GPR3k/rrGEvDdPszW7Ovxo4oOKQeBpOb/TGduPYBu8olOfq8wlmF
BhFVeqs0knSwwFziUzjhr0QMWJ06/5Yt+N6MJtuoXVOFTVLwtYD1EbVoMsfajZpDFKsQ/Y6KgfWi
AFtBjL6eNaZlQOJQDjtaY9QLy0HgeLpmmNAtnD0nJDSRlZdiqNN6Xo4OBBCQLDdswyZuGXxqj++T
oCs5AIs+frnP/ILkoEghhDLBJhbOiGUjcoGAsxC5R6dFlNqHvQBd7WHiI5jor2KrBJw1lVt+LXL0
agRnyfRH0xA2hjbW1NDYMmei9N7rsq3TJV1/DKQGYiDPGfCZZ9r3eXFdLi60l9SrKQOXq8HDRA2c
XhXUgHLTjiB/yncOKcmCmtWE+Z1bwwZr5kmiTNvMZuC/2JJ6Jxy3JTtIWGFIdgUrraiWqpHPHRj/
gUP8SiZE/+JpsTcgvukKQ+bvlJsbVGbBH+A8KBjJ5WGT6qQTUMPe5Wdal1PeHargPNyB+IPpxBP2
7gFnTThSfeyRyfPWg0waoAjPVhTVP1sEbtx+/64Oitm7mmFYPBWhmlYPgKCJsB9vsthExovZJ4lj
qHwwLiascMUTzl4xnh7J5DpHegKKobJJ/cy5w/X7tuQCE0QE+qzspUuDKkR2Q9mhuYERl4b9XaI0
GPq+y/fod//Wk0IlpEf+7G4ZV1BROJozb6T55BLt8vZT+6YWPfcbdoWUUnALfh00goB3dUVXtu5l
7uVwyDFvE+6ucQixjKZEFlLNCyk+IhK0iQt+7LPIo+5LePVWTSwtHtQboppC6wQuMcwpJAXL5J/7
8Ujy6nSoyvMrhhaPwbsb4gsXyB+fBhlIBFoXdzdxxf47ENJvJ4bTsH3HmepUyxmWiiYrEbMwjRKn
O0DhnUGVLYleEEduQDsTUn2eYvMpRR9KNJao4uNtsqi5t7C/TRK5ohk/sT+QQuDCQZqXzf/wIx/S
c+n0qPswH+ONiR67m9F2RDoH6++SkZP+Fe2o1a49Su1fuQsHtSi5OyG1M7r/bJAIL+6L0BM669Uu
RgjFUdPup6mlBNYRFsMSxDh10WuWYatJjHsi4oxzdrqSJTN66b4I9hnZ19lAvcQ5YCU3aMR4Rypm
2jnXR+rAONl17bRfCcYK4BYKqLRjB7Yj6HNA7d0R5yiQCfgzGxMKMpoiA/BkGwul/0uw+0/k/auK
dbahbSoELeLS/LWHWxhYXwVSc5CxX3lHuNvw/jHlNtx3hvIXwGJM1XTI6cfa3gM0N2rOepwUkWw+
QA00PoUqLntaBOqdc+8PeDKAhp010ipXG1IZCDj7mycgP/0gBfhr35AkyU+X0G80U1pWQ2iEdyES
aFK/HL4cRfyj62/fYbOd5NNngR8ciwjqPa8GtaLyJIRgmQDCfXCeAAM1Nxj2vXMoSkMMZLOwnIOb
72vWrF0TZGsDDuOer4gxh13EvXXunFRhRQhbAcAmVQgrYaRkYks8Thk+j2DBfwBkn9XnGrdxis7v
Z5KzHZt5tnhybFXCypVF7dmgA0xLdyMKX/zSBnkjMKqTvtMShkG6AuaCj8jogzMClCbHBYc78lQG
BUlU314lWEM9IRQRM8NMThXA8gSqvuIWKI9N7K47nCuWajLieR/9umg4IhLaFZ/syee9l8KxpO00
EolWZ63LAHSivmCN21V83gIoRPIg7VSIqcD60HtXPTPHbhTJQlkvHiHiRvlSqD8gtOBHQ+6yjyWa
dP5Ws4uEIWA593+dHuUL0YNSXkdj6G8NMFh2nLVJ16OrwmZIJsUwacs8nCupHraNt5gGbK/Fbern
C68Twkaa9fev6Ui58gAo+AmSNuQZQfGm02Hv+e/zrrjeTOEAxlTNYFEaE7ucnPERK+EHcBE91+WH
qZuJZ2Tjk7ogGMoX/nGCY/F8+n8ZNEqdB1bn5J+z6ir4mE7QZJIG/v/3l9wpQaYvp4AVT3LLKiNq
iThJAE5IiBB+yoNT58u9xsraDw8BRFfO7/N1arB1cgJHSX98wr9hzWaXfk6B3IfW746Ho0HiLG02
QC+DVKhNl0diRTQdq1n8b/FT0Unp/RVyAL2Gi7TCXQF/3vKtPemNmAh7YNV1E1a5P5uLWsXNw4Ae
WEdiu2cTu2Jstud1tcb83o6L2THrZSLt2yJU6zop2Lk4vgGIq5CvnMAgUrRjzUVEmYLS+BWm5plC
GAj1DlSUse7C4+FbCqRcW4K9y99RjRqbZ7xKs4fj66ruwtcAUunyaWL7NZmgeknjHJx4H0ZvX9PB
BwBKpzyiLEXPzg8vPkxJFdv9YXH4syVEJtwyzgp+98MABdYK1Bn4WoD4RUQWWW4mIYNwlEsEOtj/
iaLzMw0A8fhZ/3o7bswCHml/b4JFtscrjjG+bW9EHBZgmXR70SKcDaSIFZ4gcIoOXqL82uEtnUa1
JNnjJWX6UxNXrPG2OU9hZcYyCH5eQxM4AY1Y/5/OT8Jy+uXKwKpCTuAnpaBDclUj+s4A476UPNqk
c0wOQs2CKX2r3QFeQzIvrMwi1G537GJr9yEVRvsuvmne9YFqoX1aWIM3r30VOHFQqfAAZYZrURij
wUpazlYD6spy1EKPjvdQnA2b/rw3ckZKuEao3oXKLGm/UfMUvdx2BsFesrzWqlo1uJVNakh3u6RP
8cywEzi/BZwqU6s63T5epnPKrvn2NHQkP5SYfdOC7Jrd7fLe/XtMHs8giY98ot6RiqJ36dECd6Eu
ua5x9ERNNUSNHLiAuThRC2XEK+ts4tEetkgtYBJ1l58S0x7XKOfhbmdrGZ0jTYoqOyhosvRcnjUv
QGcBcWeznBinTxp7W5XdoSefJKmyrHZHaKzon+OEt5b+N7OC7NcgaCHV7NZrLJVD1nUWQhhMfQWo
3lYuB55TrylhuOK2kNUxriSbE3+ftKs8DAgxmgW8AY5/mTttgnbpjVgc9MKzGenYNsAKnHcPl4G1
btIUXMDh76l3q1BX+e3JWSTokfDF45es/iZzUSsrBZHuFf3NT2YiqSCOWjz6CXNp076yVRy1rXe3
C8NQTV9liG2fVN7NacmZdEjJcQ3LSvLCiNsBv32YB361Qtq16x5As0jDFJKYDDF/4SgBvOyCq2pZ
FTvO65B1IvqJFeOflRiI6uoYOpkDmHuDBypvcHJQggWNQ/1rPuh6+DdxWnIdwuqI25+W6w30OlXh
jToA1Zvud5dvIRfOueUfBkSAHXOzCjMIdNIQtfHSIhkc9fq9JtAtiTdtp2IcpkT+Otba2yP75024
lEc7yL+pMjKPIchsy8ZpUYRVs3lx6GoSyndH1oXTtbHNXV1nyG74jEczkPh47yjNsVL65P8nrfs5
KefNjlKEpm2cPO8WpFmV8hTccrWsROko6PNf+0SVjPrFE5EyNTtNETJNFB+TA43lgAlYDL8hM0u5
jn556AkeN1l2ofha/9nmrhBoRSpLTEzi3b+dTx6hkSNGkahFSseUcOJBsFQ0JwuGbO/YwjVcizE+
yEL0ZlVhBwjygkUFLg/6EnjqoPHmdnzBFCTPzD5DUpDZX/2xfLudFHCLgHsD/BAWroL60Vz8Eu0G
kolpAFM5sc2vjkhAUzij9JtqpoAGQkL2SLTs4TGKwwGkKZfylMapdgnO0U9wl4io4U1rR7DvPa3D
9mR0Xpd7pyNC7ZC3SQFdNKFlAurKiPobU6dzf/tv5hu4yCUQY2nZElnC9WeyNAK4U9wH/juUuc26
yi8SEuUXlxW62LfVYwl3RV5+RaLyd3QAa25oWQ4VVXYEI/37NuSZWiPKLQT8nf9Q5QO1+i0z5ydz
Qor0jZq+yb2gcg3urVbf5kqyKYGZHgjmx7KXXIJIsk3rP+yS+aLZgqiH1GsEEbnzoTKZc/7Ocmza
/ArvsuS3Un3SGhpn+vYFZltY9K/U+iU7v4cAIlgyCFCkiBQueUZpVzi2iUzoSmywm5DYbnwHtJL/
Lr/mZf8V6Zr1zgpX8NuqpR7dmMd0/i+ybUPS7VpxfMKeh+dDpZC3gZjumg8J+RowPGDnOSJQiukB
MtYAGgbl2CQwaBM8T29kTHd4BT4poPiUFrsLBshnExl1QQf0Ax5yrE/4//svam2/vg/2jX0mue+A
EmShCWc5gvLMLSihUoUsvNqd13aLtxLt+NgWia9BbQDsmj2dOq6uLBoQDP2SkjOC7VWrm9RFUWxR
UdvpfGb6SioiGgmPnXKiOyTILJLdPXUgac9tAdmZvnfWVkzB1WCNC8lFW1oesBay8mZ2jRs10SZ6
UgzPGJ2UwhqT9/F23x7RVVL0wesigBxY+XuIU5LG0Dxi2b87AnQ5zl//zup/XSRohhKv+ZoOCyqm
2o3notonbE4zKLwTIeJO+CACtkMYARphHEPnXRr86GwvXdhC08HP1oSxiFvzDllgsd5t0IF3osYx
veu4fl6k3LCWHvkdRo7TcEY4xoadQudl4HHJMh+AJ9o6vdByA+gsUKr1zG95qldLiNVcGYSdpsLZ
XHoH2p+Q7ciQOgV6xtRuTb3WMMOyMdzwbAZAuAd6oCxe1glNYBtiC0quFeXVu1zHncFImCSHEGSM
t2yLyLis5WVFHzJGMZVIklUwIVhOPP5Z0X1oKYryG+tkxuKMiU6caDESnBB6KXvHUObB0M72XlAl
Uz6D7mlvHTf0/1wfL7s4Lnx9VJJopzSyML4/DiVsABNXD9oN0mfkWkI64/Emb5rJFBZkL+lZ3iBp
ELD7i2JlfIn0gHFmmIYE7tx+TiCNUum/T/fb7+oIza7eCR+TxKj9acp8uKIF0TmYHRmrgjzJhGX1
sUCyiepxs3O1yxywWI9gqc0RmJrFR+RhnRPqkvwr+Hik/SVIrTQx8Sa7hTeBc7m0SaHezU3aHpHN
d7QbJZWrEc18NIqt5A8eydyInqG8DkBOTpUogoKOu9xxfDT+u8ZcPy7WIZp5E5mYQtfoaUaPdnzE
hPSeQeaUoL3bbnALGf056P3iqVR/KiSXmdFkU7PkBXy7/BUQTDWX4QXBxbMSSEzVYzntGI3A9rK0
Pc8jeSgW/XmSfmF5AG2TwnNlWGj9IJgWLlAjYEKBzPmCkV/IxZL0svePKtdNjxOYvI32TwhFOFR0
h4qHX+XJxmgKqlW2WlJnmmDJVQfYchl0WEzOMzkVhqgK65f0JVL1jOWXOdbr0n3lldpGxvq/pK5H
X/iZK23Kp1V4OSYq6yjWzNWvPDrsrhktLj87PPxK96Q89pms7+8PRDJN5mUmd3IwRgwzHb8Wp+IV
xgh4QdmbxRRHPgkDd13Z4AzZdm+wqLlVbUk+Ed2d9shMiKGJyDofeMmLBRw94Ipl/S8/uiqZIPcg
3x94bUWlmRQfto84/LXYwU8PW1W1jces5Xm4fyMrgzdjU7UMbluvVHofhHKvhhsXG8Rc2lBziPLf
AQyp3Jd1Lo4UQtu6bmGmZam4E39TuYaWMFNUh11lShNliv+fovKOQyvOjReDaqcK8aRbOaQIv/U2
NMHsWoBMjlG8xJnfQrkXX+ihMS+FQB6t1cPzH0MZigCDTspCPVcr4wLmQ48javLcUilTXgRtJQTf
64nsSvkqaoxJcqTaNTmu/k4Z8p4DoEzfvf23lXi5k23oQOdWRlxls1sBXz9HGrNffxZPm9VViJ/s
5sdnid/LUcR83jlg+CMXV3IRoGuQuBsurXsm7ZFdRgVQk07gmcxCKuJBd8eLJiRnhuDVkJnxhWIa
Arje9cQKBYXh8xhOeS+4o4+rDaC9jz5pzxnup5UqUEO376Okfr7NSiFCMcVNFxus1d0kx3rhsghl
yi3ksij4RwkIFxi5BXaptWx4e/t+cxKOe6BYTOWnafN7QltptOhW7jQoNQOk9dWvZ1lsU9V5Osj9
2evcEKz4jZTcuoeJwqoQkxhPWrpyyWKXL2Q73XCQ7aW3WEfters1lXWba237+ZpFaxIc5G2mLsPL
j8ARQ/86V9ahioTR5BYA++nESWjKAzsqtEF475va7kV096Kj80ivd9qNyU2tinS5qufMW6VSLnr2
kx7IE3uJbCXUc+tkK9ktU2ivQpbRgkxvhze33qjCAT3z6bQ6HHjWz6Q+FeOJBMO3776Iz2BMeg78
K0xAUwrK80229zj5b+SX/wwaYFwj1x3LIUJagJruVg3vYRMtD4mh9CRTed+lDEzf5Ih0S/BuDH4u
G3B5bVUWGPiqe9mpVFWesQQzCZPLhEF1Z/+t0Q+LAao+3PLZt3F6Z9EZme4btJf8RYgjPHR6+FJZ
hZS2P7L6EfbDzwazuz/UDU9dTEuZiFPbDHIWxJG5tuH4qBRqBUeBdj0+XEVMPErvgRL6dZDvGG1Y
2g/45DZMQXaYOSxOaonle+ASOu33E11JyjEWZksDnyBpaXPxmRsWTRFh+Z8GBN4XNvqthauTdij6
6LWJ2ukhcLRsb2h2cDlpfaPTgVD+tBzeCIH4dift2Pf/XHHbmlvFOrmwiZia7jvhplOyjNwKzP4u
ADuw3YngJQuPUqH9MGFhdUSB1eEQSn2c8dVvWUzAErOiaQ7fpYPbsxDhxy7Y/LiUXzeJYUqUFmgF
VwD2t7NjWKIzPknTmrsfRp5Ru+G4311vFzjp1SyX7iYJC7uFqlFhFVW+3emgu2RAmn5K9SqrQ3sB
JLacycMoNTTbusD4g6pRbWUPaGOf3zwmOurpExV6edP2q+uVECuaHO49FCXxxwyCRwPxHYsO1awa
KD9OcW6YTdZQYC8STMTq9Vg3IM/skdzPHz2JzS8hN/udlCql5r7UVbvDvy+Z71Ch+rwawqZiotTT
K1Z5fWgxvmKm9alNXeMsw0DxXXQypqDMwKCeI1yvP3o8FPb/ZenYsGKgoYbgV5JGWngbdt5euqz5
TQXSuDJddPx429jEBONfQJoQ0yRQYgN4/hSIyetzSS36SKoW+Fw3C+78ldBz/B2ZdedkAJ9+1MRO
1cmltmcxB0mp+xpimnfSYjrkEREoCtJ9nESvSSQs+5ikJ4cLurj+vYPJmHl50FZ0/U9cIXK9vNVk
r8+kbyBJwJYVZl+wtSKvvsFckfbdXPnNPFhDMsIoB4EUJOrgXN8iV3FYdmuNeKM7GIMvc5jUvPPp
M+ZiOKquZhVHnuO5YJKfwFt2ivM53rMlldH3TUH+e1+HumERdcZ8NuwuwsU69gP2JqdFjiCFCQ+7
u6oWUH0DK/gRg+jnVbzoIYHYcNmHMplAvAaC8fgxRCuPl7Wp6N1Ww6BBfioZXNChHqHEYKmifq9f
k3WpzD2yn4keDyRyBNIyS5gFCpEZJLpPFm4kAAVc5AaE7LTN7KFHSZ8oFRI02t8FddmmUqGUSoRp
5r8mA3qIIDNPQVDFTqCgtdEX3N481+S1wzBJ4/lmtNXQRelM9V9IF6kFC/FFyFT62rmu09HPtF15
mx45SJnLcDMNOern3UZx7zTvI0JdOoy3AxDB/sIf/rIMYWsHPQ/07tLGqVNPVUmdoNyBiaxiwX/7
hMZnru2uU2kftHGMW/jDwvKEJPs7o1jVtaVmtfA0lEYTuDy2yt/MYFHxAsKFcrcs3rS57gS0DAEP
7TUJyM6d+SecXF3kwABSSceHqFx460UrTxfqiKTNMMzGHs0cVC8FNp9setD/lk/61YIpRHz9nZJB
qvr0bwG+NucrD8lGuX1v+BFhGDU0Sd5WhcOJk4RceAHleEOBMGkP36eP43FxRW9LhbnEB0ZAIKfg
HGTZx0h5wmhb42x7pwl0Tgo13kgTEvf8BMR9I5NvNW2rdCakEacBh9puYucGu65XqGpn+lCBGvgd
1oknkjk3JUKUAC6AcNVFgSc5RMY755Ut/fqG59LL8izjs3nvlP4SD1SU2moqe/23kzsKbZS9rIIc
0hy1eIkXwqc2oWPoaeAmOCsKkP6l6mtaJoJG6sbzNZzx6HQIWfdcecQSTguZjWP04/oiSpB/49xe
7Qrxz/qX61R6BJ79PmVDkEbL4nx3NdmdnVdMLcPCj9hNwyZJrHKlkrHuVMHSfYQlhkbZm/IqPFjB
IdgWLj6u1jx1HQZdl31qMB28LvCLhKTCFoF8kqP/W3ep+jJut9jXD6PAp3H/Q8igDrCaxVYs79Yf
5HE3/bjE/0nFAS+gn7zQ6zfIjurM1XaS34IcI8h5GUVdki6OdoveX91Fi1UXlZpesFlCKOavbQmH
VO9tVTJ9OOdjJZpnCZ7DZf1KsqqsdNCPePJV6QmqhnjB+6rvPNVk7wmfyHTeNHDxbDq5kywBodGg
7CT4G3h/HrSZ1nvqqeS1eU7kSOnE0n5eOFVaoP5vb49KcWFZU3DcofARTlX/msDV0pGg1HSZV6mo
+nDOiJaO3vN8YZB8QTgvBLA61oU2EW07kImpbqWnnkCi+YHczjxavTI0hrW9coSe4Is5pZyszlEU
OHxPnjTBoGwqaqtx3C8nGK5j8J2cwTMOoLuIAMaMwSk6gsUthmSNGT3o/o0Bm+VTIycXF2Ggbe7r
7NKQOGGINkKUIjgJOkDMzTl5DHG4+nnghziuC6ymvCm/mqoQgp8GnMixd+ud8DVfEo9rWwwKpcvk
1kexeHgywN4y+35syUFTXR0uFfARPZ7nq3oPQrYmtQGyXavpvQP25atKm0VJhoCG94oPJVtuLGHU
Xz941RlX/9hoJWJLwPT5oc1Xq6pJxJs0uQMW+6WXbbAQ0RTLBI2PwcHtHAqXzODYccxsLqZNLJjm
/NG35GCh/F2vXpYdDGU64fKIAHV6ep1q7XtVgoJqMxz8Q2hl9Z7kA24ffs032LY+obNvaix3++oh
WfSbm4YJFSlyDw/9+lX1toehqrWJYSWEY93YSiVcv7tIXdDg00QPMPZx4ji0V2k4cYy7Cx6sSrDg
C34/JrKPlg1lSl4scdREybOZP/9JhaEapwaeHXdpZUXXpoRm+yryrB7aCoGTW+03x61AvK+ZXHyu
8nrsjuUnlO98fbjX+ImvIi10IxCPZWI3qCg0aZF76JbbICMH/bnCw2E7NmqoFvxHFdT6YBR18lsc
QAHhlxyskRH0SUs27mBQqclkW5bCyxZrPvADAYyMc6/jjlQJP0pHF+qt+O0LIwfDt5c/CEJlGUoE
Bssd2MXZfuZiYAy/lteA8k2T4gm3e058/2AGA6DwJbDu9W2zWsLKLPPWDCP6uhAhr0j2FF+CXzKK
4/mHPmOHc9bOl+r9Vzm1KJ13tqO60AVHCZKW3B+hLChDf4NAxrjreHMiTazaN5TvE2tAyT42922P
hQBFxANAliOX9OQ8Dalx7pesmjtJNAweQmxVlouzOShw9qJBe1j+T7Gq756u9gsmrV58mbh9AFEi
JJs62Gq0kPBlErkulJq0iT5EEZOI3dHc6fnfn297OFPV/SeO2GTeO3mVT/7hlIkvwhy5aCZ1Xc0G
m/4WyG2tG/qouZf7ekrSdFLsWLlQWCzfWNlEoCf4LS9KAnFAsJErrZvFIa0NMhRgD+/KxV3tO+HQ
FHqswDF885HXR7wk8fiRZNiQCBfKXNRhi+qWHEt5wuIW2X03SCy0VLMQ5peE/cO/uLX48FLb0bI2
bEeDAv4zrtkVfYywww9RC5COPAM+nXAlJs20IVjUlnX3StRkqZJ2pMt5pS4SFU3lphDpvvU4TAdY
G60ufwogRb2Ukp2gSCywJpaQwLFAvf0SC2v7cNdnhgyH1Xsl8XmXsb3dzA70v0J4lYLVehR742l0
jYD9+diUGTpeKxlFBhT1Lb+YHH5Wj7qnaynE7rFVG6ltmRUzGFUPjspln4uM7BZEtfJIEw2ucH/W
5fr2i6CoYwI4UY4XOSogd4amPKmWCy0tvF3yo/Z1r2i4GOK+Kq6keai+WE6iN1mME1szroDjbAba
vLafYk7bZ45JTx41/Mot0h5MObDNAcdRTRsL5g41OCkaIrWtpc4rPyoyya7UfmuOMCPAJeRWw2sR
KJYqad+2NwT1pWTVxB6Cclonw8Q31pJcFmrcHW8h3rzlQkC8esIlQ2TnJW84nrh1GzOCtdz0S0dZ
2tRqDphqYnveF35fes+MUBYNsYDlnil5D6XdLCv+N4Q/U5CbgfULjWSIEjsrJJ/DrC7uOjsCcuAT
7XqEd4PniNDmo5gD5fEUkKhK4ZcvnHYcd7w3bHrJTzvHj+Akkwo/LpAyDaTafsQ+KcMrcbvzspTD
D0NdhND+tmMuq2YUnFThJYbDDuxvhOn3M0WwudDsrwcAEozmmRe8UocW9SuCvAnIsh36Trpf9AS4
6t7WchjZjPNryuFHKXKA+sfBVXinxt1dftNj7PjJzaFFh9/YUk4lPQ/JBjGdckLHHsvAXRbL7M1s
q2YPzdOa5+IEQLgbr1AfxuOzUyxJN4p09yTjkO1gmOWrBUb7gMbv5J/j77emtwxXBzEZQVnX5AaI
bJi+Ypgt4lhYvp6desbC7K7k8cS0dOSJOSd3Q2hSZifc+bLaohFEYiIFUEg0vNBTFotPvtc4u33g
yeCg/9O8Q/RL5Cr90sNmXDuyjWDDL0/R/BcVwN/OmW7rerLh+i1JV5lvkYmpRx8QZU777MHTsmwm
GfJkW6v3gVEbmW/TEpjKC7oOCPuwwH1MLIJF0ppP15c/u8UYSfeXkI3ixMwKQM3cKyBEDVoMXhBw
vQNoeVK5O6nKODSy2HWfIiIAtJQuNMjzjy1MA6yygci2JFJEIQ0vAw7y+P0NUuaiFrI5n32vRc11
Lf9/0j2v3/wAPyUyr/XTZJ0dwGdIboSTop3k1IY4Yu5bVRJEsaqq7zQ/WoXS35E2FDgGJeikZofb
adJnSSMlqSJCfxzqP3b8aA3N/kDGBx655PlJnVFg8Z3GLNPbxs2e2ncre6xxuQUhzviGddGjj94v
0cBcx0aTWEhfKs/vabal7yhumPJ7d8tuEGkBWzcP+M6QWPTgFc5hZUNYi/D8O59BZDUM/+GIjbEg
1y40+laCMf/gcnkAdlpmtDYIigyEhiCD67O/KFLSu8C6rbE7nuoXDZKc3/pjwX5/dB63H4z2zV0I
XhrTHJFFRJgRhUcBaH590NwbErSbwuBGftFAsGffwGr/anfmCLz49yUEh2TpR9FwtQtNTMjKfAgB
7KqaSBxao3yMPMccbCA7I5gUGZb553Bv51t7x9aULvqeWaDb9QW41vdGQM1uCL/whxLK8iskiGZF
UsePPIhM5Z3mgb5c8+YooZ7VnvuAPo6uklUxzRBC6Vi2V43v+EgR7oORGkTS2tA3sCRQ1BmNxx7i
O2rQBVUSvFIThLaG4I9bOFCe1bDvMRpVedx2Yk/2fLZqA5eTJ5M7pO9yFqRvODr8Gx07Sl47RDY9
r1vN31k4hA+AbtkN8ti6rZR+q++CuNPErolsnDnzRL5BxxZuxZPvsiDPRt/9ZvOz33RTYuerJpZe
ZO4zuMRDh9BaVlWNuMkHtFlG6ZHeXZ8qY3h2hSBpL8MCloYcvUnqufSJ6AC/njIbxpom5TKd5x3B
i/SoPlPrHfxIxotdbW0AFLW5H+UJLAJRUZvb7zodZbfu+iNddYI1V+Ao4TPaJF2Td2Xq0eKep2L+
EgevCs16qS7MPrgvGa+TuXcJhODOm7X/NwWUkZA0WiOkrhIawdssd4Pz2etGjrmRdzwtUx9msFGH
i23/KqbSzxSu8jnO7IJ7XPHbUsZARohZNI7WoYH/Eore8du6pPA9oKvLhoHVA16lbgQ0kfnjtQIS
74d/VpvjtobA5jZNyq5opUV3J010ptpLrqkwZwSnTd403Rt6tUuiqICoDZ16M8ifms4QvdSIuyKC
lH2reXyvMyMpH/sbQDg/oPrD//9yiZ4UchWGO1r1WGfZpj3Ya661RbyvtHb+L/PR1IGEc7rKY0Hb
YbHKs02okONiG+O9NwEv011O6ItgkqAr+lc07Ydqa2ttlNjZ3ui6eucy2i7U3VhickvbIG+QnG+R
DobZBAF6Ebe456f3yZw4xW316ppvVOs7ATb0DYu8ZWQq5GBBfC2gP5+yua0SCgmDwbntbbTDCrf7
9jBKEnMtzXp9QwGJ4opTgCMHOhl94U4zCAKSrRDMNPDJkbW8j0Fz1hJjy+y2wDVbmo5cI/9rjatg
q6sB+MBZkTdcdKrSs/BUAh0s2khb9rqX+ssv9NclrX1E0rPhXohYnUsCc8WBk4b7/SnJS+Ox3Z4A
lOKg2i2kbgV5Fg7deJZn4a6ynbhwi52ftD4ak50bQj0tdUQcBLkuuKtYiBU1pQIyCI+NT4XARRhz
ETNqqunmyc4/XJg4SXx+7c6ht209mq/uDBYpjzMxM3tpW23lr/25aICzz5/hD78f5kJfbg3j3LQ6
GsepyoH4IxrxqKTeb4DKwIt/YaeKFAkElm8Y+9dJUbR6GkyVlsyQZ/xdlfN2TwPGzDu4R52Sep7t
/8rtvBUOXzLuyTSh5Ho4GBl2cW4it4GX7HDg7uuITpDn4jKMT5tdShZ77PYAUf4fIPyNSyztci2X
jvfoJ8lPL+w69MTX/zz1Yg9/gPnDRt9AfJAoTiuTn/ltFgxh+mnANGnKDMFZaAOkoi0nQW1skvNU
40ZX6O2d2TAofLtaHd+43aa+6Q/NS0DWIxcLgBNpMcsTmR6hllKGnaJ3EP3MfxEefEwNjck2WlyL
TSJwEe4Xq+sm7Q1tHjBimzLb4xYbtM9PvJuuEfzYqWtqojg1m0bhvDu0avDWKGp3e+Pz6MS7Xg4W
j5w5YKAoU/Euo8NFBV1esecLr79Kh4rcmv0VCpQY/xk80UNlZLPa4XDKCJ/P4ZhbQxKs93MYjZzj
m3doiVNjBTzyiS+Des40kn8F3N9oVLsGfdoizAoHTFnmQ/u3Hjynh4VKTBVS6fv4QSe0F5V9IWxk
6EBGt7ZdmuUedSKgIYo810hM6/xlUUuxx44xPqDzRwq+vQ61ZAZJRPU57gknhFyRJMuUFC/QQXtO
KQed1BxKWPZRuhk7kGn5GJVKXFzRxCcTt698B+Ubztb0fEEC98TtZ4TxHcML5vQOhc0sLz2D+cGB
RLJjnGNHoj/KXMxFgydF2IE5ZeRbhfYt9G443efRNe0rhTJlXIy/Mwi8be94Mf0op3R3galnrllm
US3qMn4qxOBwiUNLbkZlLZBTajYNHkpD1ZPt3nrRkSFGikFC6fr9259dseAEjFcIC9mnjByTgvw6
hyKsm2RvCOelCt9yjfAUaXQTgOo0z8dVBgzt8fnDCrnmbDUvh8ZXFH1yfMiKBeFpV8Ul4zMNFY7E
u1nn3N5h2NaxcKgXoBoDAL+NsokH7zcI/MMkFM0KEzgfD3+lkQlLXcUFFBoF8Ysktpzv+91DV6VD
2RLuojRVwEb3RvHCWufX5ILq/SG3XNtIrmjO+UtCfXU4o/Uro+apvLbA+hMgdJy3ohAI9ZwxsZRA
0LIUlJDHg88PHrLcUjJbSVbpgvRVzOmvjLgM2xhTvZt7vSPRjrIW70p/5rvB6fl9oUgK9l/J2/gn
+Kub8Ih4CQnN6xvnLfGFdEGDssuYyLwYubv4W1VkWgwRXRLz6ElhUC+YiaiIyL3AnN+P4kmWF8LW
2dcEkMsU32hzVY29Px3oXTMVZiRJ92KceReQ26AmIGWG9GUJZRO7caVNaznJJ6AM8KNriqwPj+V9
8hbw0FUbI6eUbWeRUmOvSm9iKQPz0XOKTBePrCBmOKzNW5aCLboolBnaE8ktQn3tN2m743HmNG94
dFST4K8Xwa3HOnI8paILkniMgsmCUKbtrWu7VlvINAuQIqlmiC00/xnKx0+67P1ZwZlysEa/4D9r
1+rzIc0lpqVh/nKf0yTJ/0pgSfOkZGpmTmYyyA5JvX+6sf1oDzUJXIMPMWsfym7bV95QISyu9Olx
j7jDydgBwZ4eWWpZbIQqPOFKPtz1p5GVFj1Oxm71pJaFDTsf8z34abCuCcnBT01rvl77NmxO86UP
kFPhtDC5SDlexu3QIfQHNOrxQuAR+jYeopIyevMrbVW1aS87n/sSeHpNK3kclKz4G6RPjzHCA0pe
Tt2YDHO2Gqp2MDi4BWlobVWaJXRlikK8CnyippyH1VtJFRs9PdJ+V9ysek1pFTEkEguf2j7KIYnH
RKp/oOCv5/W7DO0QtWYWSQdyD782liLcCFYg6hS9GBY254Wl5HAEo6DzoQdR/TChrkqTvMAY2jka
WUyTyiuaN/vRZ+LwR+eTumoW8WSn3pCeboZGjDvSmpplWRmxCnsebML15xtPr4j7VY1xhqn5Wy5j
xL4ZP00OVwgtoayQkSNDUxmWD8v4OTTD3STUAwY1xH7fGUPIWqZZ7ORuK2BeixlcsOS7/sx0kbqN
OOhh/WB83hbOPKu2ZFIopDAsSqo/tgoaNEKcCv/1oKhMYdESn9i99mkjTj3IBnxkorMIvhzDBN0/
4nZCVHgLYIhgsE2zfSrfhte1Hde173hEbWtYtpOLkvyinOfquPGcupJQt7FZRgGT5gfQLL+bYhzN
z3AK5AnW1Sl7kMk7vb8QTDkUI7tViFiwSCYXQOas6F3PNx1Qk0w3lSJEShC2KAi2s4ZTBB2SGj7w
HN+lq0zFmdebySV1pJdC+mTuIG2voZqQoBLP5qrUrgo63Bp6WMkq6E/o8/K3WaLC3+MZzlzYXy0d
l2+EnstTq5wJMDTjrEXfLjtDDGh7T4VuX0dEQILek7qEjUJ/ats7+2I+Aq3Whz+q1Lgr/pq91Yz3
C+dMiBkp9dU+alrm2KryR/x7B8uGi9GnnX6iSVnOUutONtkkwUEH1TEMC0A1tb2DbKh7vRzDRcQw
KI5uHrHOFqqw1+UeLjZlYESxaLk0E9FMkvvbEfP18zK8EwGsUGDfcjOLVHvPmJcciud/pxcQtfKe
1av2u4yfMp2wriAWdjDwqXIHinSUxVtDYcKVSERyQnfvpDl8dnIxs76m7AYASf9r4AJYjHqHMiP/
j3SdTqFBTMgGwrYoOCQxXkPB9kxZO4gUC9KSowI+d1d8hBk9FnFegAkjPhouOxhLXWkbCutIadjy
q2CNx+DOUUVxmEpzF8Oi2R4aZ2PBHKq8E5rVB3Mv5nBrvgYzsum3ipbS1WQq8pPVB418fL+tjugI
+4wcNaQHt20LQO7/JHo4pDQ7zKAnbx5opMdLWCUuuvBZqP7tgMr3jcMP/Xb0alnYb8nTo7nWDprK
maU5eUuliTAsgUAqcPjW6I+lBevyaV37nds44z5zSMlCQaYusWtZtXrqS6DQi84a2xeAGkxvPYmk
pwGgY2BFwSyc7t2FnY29+9OfyhI1gHdXr1RxI427pkgDsisgLrswBQFSQioIWPN1jhuN03VWUSaw
/5HCRhatRCfhmfOW7U2OqiwFid3TJ4tJ7TVgN6xi2JpNtOWsYcUS0dY2X9gnLRHP91K8ytFgyIQV
naK/z1jK0d4a10jOre5F5bxSBIR0N2o+LvgwdU2VMbb/9ypQnGIMb2DeCvLGBE+5zWwNrj0+v8iD
W89wLjLDpEIQkQwikqnB8w/nhWCx6pSV7DCJya0cr+iD75bbozVnx6OJD00uDrOrQX6wKcPVMgym
OZKcXbzZiRjivvOQ9igrBhK6jp1ApMdj3PjPFVohGl2JKRmWtqkI1e66rB10VQTLRwU8L2pORUUo
6n9oMN4R2B5T69Ij/isoB9E+dsB3JrcCcqyIDm1+860E3eymTqCLWZqD2p4gK1p87wrOJE/ZK+E6
5NShOkfaSZcNH+gWLq6qXaIwxjBaQTOksVZ7ZZgzwCtFMXPSU/Lb1KhlE7tivij9BABh9yiF5tT6
ZlXDjfZGdL8RFWPbuis2oAU5PtYfCBJ4m+CRDkjRrFpcCuERYvjBp/ikovQa2Y+0SjJMG3TMPDPt
jskOyHkr9BbKyhJxqj9h058IweY3Izy9yy3oUI7DJD8HGkWEIwr2CsuvH0mXifZqLQmK8DVEBXEG
fG7t9PYn9XHMDUO24mCNOu1qBaTb7eQm1ZmB+yi9Ed83WqV8jxRb35X0aE2nU6TtVx9YadIjKZX8
QAFsoxFTds98IgqNyNASDC35AfYGqFBAsYLcSzvNhYwzePs2lOiD3bpVPtakk099UaOBHOM7Z3Tp
5WCzfLwZb88DiKrTq2vxlmePVmiqNEfVCfSMlS0uXwDTODbELQs4WS2I0HOcrJ8YZepNWc5XDIz8
B4f8I6RZZs7GPl1/4XR1LrDEzQp1fbE5wG3OuJ+48m8MFuK2mJaA8QmbRFZeKcODjcyWbvEGDTW2
zET6L01edZIKNImndtncco5yc5wP3F1Nw1OHwjam5EpQljnrMDUAYmTJBAT7ZeZs+ZF7F+4dk/aH
NhmZJ1bXd8XlwJ3Ghrnevp/tBxZItflpKqQZXHLBidklenPS26jclSbKWKpEHgXDWvi/ntciwh9V
xBu88YTwhaNzOh1nWBuefizW2qvIew3/90Px7OKv3eoEbzaDsv8bnLD++/Bz1gMFJQJj2k/PPQgr
Fp/SDHGxd2i/3Rxcmf0m1kenhZsEvsh0Fx65i0QHRg9GqBtkCMmXw7dPXA5SFiWAva8MZYKciccU
wGympKrWFoou9L1ThwuGYcR3987E8eLUfa7dkzISZs+daH3zLJkrNkO832vBuRMSuNmGmh69Cg1o
yNYlgwuodzsOWtx5GSwQ/JHPSlvfCUnAD/axf/ej+CVisERyr4L+AuPcjolpr1v/PlT9iaUEFWRk
J0/6z+wwUCtAoNtA9GE05OKd34Xlq2qN+OlwfwTqVYQ1nz2mtU34A0vRmnWCrE7+HNZcZAiMG853
TkzqpXHlLEgrDssX0vcWw+IYMkDGF1wkU+cA6pEFkDSQ0uakz+/26w2UpqHrzHbe3xG7+s13T5Nh
WxcXEjmlEAXV9aS74r3yK6KTEcgb/AffViIFamNvstYSGmVzvWWZZBcEPPWwKZzyLRCv244Sq39e
Zbqs8/MHXREG9dkXCzNymqbBEEWAlcSRO9K/WmjqasvxumOoXDNPc4PFHsV88E7X5rN8zpbv7X7k
QP4iLDn6nDMqvwiV2R8hTPnLend/uUyLdB8WbcQmntaSN556ig0vZ8uvjFij1aV2ovMJNoa06B/I
lEjTLP+XM/qvpaCP8O4zBNjG7b3BO96hcxnLFsF5kwvq5UPlf86CBgJUuYc08aA9Zp4VOFxgmOk2
zkSv0Hg3g4lRkw5A52gP/TQjKyTq1Qh+B1F2OVnRC9RHX45RpYV+87v74QyPnErsLBjgDUl9Tk6+
7tyPZqLRNqPb6g1gPDdoWXCmFxF4gsjJX6JTw9zTUGXQarGD2HHaYTXXxzVT85zwAmXSBAEb392P
L4QHHi8B4tvon48fwN4j1NcjSd1fqpF8YoqAkiFbTrHDy1KvPVWRRQFljx6qGa0LyNgpxokVo39d
UY00GZjcczr0/qWdKZhKLWRHU+R53XOyoXuAThK6tYvOVXfaRz8puEJNNj1wCm/hj5A0g2kyCkWX
zXBjHqiNFwRihvfSY3K3v/HdU1PxUTNa+KYgUVtY0YO5H7N8p1bNev4MGussOqvJqYIItnjWMDU8
GLYhp+lSMibVjzoNz86pYd8FqpgI1yk+i3j7pJu2xzd3ZGnH8xX+7Ef2OVBZd8zheVnnlZlttNRb
7bLLY4a3JxLsmJ98nW9EXbPPBXMdg/3+6ktGORMUF6/h6HQWdW1IIZCVycKgC9PyRDZlWly+ScuR
ZXgzIUou3F/AxEyls5FxXd7sEpXL6ty3R1SWJe/NRPK5/IFkwoW82P6Nx52r+DNyeUEt5SLrrt3q
sNHwGXmYEZSPNyIiSSAUFVN9sO3iMMpo2kdLRVmxWuFB76+mQWj0q59lO2T+msz27o7pd3/CGHAJ
XITy4nQkLqUXAjgsz7zs/5DsLKgedUt1rZMS1l+01aBf+gE/r0zKi5k2PdBPR+RiqMpeb/q2WLGG
Y+KpjIY67/ajtPSUtiVus8lQocCbrg+x6dB0SS2PJCIG8lhT3rSmer3cwjsRW53bLWKCzULoPiY9
DxoB7QvYm5+zxDtw8FW5poUte/miT3jZgfswSVcIDtL+Z183xnsMkhgkyKKhZ+ekTXinBrhgHUtN
9VxCmdiMvMlhx6up+IwjIRieqed/izECqw3ix1uP759yh4uFaKHBmk1my565/H2LtUyfZzrAbcl/
ibMElzmPQm/vc99y8l1T4F3GBqXG2Ci5vL9dp6kcMJ9t1hfkKonY+NBz7yOofEn0uwuXmkpuFGNJ
JftmKMH+OIKT8FBBTJzfukMcrZcAQx3dV1JeChgk5D47Am5OfMhdPwwTbxFPbtfQ5m2tpFUSDpMO
HBWttFNq+k4MT94OXooa2y9yAhV1PTEQRqJM8/0BmrjVb6FrUOnraeUD1s845Y+c/mX5sMVr7KbR
qdSgTaoUI2SNNJFlGNVvmvyxmUW9Z9FmqpSFq4hS69a9cQiDLGkgiS5kKqcgmqc5YRiTrsgOJI6x
WpIJ7C3Z+xyqT6d2tw6bxxaBXP8JanaTFgb1ERRrYnhh7Kgi0/FOo5Ihacitdn8qKM+1tI1KW9TK
kN1klZtHOQxT4I1SVr2IfdAMMtuO6a004aA9h3LVr9FPQ4v9LhyI7TOe5P50zByCGH1cEKwX8952
H+G55jnGLdHneyYHfqsP6rR2YxS5KZ6zG4KwT8Eo7+iFaJGH3/LcvMIFWZuSIjq6dZp6vsVazC0J
szUp27TGP5KnRSRSrj8AtMSVhRjT5CwYdepWLyqxVba4sVpqZwhWcFvcl4Qbvm/PhH+jPOstjcdR
7D8OLOdBKShO4jifg0omu8aFVkT/D+dd6o0dJyzfYWDIRLP6R6yy5f9OVnOdYSdOvMVSqUxWnCJh
Vd8KxgQ1TdErUEv+gpnhjonrQEE3yOsoUAdIEv5F0s3IaZwPykoEhxg2+QfyUS27sHiP/i534MPD
TZ01KMFtJQ5af2oqHqE4d9DCM4Cl8bRCGSex8Aj63dhcgWIac69tVBlZK5K+0pysCdNFfiCg7Sil
5X+bS0r+30iEWUirAYkp2XTo4/ZVJSn5qiOiJ+Yhi8kHcv60DJ3PRNshU7jhyAr90uJbSeSGOskT
zLbgG6WSggpWbplJhkAVTrmNpySf6sOIsQ9qVPI9lZVHmqkdA+2NNWju9Bq+1doi+TR/7zIAplLZ
cC1SuT8jjTlfkNTraHXq1lL4nkCLpmr6BtY2Xev/Vt2khCTlHt56HZEWgvcvn7ptUDiIolOOG072
ofndNHQQLBdsYce6+GTbFXVrP78umrr5x4ctGDlBuKp1tL1Dx9QSRHHWgX0WQV3YBcBbDPPgeEf3
3H+8njFlC/NuOLxOZygwNRs8jSjrQMjzq3KK3ne5niMTGkSUK0D8QQtl/iRebLNdJz4lg2NtGeIs
yU3Su2m0kxB957k39h/3eVgwLNkl8tHaRe+Kber4yXjkXRPDiPkJz9Cy75cigzi7ehXW9hKOImmd
aQusvZv0nVhwHtCIKKGyTSPzLCxmAXIloqp7VK1guL9FpDq0dAaDbVdYIOw+Qv8UgIz6H6qM/o8l
PrbpnEHpFpSpdOMUP9RGXrwsDlw8fB/rJePh2Rf7Wd6hqPw4UVB1YeQ1GbZ71xfqKAqN4/beSiqI
ZeWDKm39tnxr5g6tcbqw3H9vqveQ21NEHZKokaUkkfvbpUGS9DjIiFTPO7j+n05Sy4PHin/Vp2LC
NzV4/8iMfpMzD+Hl/4CxiRJ+7zFSMy50/eIKmKC6aMZuIXGeCjyozka+8lAEXc13+3Jy6tpceoGT
qhWBKMy9XxSoAxt/y4bFdcur9AYr/rpG6yLn+WTGANcWpdG8A7iCwHkHwnFU0Efn+PL6YrptWh3Z
1EtEbebFqQC553N9bkQGivwPRyKHje6sXQRgbnWdM31t/AYSjT+QJRVHt74ZDohpiq75k60VJjhg
CZ2DQXRZNrSHJLN6sQK9+uZg2PO4RCDPfX75E3oOtRmX2SmRoantcQeZS4SSdKM34YjHJaT0dIEC
XlEMEj3FtL0TsStz/mfpfqxeqNegXzzNixDscJ1fhitVKTHoo6aw1l2fIk2B5x3GI9B4FqDWwaoa
9INA0CNqo4j45zWGgC3EYAUS+t/t+b6TRlrBQlMdfv5QftYo5o4UqwDz5w0XxRURTKSJedwPvT4e
8jdXVWo+fFWlWvTZNyuRfFuNRj8x8e8O5gHcimyELjh7kZVVi50ZJEtGoxVBH+PguOxNsvYMi8mV
mVdQPkLoH/xOHwHqheZ0Aoxs+x/nk7h8g82YdSAh5TIGFTR/7YgpbaFHN9wO3JfBFJ7nBPLD52lO
GStD+fTagAhO7hYTZ8MMArRVDBHMZUiwmn8KP6kOYX1vUm+CWPWozUUCxl2QDEoyl4Xz+RRHihls
NxCDD/nIy5mUYDqqqXOTMPJXv0Gtlgn9J5tvEO7biGSeIEjUSYtuvHYI5tW5aVm1w12DUr0GAzBf
vK5oBYIcWLnORsFkAXLyWd7yIcHgqfwJ8EMG7RyRd2ath2Du2MGa9ypXeiIfYX/uvBJY9pbL40RY
VUyR59FJtFhfcr+mPo+quQ418ZEkxcNM1KDTF74qpXG44M6L2nFe/f23LG9yqeCBIXDUMGIcHmFA
WYVJ9Uk0rn4I3Cci43hNnqzCdom67qm1uc8qUFKHo91PUjz9hT0R1rhcmJSFa8hr3p9a6VVuVhUg
mR0/DfnQ7wB27xQlUs+rJUdQBLwwTi9L2pt6k+7UoKYk5dRbyeD+UN7F4UL7GSCTW4pCURImg08Y
ATZq4hxmwJVn2M//JDETtT5L7GXBhx8aZg5GZ031UFtSIZgk0lUoSq8Z1qarSz41T3D9XRHTVIES
MkB+Svj6hOusKaECMW3TIWnD1ES2ah1aKghu23HOPfpn4qgGnNS3TyfmV0br0CiA5YalSsz5tupu
h1xXmupVaYnPlCxsPkP3Mi0mxKeNAPsK+zbllzKDMVRxsUy6mUYqKQ3Bh3VdHX9Kg2J0G/0Zyp4I
D2KS/VidzXwKLcG3Ab7C+MoQCW2PkPlDZwuCeNWVarVQ+qIWuGrm3hlxjj8bRWnbrXpgJwcG3g7x
UvJMqEAqNQxnFyx7mGvvrmlfszyvcYKyeGfq2XnAQG2RCe3sR+4qhL2O+u2ALtgv01/AhfO0B8a1
sQzuQ60CjxXe1edR1CVtZXRieTMCBPop7uALdSETqkhAU1NXCFfG7JcxKr/HQairx/kWgElyn20v
xczTEwWeBjtQ9WKc7BdO8udHL/6J7deP+GZdoVKdy4EsFw+lF08UlkcyokXQVTGPchHbb7jkDwR/
4Q9p97/6EGzz+g+D3veTZplUgJaNtcto33gIypQh6KtYRK86eHEQNWCx8bneba5IsFImpRtFWEAq
VzPnDNF1xQFTimyNvQeiVBiR3I+Snts2rAIBk+SJEycpZlKuSh9ttqRRrlmSLrMlHQRAegkMuynK
N/kq12Ysy3WU6w/pHQY+KazMCxtlNRnOQQCnxEaFMpeCQTySXk1eD51SYNHmJdQnNlmpuZ1H7wcd
w9fMTrz9BQbuJ3C72AMhrWdgn1h7zWV7igQvv52TQCh0wWhmHnu13dZ8XigBrde/3K2W5LXzLLxs
L+hBhzsydPg4DMIXo3xFqxKvUnm6i6qQkTovX+8XMQoBwqME7gmbc7EIxXXHbuKYAk2BDYhEtqZB
hrgHYysJUHj6VNpp2LOWAeG3+rJGW/7V1eletsdYVrS37VDph/d+aiXy06ySo08jMNNAhiZBtini
vJ8VxOiJIXKroKa3F3+tlbTmBIL6Z/1rGSWDO/+I876Cinc8ed0DHhy72f8mipZE6EKe9XLBuATN
ZlsybhkoVpkR73J9xayjoklQYKYw0U/OoBlxezMMd80attFh1sO4RlMLc9bBOEupCUqrp7DHB1oo
rAFbC85yFdxTqQB/86xaYbe6Bd9C81Zmjv/sYYcvO1Q1PJUKsrI4SQFAWhPSM2V9TUn5JXMH1OLD
YpdXNnBf03Sw3zSnqWDvZmc8a816ZeLnHnaegl8ckuU6OB+bqQki3gv1ot5VvuyigtprssA4PzBz
49VvhfObzTXCCV9MRceIzpAhdvVjm9Ezb+N3z9YoVlBCL3gGES7bSTM9EficzZfaD7XL6/WZoQir
2tVqe9H9XsqlPuyFoLWRKTxmp8ZPkfzbfLZpD1RCadPj+QhQjS2bkfKkHcofpFyBqmP5zRPaPqHy
JGwvR8o2Y/1BtnZfH/WqOvq5+Lgyo9/oX0ac8I7WO46pOyp0y20d740LGPsQqrGaKnkQZzSStjLr
0F782HD0sWL+S6AziemjzTaxilIkQbp8QWgOIfdchh+2N45ADdJvvzzmpnvBWjaHNuezrWXAP7vF
VpCaKNPPy4d3Sxl6Ft4M0MLVuw53la/YoBjfGkpyQlB83GKiwxRykD9f9vfV+F0Hsla/RTY2Q6pP
p1oVd2AsnLO1O9LDd1uEyvwiaggPca/eyrTRGtyeG6dCWeiP+OstewkPmZIhb/u5c+sKQK2jvKLJ
kfUW4oRGXCLPcSeqIxfvCtkwfsa1OBy4fG54n8ZL4Mto4GyNjBys1S1awOr+LxxZcxt3S17sy0ak
zTysE2+Zf1Yv7ysEUtjDqrSJnA3cFxqz0jP2F2EXhIf/zkkFzR7L8m3RKscezsqUwfT5HAQY+87d
v3rUtyJwCPU+BVB6SY4BPuhwIzZn18/c/oyiuTOjKnJj+3+gx69lhpmip6BOUNHxlspQ7xEA9cg0
9I8Q+SsFFqm/pApR+cmOfIyKmEwK6ePfFt9q2cvvFEEOSbrJyPicWYwm4dOlAg5pVDz4wh+YH8l4
CZdRUSrN8cci8O9wtjI+iqf5RlNYMu6XZDUKWwQyfV5gP6H9LEbZnUOPJUc5GwwzyBDs8tAYRiUN
rllkF/MVfdqDplfryZ6BCKtQ1k2tDpmbP1K2/Dvyl2h6eJHPJs3xselcrACdzLpqFx5anOpUidNn
nKOH08wutR73z5towmK0ZvdjAl8ikghiD1mKZpxVGDqPQ/y5XSkeInUxOuGjs7Ix4UJT0rzOeOyY
JyrguCeez8jVRaouWXFUAwP2EMyGaZyio/tsl6jw/A+uUwjgAy6tfPwR+BaR4hZYnBZdY17qVfAE
kgiUF3tadccXTDKq3RJ6pHUvAOVT5K+sb2SUd3u8RwQ4gsr2qdcVAg1mmsTe6q0a0+ttXOOwHl77
juEyvPJegwGHkLImaDGawK36yHEq3d0XzJCzJBfaZcRm6l/niB8PKFTEsNmeG/7+Tcm1JcO8t9eO
yF+cSIwImZWrQCFY2ePKWxuJnAbCMG3A1peJJdqurWzPSrW8qQiPt6E4wNo/xy7bpegKPgTSFkiZ
LUnoUyQPwKlowMN77nfH6gSwfJCIl1+wP3ZYAUeHPgsAU/7b9ozixnblLj/VDY6izQYfb9ITAEww
N0rGdKW//gnP4aQDEBwzGNNjKOk49eoAK4pCWznhy5clPNMMiDlv6hn1xk9L8JiQ204A8oLiy1TJ
TgYRCExD0XTtz8fSbF8VFr9xiUrY9S0BJ2h0pi7i6kmXJYgsLKhKcxdPmuDpleOBKncM04Zls1Ho
G+4WuqK+B94SqaY/skXnQq/DD9isEefp4/ClYEtc8SSpI2DiZrMmOPkOrNvPaeuTFfLRIBBoTTwH
wbX7jvQDRx2O4pFTEWT1mS4rS9lwggQ25w861NP4LpMsT6GUFis1+0ZFDQ5row67cl4/5umTCcjX
GY1vHw0VWQw3636lngkqjMtawiYLw2cuh2zfzLVHEhv+2lN54zM0V+roplNiXI8rTYx9Lmx3jsyN
Vj0UlAhraLUUI6mezII3a4DgofSNRHnaqLEvEEvPBzIl3rChwFkvYvqImkPd7Fk6YyPia56Ik3xt
YopSiiinzwRu/4M9cZVXXWK4Z8yyFOg6qU6Xx79dRqdntxda2BUoZIH6EnBlX6qBwsdPWwxZMEsa
fjFStgwMYLHI52+qrcvteIJIr8JT94z2LQes302nncxi7QvQG3id8P7EmqFBPTTf0mN5GsDKHCma
+PJ4hLfdNZoaKrMYjUTjx3svNv9Fqw1N0s/foy8ElEUV+86tQKuhxAEBOcygzdXZxJGzfqs1j++Y
qyJ8NJwkhRQ0mjArG9RGIHyxlbtfb38htQ23AfVcd1Uez+91sWOO+RxNgiwZzUDmKVUwdDJdIrpY
3BjIjv0EiLxJhZ/5I6bYqs42ROmrQz/3agwpGhqJkvHwwEEoJusTcn3yEK2TUy+d/jTftssHuowk
fZ/Kk4aQxxUd8LZNp8pZSKWhY27PcQKWbyhaTIcqs6Ksza1Wf6K/sd6TrP1pRFsS9mnbKdwcgoJP
p1bvpn6G0CjWDPA/5rjY4uCm5orQcYhbTQNz9ZwtMjXvIuwTl+E8S7cImymZoTyNc1+MBYrHZuVA
AZeim0Wb+nysSUMQMWpRri6TKLQ3FENqoNk/cq3TAWWsa9fubOLejtmvfoTB6rbB+E3o9mvqC0Ak
vITmW60xz5TolQUpAzkvL7HYxov+jEb7qk6QsZms2VFUxMkoVeN45kRO8r7dgp/YCrFAoqeQOno7
jIipqPl3bP44jjB44/bB7jQ6qlvfbBFzHbp64tFlRDLn6iHHESzOWL5L/gQpvTVCPSA5ZOGC9l5z
l2Ule8yfF7iEb8NjTxJ/XUN2BvMzToKE0lfXcuBpGkkZ5NFM9FCbwT8l96qLDqvCniCQ1/SisJxX
win/UM4J5gIXfmT5AWDYpU43zKhPQfljJQnAeKwhXDhqTwUgCfldJtEGmpH5GcpteBt/tRKYThZo
GOaEtEaVEVrKTzpc9I70HPCXc6NlQ+A6avjL7L6V8l5REl8+4FDyVxjJKNVpC7A1jxnGcfiAVcTF
wg1I/751sBNvFP8kbopa9wJ74xV6DuCkyxyxhs+XD/Fm6KZoRmWM3Bswx7LptwVi0t80ZAS1I3bz
EZAJ/Idlh5ioYo2/FFZLjr/2CuxwK2iVOCbFFGNiaprEu6f4yksm1KMXEx/2vD1HNbwUxMEpSHGQ
6FKSgmF6Hf1Hr1rV3el8n/7yguNnPZ1I0vTFv1jKF0S+EziVmXtJBtbzFSUKXqUyqg10G425j9tz
/hDSmOzjsK117uMPR/F+wNXNvmF3RQmieT+P4HPbyzymW9Q9X3jEmKE5lNMS1xnP24gc11WJ36Ag
3fRMzl5mvc7xG3c3G/bYgPBdJiL/QCEipTQ4Kf4aPiR1zCdvLNQWl/dh2/mPsNZNK1JBgCYCGIh9
V6/PDVjMNJV5whM8eyxcyQ/XwGJRGtgMBekAzW/DNZ7QemE7M4GRjMjz7x8Nw5EfbiOwxIjAZNJZ
iKy2M+605TBemkaN9vcprK44IBsPu6w3flchJqWsrulmX+kTVa0s8r6/n8k86xzVW3USqwUeZ+Ta
/z/YpCoLUQSB5kCKZ7AhIe+1/HQV/piELXF1kGYXklixaZ6gaXdt2YpW5ShkcDQkNHEEcBAcDBBM
l4AfAaeB9dpNhKC8FdXqVr0SMv9mXOkI20jlUM3jemwcLozKLyt056Ml7PHcWgieBhXf+8680iO9
wz4/hz2xTReq5bblOzIiGRS9mWSgrBfwHoLZSAwatQxDzIH1b1O3LvZL4qsIvh/ObE2DzjC66nAB
Y4wuDHiLDigQcwVkueeuu7mjrCH3ljr9gqlN5noD9q5IC0MrJbu0bEx3gCNDeKVpRnIb1ZbDRWkU
nl59gCNOBI+Kui4jxNseOeNMV/ij7886/YK4EuoC2JcH6BnM4yHeWhS+kEJmi9nTyBD12aMBjdJH
yKkd5iYaKiIh7dozwBhw867yuQdtqJyhUkqwEUuBqdecy3QkFjRcgzBNMxDpD75rcwMB5AqoO9VT
uDGTv9IIPXUoRb5tLYjDcWFDfK9/KMPOIgqeqQJPEU/ieGyfOWVQqMgN9G9Ll/4j4QuAK18He9cq
DaLXsWtvi++3xSD+ZAITCx6DIyjsVJqvleryJIUuzp7C/ItHVmnWp8QAPwxl2ioJTJ4ijioS0hNE
AG4zFmc1Y4lq+uoXAhDEQCActt9+W506tqMCewXbHM3woqcb+wMKEHWqJDT1zMADoshI02pelHIB
EhsAdCv3iob2M8lTmftyGFVlN9/Hzho2W14bQ10HN5KhYtuHOiKoqQqX5YC0a+XOKtIAOPpNbmth
XakUiajDQkOU4EZARCTYjr7fjy+u43PSZXPOt8sOHuDusbcj5fPs8o8J9Nks8V1HSBuJ8JAkBQ2y
PAqNEK1nGEhsHv+kucCmU7Zj07X6adUkh34O7Gu3V1NjmE7y5Ktl/98DBAUVyh23EmddHpeCtonx
lzSpoQ5279AXeR2p0J0T/vsqNOU5GmOUUEbn7XCfGNzl4vdLMuFZWRjYdh71T914dbwIMPRlsfJ1
vU+0b3+EdvjzoCjZd4utAVKiIt+SztQttNCU6UZNcxBh2R/MRqrRVTBbtMUtmwTBp8NJ2Mliu9bt
8bO60lRwZcaDdqAqKR4cdv5KGLDeTUBtlwbMfi6LJ6I642xet3xGtTlrXcyg6jI7y5gxGhcCEf1c
PqbHCidd8WsLaw8FbwGuwIhNoZdswRikditvyFu9s15TlDjEpEWGJQC0RrA9tZ998IZAdDTdY4gv
c3gZQWksQrJNDm6CuTDKkRHNWxgPc8ucwsilx3GK+8xOGt/NWXOYI3+qNf5jmdzKgpCyNq8hofFw
N5OtphrfirYw9Z4wpUK4CeIH6V3TvpF4kmXi+EyFG2RCxh1t5oAIUSgb/KEUp73FLO4LiSLnxyIu
v32KhHyqTUjMrva0VQRYsKO+IBaQG7InuNy/VSIdidbfbFD27yFGE1qqwpMw/TRgNHobcPRojPcV
rlrH25WUaaobsE0sY1gkrKg0MlClUd8k7paVHbsrV3N4f/e0CxQ8oDcBkSh06JlzVSCJOly2Mk3l
AP5ah6Y0OGbuo6YcV3WFM1+fA5tu4gwpoZzXNk2bhI1tgk7uveJhKAubA3UJHzn4aARWwN87sJB4
/v3qcML/ckfPzX0CZ9PwCc93aPp+8B7hh3FPoTbiH7L4ofiVtZ3wd54WqDWG37DK8CW3wg2Ah9S5
OLNQofuwLbLu92FQiBqB+9nB/vesvtFL4tbwQZXI+pd+FZgtxKXQpYh8TAWgPsWLnMT9JXiCdjdE
ddok85nyU1RZG6infAvfRaMJONDnQ4b2Qjg64QseOhvL/ud1jNBubR9mwavltVHNSmF5xWdB5ep8
QRzlgjkFRxnCFUyGNOak5EUaT3M1iSCvTAXIaIMdqXYam3kA0nMt9bNSuCjlUd+cYsq2SjBecQkf
iOTa58yUfOwsNruQFiW40w7M0M4eTzWh6VejpE97voIzVF7ZcyCEXDA4k1C/wCHA72HJgo3uCH0K
X7irJJIq8WEJosyBz5WOb2ZqmmDzGc9to0DtINzWC0DaEsucKEHHi865RbyLLzh+J9VpaKdocy0l
5Vvo1W39p8n7y5UQ0QGDGLg5i4EwQJlw8+H4p2+cHT81jGojb3hnlCcT9kmiXJFHMl3jnSFv8T8F
DLgqYByv0D7nEQ2+PrJJpFvYKKeOiXMe/yqTaa2Fc6rLtuTqLagRDoVA92WT6pzzG4yZSMn/w+uf
/s8ZIIrfdLy7jMG+JmAIgjO2/l0AZT4fa88foBouWETwR0wWWZm2357Y95QbetvyGfuH9a4ilywi
oKoHGeo3H50BxHKfkqWFki4kQGRApHoaGd42c8wk5QOwv4PywsDSJGBkIRhsfwMDbiBjISDLHjri
xv+Gi9L21Q09iTILunNBwjVk1pUorO2eDO59sqMAbyejl99JJSmV+NuCelWMMJ/QBdF873b9X6+9
fFPwYSbw2/qO82mxCBqJf44LYmIPQXYT8mttWxktfD+G2rKlYPaEyhrkZ2hncHwYBMzLpDpwkCG/
U9QbHGrowmDiDZBQR5ug/04JxATryxb4Kgbg9D0W0TI/dB4ad5HZzybdKu9SEM+c6abDde/hcLG1
Zf85JAYE3cY8fHWlhQLy9Q58DS/qw8k7SE15BLxPGco5q9Vfj0Oe6/4GKMHJncZGXngZmpQucY7/
AG0Ne2WERxXadRCUIM4+b8id4Fdzkpj6kOJmhO/iyyaAg5MOApEeXx28B7tDWQ45wKgqGq4EvsS1
LrVjxoMfzFeW0AR5dqT7sK5RJjglSRMaT4fxdgOugdmJUUsWrc6cIbNC7PtnN75yFUBOkEyKtKsn
BF4FU+NglORGdW2tVYDQ0ZZqJH0UJ75UpnkmTJ2K3IKpDSeyDBNWbv8alCbSTGXcm/0pUiOwkKVh
z8cm8Ka1Gv5CcMd/kgquIvoT9S0ug2/NUN5LK/kpGmXIUEjdRj9Edmi7Ji1qblkeFwBm8Svg4J+f
8kW+7ivLR7lJLNvJYyFwLCzZz0OhJrXNUQE6kqlZJxsnWWHXm4qv5D8w8Ysl+iEPHTgHlOIG+w8j
nn3ZhiYmiM/kWTp1xSX+qxHWMRxjrtk4uagihzrX1FGMSE4GJnp3Mfr5yySAqTQwMTnCjt0p7S0e
JGEfq85XNTaUhKWhy2C4JvCr+ChYbTEYc84rmCloWxFVNDHrqOcjUcdaYwznwKO7BOaGvkxMrr7A
8Orfv0IdCoc+j83fwEAvKtD46eZjKCa3VapNcGcY09g6WvIJe5SRCqNwOE9urtyZGeyA7ytcsi6P
68Wn0C9BZSDBVEwRF9QslmKPG/iHgr8hgMVI8fscsLqBThxQBZsDoQfikKcSv+3jTThan1Xil4a6
kkcUlMtmMyS5j8Jr5yTn2jd6Lafe+AMy5c9kgzzdhg75U76SEvAZSFG1j59IR+7Hd92oBU4OEVb0
Tmar6fPhRSlEGWYXY4cakg8PEQUlOaGWlIGzVTBdinkBHNc6BKiVxijGq7N985rxDROhM71HEHTt
d9InQEi3m0QhkMQyVGptMjDJgnG+Isjj5N1fsX3FB+NtwpaRsh+IILTue/hq3et7WL0CztuoWFag
hW1PAJ/4XZR+/5M4RBp3Sl9n92TY39mZXn74Q6Q531i2L24Naao51ZicN2jNohipjTcwic2L68tf
KJMZqS2UUCZgmWHRHadrq0d63tTV7dPRkL5hxvguWxlCPaRrlY/yAZQVevA1z1HCR+S5X0bXOsvD
4CBD13cTpWFgXkU+FD/Z5OeogTzTPyqJZfF36ptMtdcp4z7MRix1Xjo9qowrLjw9tpx02anYzXCF
rGNMP0D5CiREsG6x6hgwR4PAObYmwSJ+/5Og4a1UQ69Gl/kv8Hq5/Xt2DeycmVnM2sOGGOhC0l8V
FezcFcFO7NLaGrHfVROv7FGmJnHRuex2Bp+m+KPWswxVIMfX+0MwcnXauHSyuAjZoX4n+HVBeOMv
3xRlOWQFsWVYXXqPggJ7NqbmVjy830AHEjCgfBepX6rWF+bNOpFgW4oXHNy/VQzsuuF204NhnFXW
bfjYsSpJpnYIyzFDGHNEfPjyiObYApKByT6Hl5ZIwRLG8EfrMvMWOpz4caNt9CFhfeUOAu/2Ff9X
N/uJDFWCkh/r6zlFrC7f2rrONgGmGlftUIbydc14Tu5WUkXyR1414YhKIDicElJ8hekaMpGvJhRA
ODhUnLRDnCS0E5FGrdlm7tld5+phgII341XZGQ7AdZhDWfnL0+/xSFd+MCXzT8i9oRc4dPK+eHnz
LhRuegue77wTqppJk4To8eMEcpbWn1QLe3MDIKBj8xpk9POFJgAr1Xg/lYbezhSVTwg4A9u7Xb0J
uvLw3xwHP4F20lQ3zqRcKNVzZk9ZljxoHOc4LyD779wefDXADUscVED0B3GCcNdOkvGgVchGXMvY
rJii4u+euwnZaLv62MIE8o06pHtqhTUltoa0mGncH+qBH688Y5EtkoM9j3FC5CZVCQ55rs4zWB3q
Yl2WXC7qOaOXkfot+Ju173hsvANMF2/tigENpNDzpLyeQHr1EfNb8nh28r7xeZxU9oTEdz+yan23
UYJOoit0ewggeZLGMlEX+IPfFDAj8TSXN4/e3eXZ+7Gk6NFR5nKj3I8zdLwjMv3ZvNvertxPNcnq
y95nOnKuuFnUzitdo5gTZqFTBwTKLxB3N2MAVJX0FnA2r6X7YaZg2TJTQGqcqxlAfbZ2p+A4u2bv
0wS2Mwc+I9FayZnvhbe16TRI8Lfto8bwclyydmcKhQKQGjHXFIU+ecJg0zKd97I5xacufKBb2S0b
2B3AngHAwRruCkyz1e5d1kXk6eC90WjGOB/y0+8XOMY8wxN7HF2OWAgdkF4098VtCunimJlBqLNQ
FFQmwlJRJ8anfnsaSBo14AQNj/dMW3wFugbi8Pnif4aixzsWsoQ91YQuNaqmvr6s++cJEPHteomY
Fu34WkW8qYoXoripqnrz7xSE1R0/uhS2Qi1/zGzc0CIRAkXWvfh+H/B8ATvruzYm35Pc7kAWSUOE
vQAMHrEeKNqkvle4j7aeU1mKH6N8Vu0VbMF+8vThLuTNb+OcvuzZPb1Y/oaYeZg8zcTL4FJZVYqJ
xctJvTkCmHjFb2CjW1UMgZ6MlViT8T7o1JMLdfsNCELKV9olWIVoIyXUIFvD3rwi08nvfp4w909t
bYE1EH1sfh6YREQ7m5Sz4IXaDcfqB4lMaiK8MmXE7oCRYUxXjFtihyxmMWffDEBxiRC/GB2P9ZzB
9py3vq7CA2TBBAi2ZFgfUm0dJbIyqU9GiEBNsg78m62ooFze6p35EcgjB8M1Ort9HfauJJOWX2aQ
zJ4YMcbUX53hRz1iRmwsUfiewPnM8oRqo9nZZcsbIDAk/n8zyc38jWukms/xgrWQypFUDT2YqGpa
3OnYLtTQ5aTJZLxU7PEw2ziT2LvAVuJPPfcSob9XfOT13bB5Xw72kkMfVQJkSo0e2fPK/N1XvRtU
r/dxsN5CorjoJufn2qi0savNFJDiFfr7o5/Skypuu+EyCnFUoxBUyJF/CBDsP6wyxiDqj+Fnyx4v
aL0UJHYq654HUyWc3gLUAG8x/boSg42RPmBIZYTgddCdomgRNHlTyzWsd4UM6/HPG4fvKnLHiN66
Sq+FJRKipACrsC2AVdRjVhGwO34GkRDtGmRiHu9eQhtjVDplMXSK2QmZmovQCJnoaZMR4tYlE4G1
pymaOcmrgT1l4CCws/oRThFf9r6+TdW5W9VPZDOyV8izbPPxIV8oMCM++tVwAY0doVyLQZtRMcsp
XcRkyvIcql4hDadMM95jl+ESmay25B5b26sToU5BvQrnPw1Gh/Or7DbMbpmofNadg1zgA2OWba7w
o3UxuZPXQWIydOtDdxO2klEI0OjFqcbYrJ+GGFTPJc9DpzU2kZhW9zzYGtVX5LKHtqTvJd7StIJA
aMcZ7gpoSVYy9wDbadQUglgKCcQrWrJ8Nv6YVaeIxlL39JlTB9VPE1lZzBS+uZaqqt4g1iHq9tbI
Ri8hPv8tsQ2GTqsVJJSbTd4loVjM1JfW7/nach0PJ+4eXnp3If1iAt46FHfd3Wy9fFOkBhw4cesW
VyTzcWWYl53638BmadZgF7r8LhqIRBMvnISNDGY3F2dWqgoPTx1T5FHXxS3PqLEQ3JhVUfa6CXMc
t6y0kIZKLOAcYCEYXbUtuUMMR88kdwfeg7TYsb4afayqJloRqFdgkCss3ZAZh4BKXMSAlTll4T/h
JctEeaLnLrbvRizsr6n2/X3b+ahyJNsO40QuD/pNHukMLIN90XvoxX9QFTN6wPufH3J0PgqHvXvF
eLgaGHJVmyjsVOgUU+hug23M8Gtggv8FCPgB3rJiQWbHF3C4qlOx3Hgwsual5xGj5FyI4JfmaxIX
Wax7a46Vbq6tw+QCC/lkfmDY4CZpdjlWRqxJb/1LRSs1adt3vVbpX484ITAaK78TgNWlb5LZ3S2U
Wjl/pAh9no4I7C9MP5O8M4jWMstJUrP1QpMUmsTANn/PdQIcACExe5+qTVOSbxi8+UjCOjsnlrjC
C3gArl5FIIj7ILWYviEaSetzIN3P8mdda8ZorG6SOdR4fJlPdcEQpcl57Af3D36sVBe3MFvAAVYF
0DKBnrqLjeAcswM5NpqW2UwiG8ZkCGqvZaHKcZXH2/u0oC9/XrzYRoUnhzk9Kwq/YxesLIGXF3qP
N+XL/fjU0p6QP9ikYLVq9CuW38JypwVhM/ztUy1gDKnJdHwWYIK88NL2B9qP6V7virKZA9pXp/BT
+2e/TMnDZumb8kEUfWjS8914WKlpfARq7c35htIgKyg/bFRCRAj/w1ZU6EYF7IR97EiKdJ1gVRn6
jDYaBa7VvUs7z2ovXZF754z4O2zUGTHklQuKmZ086i+8Y4JD0BaMQpP9gOhkAc9TwevD5dPegrrR
Hv33XS7IY2Hv5ykVFC2ugfiMGvtfpXPckVPi1TjYH9O6zoGo0g4EPObyPW3yP+7Ek0hIy3JJPhx5
FYyAEOwfDCO0rwPVwihCSxCxmyR3lx0347bqR8XvbXi4xTToZjRbOmdY1c/2JBG2eq3LKTxXBppS
cxcf0oIJ+VNsI+klrL14zt9yxgslRoJwI2FlJVmSXR7AKJlSe1IMIpsqF1dUva8MX/qlPCEVzQYc
AI+pc/Yi2sCkEkIttrEiqkiIPS7mHZ0osgnkDdwT2A9/zl9gAMswuxxjNHvN98ey8g1aeFgz+v/J
PTZYUKnb9XNwzqpE+rtM2IKz2ca/n5qLGq8MvR9vdNqjlpoOEWclemBovRC0TNPCInb59Im0ezNc
dV9UxeiEXMcVEfnZi7jukNtOcGgyIcvYcldxtM1Hm0EL/aPoSXp7T+esfCjWvgzJLeMzNp7BrHuz
L5b5w82KZIOQIHGQ+UzXSHNVvG/aqrbODdK0jsLkyHScfyQ7Fmpvl6fpEMrxuclJM5DNgFtah/AM
vZ+9oQ/IioIR7ejXhaAam4GvJq7qqG02GjjZL9PkEqQEilf9qbNpLazl86GCznAys0/WEgDBvJIG
BhhuI51croiZWAtmQqTM5UeoEa6Up58Q+SuJngbWaSMG8IjZfZPS9djjj4+tFhuuPVG7l2D8UPHq
5JeRz1Pqqc6kpwEZONXUpb4mTZSJxaJNXEPhxQyC7SnBse+E+gqoOxuiMscbFfFKQVR9b1kKaVQ5
wuni1FbVaec67Bg2PTgj4ku5x6tObrPgx5zNlZDeo0WwwzTibnIZ9co3mch+3zmWcyfJ5hsqgnrJ
KMYbVN7pJX5WWepIkGoBeR7fZ/WWODhHfFtcqeHr1/T71DsZcSCX8pEJpz438LZTaVzjtWnkqrYe
LlHNQfEh/5pei4JVaZ/bHgI8iV964dJuB8yGKsiwamQxejEq8NdvKey1aZnArcGeeXjSH0fVWyPp
nyhQl+UiYibo9fEQVqKKWVsnMiY6oWB1yQVzVPYiaEFrOSZs5dcDoU8YjXQX4XKtKTTHM0BPtSnL
TTAUCQ2r4C9KtyOxltcuu2seTZYG4IFnmkXJeniRbBN2Kv8SDzjXcUmNk/ENSgqBR/rBm1i7q+7l
8sFQEKj8MtEz+EorofH9PXDK0ke6ASVXSjFXhO406dyRURX7P+XpLahokdvYjQbk444PZhfs3bKd
WRyrwQFO7jNgOTpkQ+0LAtKIFxC+WGkqaF+NDood2U2tEsevYuFE5yzr1SJkG3YAMBFHH//n8rW6
bv7KYb1NZPvNaCl7p3RJ53WiR9Et823BgMvTjClaa9uT+AGhb1fubehERZSOuZMc25lQysVQVXhM
VQ3k62DVIr5xrnAzVXJemZzg1Dgv40O5hwqDEPGpxpe7pSKyHzgOij25uTvOdKuvrvALZV3UoAQF
riXYgNNVU6BV42PancuuwbM+1Ka3wKli+wBcgHZem1Lq2uv6KeeUpI3ni2HV5bdoFcADrf1RayZM
ScaGYJENlgXx+SRkY1DWv+Osld9wAHu44fcYiDihbYa1uvbXcaCCmYyGxsnFAuEfdd0Nzt1M6sLJ
cqLE4+eC+Bp8nQufyJ30u+gFWbMhRkART6QLi3xr6GSz9uycg2YxeOmakiD2cK7XGoczsUCK+6B9
/ti1mnNQ4UENEBbDa9JFKs0HTg90yJ/d36sd6e4V+2CCr/ZfF8ZlMPsHgw+4qhmdrgkJTkSOMhtA
3tYCd6JFUFYTGdbI0xsl4uzBnDCb4OzDT+ZHH+4CuLTG/oIwIw2z74vCaBd3+yHBTbgKaB7UL4av
mQFf6CtGsopGHPDSdiDcvSAnykKSEpEn8ukPjVZgkXf1jBRWGOeDs4ODbNMR9MR6Tq47H8NrDmqp
+YdFEH9O0GL5ZmcyJCwaSAWwJ/p/tV/iTKRtMuBOG8jSkgBz4Jy3ZBUdtXVdV0l1F1lJ/qhxSssr
czakhRDJutgE0KVJxfzt9jzNLneduRSTRhJyj4TFIbZRQWOlG8vW3EpjY3tkXsRLI4fBtaz4Hrlz
mlmkmqbocg8JYlNpegsm6LI3RBi3df7nq6FvSsVbt9XxOuP+1ZndygpiUa6gEPp8YqINz5JW8LgG
uWRJeCrr5RNIKwep7bPoepx0nzkImJa5rytq9V11raLTVcFzVlTEzx6kLZNevRH+kpycaPdkIaBU
zi7mxbEaZDxIEpJCTiGCR3TiLtOG2tysI0p3YGbCnCeG++IvC4rtrsWEcxtdqlh6NReW1zBOnjh7
XmObg3bT/RcOmlOkAUA68siZkHGA7x09iJebjdvE5Y03gsPX3yydAlhhetysJMHK8K27TWJBAQWV
wIBSc0OFpQpkT1g3JpJWqep2CzuYP4u795Z28Vla4UeAjBiP7nPIBhZNjLzkpgphSlV2UIYTo2/I
rv9ZWzf/dBNH+2AC+fOWtL8V6q16rIPN69VIcYXMx8PID0lIrSqdT9bFSoJGv6FABpf9Oy/DPnKN
g1u9HtFyHaI9SiTdl8aHvm7T37LC1piPN1M9mZaUgs2MXHriel7v2CXvh6og09C2gNTrldzupNOp
pPEDoVk5Pb87nZGkhbLBb9RgmaYeapwxXiCMHC9PG9AGlYd5LunYNIqEMNvBtbRwDL2JkYkh3/zp
5HtCQlLyXvzyepfSB0LRPAC1/l6vK90F3qJW1rEGwx/yqbs1IUV+uq1NCv3dTs2LJccUVslu0yht
v9z+9PcnhLtEI1WcZGtFvwf8WFU3rAp4ZPyEkFyoCJZrStqz6iZUHnhZ4ayp31qMpMNxKKgVsDOh
7/JUQNKn2fpNKZjIcQUf7E0FzQ9cWdGjQPQ/bjOVx4kprEpg11NPDdwNfkqjHqsk7uJYkB8Qb6Ll
/udOqqaMHrEAKzu2CbOJQ3VXl3dbkhFsBa5GSLV8VDSIddPFqZytYp4v3HYToMNhE2a2isE6wah4
ub4ZEd2X9g3EBNJyPgWbxeF20wjRyNaEqYZDwl51r+JTy/N5wUnnT9K98DuRAT0++APikeNVfGAu
LFn2nHRJvISPa53amOnDHeT8ULGGgvU6Nt0tBDxYIkhPO3R/kLWcM/pc+w3vzLR8k2hPTHhZ3FrU
bgYlcH3DG6ZYA/28wc+Auyl61w9yr829A69zTeSqZtGwaNKdMXxlGsihCqieED/eTrgO+GJpjdG7
V9pFZj1GXP4cW5kA0Ltc4kJ7zvq/XSa45rO0unJJRDig5uW4lkR2/E/NTIhDrn4j8XgeKegpxcCF
frxVhFbBfCWfRqixQKEnqW1o0207YiF6bh4U1Pqujy4jn3Y0bhwkscHfV2wtrSYqYO8ZyQ3lZwCy
ZNnUVbs7wDQLgPVGz1EUU+277GinBQybjm6bVqnJFs6AXvsRWYx/pbvGbNR3iBy7HNktC6hMFYU3
fuCGQlGUJIPjjuDlxUhaBT+yZjguxyt7O4kRQZ+ebnVw6hX5/glCYjJ+LFHhesX7R27+zD86shgE
Pa0aOayRR1oWVkpe1qKLxu11f4cyFYiqvsCB4M+B5uPL7gSj9kkkOFHPbpWw6/+Ez8k8T67KqviW
aCasUEpMtWZnzSdmAl0y8Z7x4lWTSKsxF+gV1bK1N0QjagASNpBJBFSYaCZvNSM07SsqM4rSqPxk
jO2qVamhs2Nkx9gaXO1QRH8S2UnRonFGuBgWaduJ7qREOG1+aE8k3ucqqlC7GHZmYg4pMCLqDRr3
vBsXP9dBd+GN+CvXmE4WWqj68bhqfFXJU/LlaHpuGyTA/csHJf06Ff7quJ/5jynHRpRh6KNfjkH4
9GPDhu6lkXrjTcAqTWSJKgrdsFX5oRYg3W4i02BwUSRS8e4exzr6oA8IdQSt++yeDy16uxRJEwSK
ZvlbZOzPb/plY6j147KsVEgox+nsp7uDB8DkfmJa9hTuOCW0fve8xETdGbbbzNVgVnQBvdkkWPwR
PDC396QI0Q/GUHebpgx8shWL2AkeZtqulOoqTc1TC+ybm6Rytyn4L6ak3RV90EGtcwzKFQeH7Hi9
Kk5kVkWijBnhM/Kq691ONz833Y2xxZWQuYnBwsOGwZA/pZl56ZasY4n7f2ofJaByxyYRQHYW8fVC
dPWUx7//+WOom3KP8igR3vePKbvv74W7Yh69XDmuXxofg4OLuTyGtxxVYprG7D6qVR9NKyX7RgqM
UImnqZf2HAnmwj2ecKTY7ysVUYc1xpvljIj+RkEwLuNvIQagtmDX5tCBb+0LUKwMs2QM7ls3XUii
Bh8Ov80UnNYyhpN88rVCu3l0AeTVpjlgIrn+XK+9Y3/76OmQeJzXCyEKKQS20UYES8+RQ/fKUmME
JcHH8LZbUHe/SPX4pmBg2qskCk327wpTR/LrQfL94ITn0zqRExGtegvHlCIYnrPLeDkK8/F+l9Aq
BPQVYIxxwpHKkaRzGOuGhtDRxSspMxjIlgAjdXBsd48zMBzloAZRQuGCzyIuLG3EWEVjny+Sk5ZJ
mXT6bVT3/IHLOzHIvkP70e3prfsvgGnjVd6khuQ0YCWQw5rYlKwX8AHy28xQUKwZE5+kxhsPOx2e
3/opc++pl8mVokAo4wzu0JVpWaQZ8IWmiZQ8Cwl54VkPRP6hdz+83wLN7Ni3XuiaFWoNS1Xm1Hpl
jAGjndS/Dk8wvmnFU5qVhxkGB+GDKcXp8GSTfLgoQmiqiKY1a5Vj/u0wfbd/YNt2SzmgU56St3MC
mBnP/oBcTAzPcUY3N/lCO0cdcpp30X9/g+MyDxIv4hNwMdhqpDydiYTKc0fa+hfRn7aCItQHRlB+
OK7b0pMd9UMUJ7AFnTVT1Ha2w5lYOAkWCvl4HcMnNB1uBahNzz2xykG3VvXWNJzhUmXfwy6zh++I
k0b7GrQMwyWPmVZoVGpGXSajyB9tXGfHyRMDigU9Sk3NQR7dgY/L8TpiD3HlTwuU8SMhfYyJ/q0+
HbjFicnFOBevIUiQIaI+Cleat2x7pMfGC7AOEbIw+XT67HECcTjXIBaTCcLe/gIJUEbNQfQOkDKP
Cjr9PdAaL2RQkICcduRDdIRExeyKhRplglvzpodgGesKmPpGepcafJpLwRcm9ENxVvv7v+jMWxNc
lQ8gRzOqB+TncLnKtort9sQeWST1qImPPYlI9YOc4BoW1Ylfr4Kljm9HmCWDYwa/KiyueVSUEqJl
9n8Ic0OK+OQ+sYYK56lVJJQL3sU2ZNqA7N9afGVS7VoCGnM+8eEVejFJD4BPkCjVvQcSXu8fEFR5
jlH7HpsOPI8gsUgCHvrdOmDThgChEKTjPu6ZZC8bo28kBlT03YLEuL51eHSaQIepQQ5huDsrFQCN
l/wyv3DbbJMTlaykcwqtXfEbRr8ZwuvI3EL4qtwZUByWdABmE+bn19g5Pr/KlhidZVxhUCAGCLZK
gFmel41eCbZyhic6yH8FFk5B3f9n9vzB1Sc4TvpEIVJz8TP6ZXDhgI/yHRUu0JUNBGZq/C9IeKpc
7ZnBnyus5MZCYToErzX/GstL8LDmU2Mqva5D3DNHS8n0koHj1tv7xERLw0V4niOmS0iIesUwlQ7M
XyxYz8XQABSVMMDOwwok4NF7BASkTrKjnUzkpvCmXsWBq8tcfGGBMXJ7RiuQGjVZA6FOuekAE8DW
Q4/RogtvPDkWa6r8KjLJn02ZsBFm7GqK+CCaHDWRSDcgMZym+DeDuMcjp9XYn9sIC+18mVxhXgOk
Pok5VS1mSAEC62hZ5l80KYZU8JCvP4+3XL8Ad5MpNscqAZfjFXx95shCsmMQyJu4Bly9io4gqE5J
O39xdGdA6u/3VxedlH2bxfQO7/Q9l/4pP0yjMcpo8pksHl3ZMStiHYFBaq39CXBW90X6i+qWj/xw
QUA4JxVoiQ50qj6jCHrD6QycskkjgFwRzc5MRwy73VWej3Ir2Mi9FXzGJ/4QLObPQzkgytrUII36
mUnw72gCK8pCPgh/N0WNxycFzQ/ceWEKXzr0JktjMCinpIrH21Fi14j8QmD5KqTCNRvtyzGCiYDF
GHbxoykU5FJsxAFuUGgOQmG3wz29rhziVSxwbqUh0cSZHZNDu4ILNFNDwWhy0TukcUzE1JNqeRD8
cgpR3zke93M+lF4oELmIpITvUOy9I0Xy0NHEy8XnYhKV7t53eeclWchCTy5pWMpRMXjSFmj+M9R5
4zE51wPlLX9A/569ynnavsV1iE2Bfg+4wnr1dQ2X5Qy61R/wdDS8/xkptfQ07kOrMCrr7ghBg6ke
bcZrc3BEf5L22Ml2Z6qdYgfpPXmWYGFPiS/3qqcig9bl+ueLiV2KYRe+EfIjhJ+/y31wR48uAJ2u
ElL42wPaGf3Sep6RvfOTxo0w+ofTvDJ+3I0oEyZLCB0cQTML3iWEyFvdRI1RfzOsfLp1EBdgn8ut
oW1cnte5HJupBlB71H6OWC5Xjl4+7sjf6f3HNXhj1rpu9uhkMvVgaxd9sqlhtwajtBohsGcybC2M
40xRX7ISS6PMMMBJSLwtBmylkHqBvLuwUA9QcBgt+nu9EaM9hwG+jJozqx8QWaNmO+K6KxUjC+++
9NCBhhsYOkMUzoSFz7SRIZoGx3VxoBIFPtETo/SWX3jea/irleuRrtF9wOLee7cTo1rtWNK501+7
hwTqsu5IOKt/ctcD/2rHRI2GyVAWR11WiRswji9pDD+O8Aq8wtZ/S3lJ7GclSgiBL+fnHkN7VlwU
4ruLDzrWDO7f5niFpaeIHYR7FgUytISZPyVNAEV9VDDkP5QuOuvRBNRPuyp6cbOWv+0Dhe0mw3eo
DQ6UcbOwt+t5pWtplKa+/YlVPJFc+1ppMgv6i/+bS3RM5Q2v+QNVE4KhI9W7kkaeEudyF+XVfyVl
I1t8GSBvUoW4mQVetDQtz5qFPmpz5QjP7NgWZnOs5klOVIiaTa2NQKxSLM7i6ps5lBZCoD4Fl7hR
K+KE8F3sYSdUt839HNwn0wnS4PIPs5qgeVxiFSW8cwJnuu1pCmIMmKrNQq7Dkj74ZaQ1r927NRtV
8mpnXDJfwFsfM4Vy0e/LF2b2FYWn3a+iLaau1w9yEAFA9MLzJ5hEaK2IJmC7lY7C8KKcp/JHVov3
6wcD82KbbzX+UQOM6OjWmPAHFzE4ncm5cdEtaspXT8uYJ6VWDSvxivDlllRZjIE4Ub2vaZNPzrvA
W4wPfP4JFWJyFloBg7sow+ASDLkquVAbJ/WHr+1JFvwlsxwledYpwMJgb9wl1GR1T42lBen01zVt
+iUtdWbMYJWjh5GNwy1HBIpFrC9PrD4eEUudMa0WcVd9Iy//jGuLgSGtF0vWq4Fbu7dmKofXrRyU
4/gQX+Re36raNPaL5qPkLGY91+uoTfM8Wz3ZQtudMrFgBaAn6Xds7f8+CV1x/Vph8XchNnbcrGf7
oQ+zsciSMXIgMSYE1fU9DukHB8Lz5eR45pK/fBcDQf9qnj/uwy2n47OpsS2iGn/xl0FWmfDKlnjX
vo1B46kIE2juFKFWmPc+DUHvEYWSzdbpu8YHbGAO8lJzTVl7PTGbsHuT9bpDTbQ30O5b6vhQWmwn
6LaWfby2AQNl6d1chdSP6oQDx540Su3m1oCUBHTBbHVrsE1xMqODElBjpTYWVfzptGSs/atigRju
DYKDVtW3kQSfqkZi1Lic4OHwDsvhhO7kGk6i3cMDYwClcGHlwanxAAxzv0KV/V3rni0IGpMYaZL8
CLHLGrZXoOmyciIyk8wTPw9BOjB3iv3G1y8WuJO/rI4Z0GljuZwJ5a2IbX5F2EhYrHrTDezp1Udg
DSkFT2hBgRMD+2+9hNd1ynyhOCnweoSeVGs6wNah7SrvEUGRW41GI7U68ba8BkYM10oQ7tdEBwrD
TrPpahKDLAiFQ2Vw8WMrT835Wq0OPsIFobSJYCp4lJnOQZKFenStnCk54XWuP17DAzX5Saj/MMJV
NF/XhluEFdUU9ecfOKRU69JBbaPGIl3QgMc/SsIj9TZ4KV//wyL8wtzSmmqydv7Xj0PcXQ/ET7hJ
z5DkL0sj5kYE0axLirDaSeASTv+qBIP1mcfQMghLQeqtqKf1WCKJ3mSmXmXEyv9Ib46EGhjejkLc
8FjJhFxyuWf8jD8NFlBhn2+ZeEid7q5p/DivXfKB5Xt1FjKCuNIsN624iJb1WwKRqevPfmE5fEg3
EiZ0LU6FyfF6/n0l+fVVBrMuy+F8jA3cxBOdw6KEsB6thdYB/Z/ImruFvWmBvxqJProQAaH4S6Y7
AshMCetzooNmk/nQNNVbKxg/0rFdwXn9anLQTgOLPgWfxu0VM6CyueE6II19s1I2EyuWlj0Q8ajR
uUQ7x9OVmGb4gEctv77/8s8tkCTfm84soZUHOUzBcf6Ejoje66xnlwOuqUdzaDkWwZfiNQ9iLEFP
mvCDPfIMhf7Bv+2MRkwZZwf/lkuAGCViEavNjJ8H3UzoNiZfky82RekpmSyvHB8PL8hXtrTZipc2
LSYYfSb7X4ZBiOtZeaIR+P+z+J7Xsx+yNS5nUYa2alrp0iC+3Qa+6aYgAWVCjKIRMQSJVdHLmZsA
GoN1wqJxNA3rertVO9gl3rv3K6VWzO2DEQtIhtwz1ZJPHQD+G4klqUgivuJKnxLAlyzlcxMAK6HY
5lDIzgelj3iDLJfrblwIWHAphCGF2khSAm2nFg3aZ9C5xJKgFtKjw+wS5OGGvyk2qQk7kIwLC8gF
oUp4eZNS6uBRsBLr85uMKlEVNXzuZiWdmV4VOlKK++DTqcf535k8i2RJM3VglIZuDhi3IAtDKeDq
4IIVf6y+9CTugDuEjiM/mJel+yvrYittWr2sG0P1NomZFEnW82OY6urZ4mE63Ce2DahBD+7M8BdA
NSyJ4OrI5QM5BtRSgNe5lf1vzBJprijUNBo+/qqHX0o5RAhvbfZLEx5kzctvHbOSw1nfGy7yDaZf
VFr1972LqB/8HsFuKhyez3GSCIpii7vttZz++meUKKFo8ZS3Xrq1iTTQDtcBt/0KHchQd5L9QHOI
AsRv4akIjCytQfvyuG6BSMtNrTRktF0NimA8qO1BKphMVtEXSCEY4l9uYRFrOSWYjekxJbgytjfe
yYMvRNiqbmnyKlB4d9CqHKph3pMzLaKgs1AIwZIzDdBGHhJq+L043arv4XLRJgqsMqg2zbkAMyKT
TSKfVYB4YxQ/wEU0w2Wt0te+ioXzHU7ofDmFINuTtmVLk7lM1dR3Jg4XpO8IJanOrv+5UwxqiTI5
ZiIEOlB3AwKtoow+1aJewbvo1RLY7zCwSe8WKOu/Yj6Z/J0pHgUu0eMOEUzi8iqc934UZ3sTjG9u
2hW3ICQOvRsxdtTaQuVfOhJNTGKvA7RgwNpIEq62COzX6LKkvlMnQQgNFs+smOhHWtNYjC+sKDFa
V8VecictSrkcabH4TQti5BZBUUMhqN7krl/TVNaED3alhHgCGiuM491sQjGjuiGKEwTysiY5VmVc
Zs1d9O9XUacRbB25FR7yRAFoIuVyS5m4QbsmFNoa3Elr3rRdW5+Arqq59Y11DvPGgF7Uls5RSHaD
IBX+t43tj0ee3KOClw+C8psTU3EJhltHnD9PkxuQqwBY2EKn4q8+eOFAyRZQqEVdsSqYrlvTaBZZ
z6TJNXf02cqye94jCMCX7sXey01RBeausnvbIyJnq+S3gRy6aSUk0EGny5sIgeismHYP5QlhgNuQ
Lcd6lGJIVvMdZMoaEhkl1rlfMGh9BNuje+CG6bZH2zpNEN7uYX34mZ4nBVHm7QvRuA/PddCzWo+P
Osl6udLwaHs9oJ6f502usFfDhua6BNA8tMJSUKtP4rAqtFFtpjgwQuZOV+VsXfA5indYdcro6eTf
+cVVrU2XqIFX3lkrncVr4/XerA7VN5ikw2k9s0Tn7uriVljeFKHIOWIul7YZ7IE5kDkjUOieA2tP
hvSBWLadcyBx5vceXiNKHWSNCU3E5sMCB1MR0vqCiWYk452gEm3jWDiLpaB/txygB7DPp1ogY+yi
No0GqLwq3dNc8T+VTsNdoZTkVubnLFdK+kbPxCtZsiGEMxmwc5Kp9LKHSrFb9uOmH+SRUeZnkB/Z
oHvBa8fGqjMH9NRLwtPj9bwMe8bORPtnTIzx2RvuPI5OwD9Omyel+nxcSxt6+plJkOHXMq5+u1wz
zYwVmduc3IE2OEf/o1dXP5eWLaNtq4PQOXIae7h+xyvqzwdMIPlnbSmTlwGUZW/+E5DiRRUFsS5s
5E+v+9lyu2vwq4dSJP5Aet+Xsz4FJ8pJkRuf/NHdLb9VoTb8UErFpYI3H02DrkIpOWefc7qs0rvK
uuoUm3aspNPNPU6hjmpr/83nK4L6bT4PMWZxELqLWgtJ0cPCoq/XtX8ZDntkDAMQ8M0vE86cWCmf
meTis0VxK+OO3DOoG3jwmyeXISCMyVKC8p+8sX9IqB9qux9mM8MomKP4vNJZ5QTCNANgWwcoFWg1
xRfjTlMqzXv5eGWu9ddK1wpjVOy6YawkGVDizeQjLCwN/TlW1jTjcNHJARzQKoGizxBVe6MrOCGZ
Tei+V5B5viF2snfAIXoHlsv64BxD5XHPoWwcIjq5BonHFa1GjaGjPuokH+Zfbb1x4S9tYWmBeaEB
mJB3rgaYX0fdbdxf0VGOfbHvwBfJuIMPN8b4dtakihFOjX4OSvVVTELLWYBRhzzwCZUTk8rK8zYg
K+dzsv8UJYltN12qaDb9IW3NMw4lOkL5w88bhSiSDfJT7MqhCJrQkGrMPbxEzHNwX1fJmWPhpWNw
9u30PvyogzAt9lMqipFgHnZkbHLVxGrGs+2+nKceQgA3GXVr9yfQLC7Ke6GTOOFFU9a8egg7CDry
e9qptZILcA9Qee909xxUkIofu70ehuTFYjl8xUmvss8ngAdVTSZkYXEEfucjJIPkYJGj1J2v8ouL
44shLhnDuYf+sf3ebY1kUrzslE47MggNsSfShIuZfP7GE7dmomigb62OVqYZCVcaC+QizAWrSMMA
YqNwAeKvRXPMFBiFmi8yl9ETLTQ0WbUf9aJBbLPlnl5CdH1I07WZETAi/li1Kqf927PlSJak0wz0
XW/aSsa2s1t3vrLuciHY1NEPTDlrik2wKoyIWbLCe9CDlRA8QKtAXs48eITZipoM0rQ7FClPTlZg
kZNgCHQzoK5BcUOe20/aEcfOC0UvAihsabD79320f0xB/EWUPfvxlJ/eCZWNMYpPUbgLqYfBsW9j
2H5GaQwnWN2JmbTDQRX5tdRVtNDyNPG4KC1HIZTuIL7yqROaPwiuhOmgXxzrVjzOeqNiYiyZgxaQ
PbnBgEw0M32vKKtHKR63KMAbV7EZRrO3iHsCoAOHXyWqWP5ZuZuIXNTB9mG3qLacBAY7WQsbYnhW
s7oPqEzAF3raXahQ68lNRxq8gueS9dOOn01dKBIjgaU5s2BI3PGfsqb/Qs/YoCfbcjoYQxOTL0kV
byw1hHprterCiv0we+xitvszSeFU7w0XxZ+0kjXeSEo6BERvt72p802d1oAmmmeyeZA7RtKjAaz5
v1FQPveL/gUlVXcB00duR4L8b5q7ZqXV/YSBy+V4gQBhd+F6RIjfqxDlnBJ3t2a6Z/xh0ZA2lBVG
M0wwtaO1ggC/FKnfirCztK7lCC8jzV5MDmSz5pKJoM9M931BxcPnZqy2tnS3sbzsVtdO2ME9FB/A
s+v0p/4Zbn30t+eekOJOH2RYevf2KtsD6c+wicBXb/ELYnd9wuwOQ0Z0uhnGnYCPjJ+9NPwJbUPP
q2Mj4HS4k9AjEbiUxbJSNqeijVVjKic6ly7LGtm4ejynoWxs2Ibh5hJPJw4MKtIP4+T9igZlQG4K
Fyt7dqZ1HGA3ALlu08AxtvCYfmehlU+UcRnkPK+jLc+eylNO4SxMUUEIgjvs213Fv6iYlb2PmhHO
INBtPjDRXeMP5MvgHp+KzzSpNKuouGoCVuSzpsNM4qqNHbW9QTX575R6rvRMyxx0vU4yEdkCfK/0
DHe0FnLtLDkgrL4GZYCAw8F0XR5OOkRpR2osez7OqrHMgsfL9Np8oWQtwO43MZRcxkLeQ9P9MSmO
+lZIzsvUuh9pBlBZwD9W50zbVEVHoxY1NihwZcvuiuFJz2Kav9IO8kK4IlsZDudlTrO9Hum0VR6p
hxOpOi6YZP6OK+wUWxWGsdilTW1oWPRIKl4jDpLnSlaTB0+2fOCFBOjK/yUBWzamZD84gzF6JFIb
LgNyZ/D5ciufTMHSicMd1xozwFJ7G/2zq1+qpr450EKA8pXfW8+wK8Lx6QJEV+Mjp2QHYrrx+vdf
jWVJNaPXNwl8UbsAJ3tUaVR3W155mbPSN8GuCe+JeH6CkBcKJoNeJxZYrLuPnWwEwTN4Vrvwsh/h
/DM+byfpkrRNwuFskccV+7Fn9pZP0W51zkYljzg2ybdyDzo9J+1d+lcxyouyRxGC9SkEZFyffBY8
gQ8dWSgC1K3ao2ji9jEExk+u5+dsAg3mhtIiaeta1rQPIq0ybAfziumIyxlmdmPNSGsDFuE3gSlb
1GVByFkxyh9hVU2LxJ6X2xcjrfYFlRT4bd8PrDAXn6LHHLSkkXeLFuwNGn3RssGQqVuPowbnY/hH
Www2xcS+okSL/tJTFN1fpH8uIAgZzsZpU5AX33VgRKr1Z1rGgJC/7Y1m+Pvi/zSVgPOnOvnC/QUV
kCaitRfbGqwNnmARBDuh4pA1p/QNqPg2hamD7GtEfXP5z4vqB+/My4QNKkKLE7MF2Mj/J0YLTGPr
EdbPbzS5iZR1kRXQFB8Po9eKK+UyuK16FvSezPA1MgTVvoshtlfdd7mqTsC3wZB2G5s2g4RN20La
X7EmD2Me8OXCWD9swx18dAUqo/A1OVZ02BwWjRlAhAfhbfb+JKHg2XN117eUozzaZvsiNtBJ6zqP
6yIRfTeChNGYPgoCiwnZm1UMI0n3rO3VsFa1IplVtZYXv5p2TIZAxqov+zFXPISDPm1NX+YEdUkb
y99bqIqpogHUCMz71AawUx/6sWkfo2TSIcLskXpeMXK/d0byFa4dOUmodESGY8gMcNuKWQqCssuR
3quGeJVt491nWrgTgLyexaqHpm9/iBvkgLKL55ogVq7RDX69mqQ5/Q6TuJ8BgwByqsakR2CrHX0F
a0YM512q6y9eY6jEQMYVisqrYWlRfszXMn/EVwTu2qyyPOjVO+Vuq4RUPgMH6CGqigOzNJF94msx
iydgtA7TPZ3mFf8XDfKHHwQ/Ac0KG68iBLF5AqWqHtYeVTV+qJhvox3Efi9zGhjsqv0xf8ujzb6A
PDwTrPtJuUoR81z9oDmWk94kbCdiolmSuNXIvNpMjyAnepeMpzyHAkMVLFufVbY6wiF3vcUIs+Oe
WFrI5GJjEq+mH71isQE15vndTZwjzyAdntbbyW0S+dDSxlkVRQWFi2hwWqJg1AZmPMOjdcgvQnYF
2DbiVDnlWs+qDW4S2XsMvJiSZXE95iFWIU2m2kUIIReh9pxumM57XfQF45ddyPRe6UvJF/7IQn43
Pr/xlFOo8fcL2Ej6MFAruY6y8/1YBlal1ZgwCmxl0KDKyMy8X5uwqF9PIKow9IbMNA2VqhpMnNND
nFY9xD+uTKdGrEKAA1VAbMMowcYQwJHXhf0Lrd+3YVMD6Sjt/v4kZeF1BUwC2Ckz4i7X42WfdB+N
dvNPI8suscGnLNuqmecAEE3vRIoX7rj7xIcUfypfMuU8UsMIKf2ilwyIC+DC7CqsZ6oHncztbA6a
cows7dDXpv0tEmmZl5vn/PVW8MbsDwexgt4dIM9v/3ydRAtVWuYNsS5fe28XL3l8JnNwjlyW1EpL
310EnTPnKIqV20LMe/ptjTTJQ8aZHUG/H5gGwcHIy0UzeuJCjhbgPwoFsaH4PvGcG1JJ7x5SxUYT
PsPvL2/hT3Z01HxbkMWFAT+ie7KpXrzb03zMH11HbtDrMeJl6B0DZ2lgk4KyeGpiGITjCITImOiE
77aWzzGTiDSjP9mGsVy5hzsG76f0er8vJgxhKLTbkx6XfeRz0dbOPiikzjL1ZKpcG5Ql5KEfYeQ7
siIsh0U+HVrwbTmkc5t/vHnnz+s0DYEsZwUGDBuzZok7fYc93FF05bgqLk8Bi6UYgQHlHftxK4w/
TZFmhSPFms3JVy5O1BJgwi+N+sfV3w2WdZinYffbb6jXfiE8fjTuiu7LpZ0WRo9TKbZXa5Z4+gnI
pTMNq3Z1cBSkUFz4rOPs6LBRj/Bc3NnqHpqghTyMLUjRSIXGWZ0TxtH9cHjaBY5OdDTrlIh4Bb27
Zrbtw6o+ZtYrizBE9hPMtIbo3+r/FR/p/nYNaTGVHbQdbLhJQliVILntBkaFGwkb0WFBkSjOZQzo
ZY7bvH0BGb1Ytv3+B+nbtCfO1/LdAsb6aOQMhGONj8QzaO7nnF7vfkIsTk/dqjPtKPCiNfV/v9E5
lSzmDcIbidJsPpRVK4nr97oYcWaSLBTVIaEh1VlMa10707TbkL0t2yBKTeaYY/pw/f1e2CthJdRn
BMomKBYGCbcECFjFeRamF9awWRl+UuGd7WRxyEy51BjdRFiQTGfUkpMH6HPCgnkqY9yasJpC7mQN
xJBvSwrPbk5whQweEFiexUW6iwiZBs2pJZXY+KbK0pwQ/OC9JGLpVhhOOpbgIKXQzsb+kWQ1P+v+
1KO/io0xUjEhkadEy/qdAk17YvgRQRmYzAD/dLBR0zOLc1NoloGUwfyy0F8khugELCJbpRNtdocu
sudgmsGtR8u0TkvatwCPOQu66/hCyh/KRgTF5rjMbRuoccRLH2e8zJjKB4LubOJQWx2hVwFqMGQR
NMWm7V8sv8G+lXxl0dsAweXaLcPR6aGO5y+vx3D3EayGL68ozU270QqUts2GXR8Lnm4CjG34VLGC
b7ieuXGNiYo7OlbGuhWzdjENHu9tQG6/uFf7+OUgN/BQ/5/246n4zYzDlbMOT9hN33bewuA2VvEs
KpJimL3J7vCUpz4CvEDa9bLoMllo38vM2yEFEZXgUUSSXAah+9wI1x3IIdMYIFUqetj4Bkgecgwi
vPXYaHVbn9ZKK/yEooSgH/Zu9z+qNPUjzbuKzccne3SxZgPuI0vxJ1Rl68d0VR7VtmNMdwi3yR+4
6sheVuSSusXl+u9Oy/9qA8HjLLzbo/Ju5FyFnStVCNU0IFgSB+rvbS8E2Rxe7e07QUhGSCzBLaPK
BeKBXry3iZYLRECpEW2nMiWAiW4HAhrXN5kbxQzrwBE2Z7GXEsU1nLFNDlyVlkNYW444l1oahit3
N6bnOv2rnSe8LitpS3Z5LkSYx0bnxR2ePyxag/gq+nncXvoqto+T8XU3920WIPzrCvWzrH3gz53e
wKCt84pMSpRQz977WDhWXlTsU58ElO88VpIFUSGtUfesVIfRd6hmXocQmB+bvcGi9UdIYpGaUL/M
IY0sAuPVzWF+SMPXWtRq2MKdqarfV6jOU2HjDfNC899Wva38nz0GQmxUjaBXGag5uRMmMeZT9/FJ
9COhvLHFlxl+RPmydep4RSqMTH7S37xdyrajnyFb4HNwjOICiAjgcvjHVocjX7BuYb4cJpPHgqVQ
jUP3Xc1GtFgkrLw6x9R6Nr2ZnGCcDRg6T6s/WuH11g8i3ZxwUvWn5Q4Y21g4VkMKsZORl/16H5yO
vouyFV5T/KLBEm//3bhaAdTWwV9rbuVWC9Iqx8WewKTk1ACADYYFo+kRaCi/9s4K+4gORh/MsfQD
hzXBWgeMOPNKvQnAcFWMLaZ6LeULO59Ugyy6dSQJh0lYgHYAf8HKwRmBdK3+PIRpfAqI2HQ4n2Qf
p6/LrY5fq5IZ1SopkfDn2X904+Y1HQbR5aYJuRXkNtkWX3wUKSr4fy8fGt/VYyXH0arQn+eXOw58
tvfdBsNa2BPfsxC0G3vNORTaNbY2NK/hS4Not4t/vLjqfJSVB7/LS8CQF90kJydSx86NKTgFgUnP
4PMwIoOkK+Ovf3ThG6w0rIeyJxvdGKXDk69DkXnWGIA6aMEzSPoEgcHhG+XGecYR+haF9a1qAA9R
Ihi87V2QrC7B8j74CWDWcpIPO0EYk+GXZ0a0W7PRs5e1s4ewjcQPOGrI5RcjDTrvsyWj7DzGPKFy
pLpBDOY/o+tKDCWCIe8Aj46U62uifRNOu/+m7JGauteyi71LlFnjnZEVvs6eGWu0dZJfY1o7OFib
kT6Iavw7/Ub3oojtFxK1/ytnHUaZ8NJZ2u2jSwCPjOZyXP6NpRVkG8pqfNzkKlSTf/+cSmoUq4JQ
+DZ4cK2J8cZpHZQrirVFG2UOaUfGaQ7fpIiHPuRACkvlAZ6U3qRWjNckIVuGBdLkhcKX6QDFKm1p
h153cIyx2pQcAGnv5beVQ8UWL4dqkYWwTaVg6KKyWvYWN2emIEEQ0SdZizodt6tNg7AtiZNtF+C+
TfZWPA8nGNWh1EJMA+p3ljODmGWoZwtfFp2BiseceKN8KEIX8KsQUHOp5N3QH1v7YQjgqGlOUZKu
aCFUlJT/4knPJxRFesKlDRghNrKj0Us7L0N3xKC7+MNgwZCNoMm788YRW0cZY8+i4MmFyLr90egJ
9/gxJRqn11m8gXJcd7mm2sLbHTFhhM3SgfatLRPYe4tFOjuECaiAHBlBM9lhmY2B5qVoml0pqT87
qrmhYON5wGeRGPjdEPzhxpaB3bOeuyt/ur3g+Kj/HJhuNOynB7aGQIDFRtBBUWlq2+pRyrc8EvuQ
Z4qet2LCry2hQA6e7S8TJFiEnDh7y5qG01P6XEPWWirTYsogvlkC2CyKcQE7U9RFSSXXDK3mvJOs
Pgq+l1R9kUb9ZFBmQe30J9sfHjGdPoCy88CxmeR3QUr+ziOgcNnCcXlIfqUp7rNFaLonFqqwDhuI
P5NU6qkHh+UyErosglgPunERhYf9GnsFJt0HKLEraEMyGXAub5JBsGHMKBVZuzjV/2EKso3gFapT
mMXCl9zAVhOlUj73SW0LSafQ1smZBM+bp3XZ9n0oDkM7P4aCfkXZtqaFCUqPIykGDpKLYfxWtC1o
9+4IrSZxW3N5QGIjvJoIdtdurEhw78WES2pAOdfgfoz9na5PFMHrivwcCIBT5sZnmocFuQ3ImRmX
hwZ6SjKXo163py7TEBomFQlT2Kb9IIIb1IogcISwrM78uSCPXzosYwSL8e81F7RXvAsqC8ur7wUf
n7/bfvxIZOTgrj0PgTGq1NyDBhmXFyi59Ob7x4oaVWuITtmtr3tL7KxmnotoCpYNubAy9WNWJQLu
Zst4U58psFNFtYDNhraKGZJmHP6Twzdlel1BZBFVxB8qC6ikZT0LRD6ZVOpCfdFvp1O6oaz+vB23
98HdnE5R7JvN0gZC/PZv9wYPPK5tYTPYUBZdWjFqas1RHQIpnEceweMzujX/Tfw75zHNh+dwm6YA
xiovGrNDBKu/2oi54jyRm7MgOgpA6F9BT50GBD6WGgo++BSV36EjcAniDLoY+44JEseO74BrFKeI
TftBb5R20eT/Ux+sq5rZc1RV1X0y+DmZuWZgpB856goseTIOqnRv+TcE3n+RLZH1EEIwkZt6C3s+
5oRudc0VEUeCe32yu4QM0a/8+gQUVcN2rn8KpfkEaCM/swyNAH7Bf52cf+mm+54m5w7wUVbfx3s8
ZbXZeu3Lili82NQotGDprgiHWvKtIQXEsiZuMcHZfZ+9Rbr6zhFEzHImWxqihrJyOu70pjSqGsSk
OC3VxAUVbqBp+ZhxNgUAxtwcouMsx/uJseL3UaoR+DL2cey+/OW7fsktrOqIPAwd8tdRGNtADky4
sd56Kv2zUSLzH8YQRarL+oeGVW/gLkDMXUvqFH4oBj6YbQWq7him3Z1cNRYnzSbPtZElLcRdd+BX
BJbWL5rsWydG9/vxNQUErr/pqpevPVzyJ+RmjGzqZkYKuPiCrTe1j2NKaolsMBUnfGf52SbHoU6D
FlWjQJ7xgcVeKw9gEzEnvDpF8e6XiUT8ybhR3aokD2joOaY3WRwA5AhxmZIDhd8eMBWVub/z8F6b
/WlLaIpAGH6htVLhNlz1SgAZm8SG3gnyGt6bWxFUDHv4mWps5l+WfOvsJUNGk692VZtWolywaaCl
HW4SAAeLpk93setyFUtIk6FtfUrt26auiFazMGlhtieoPnqdEeZg4czET0rGtUms8bO6OYYL88gw
biiUdG7LBmTTGPlyem2IcgA9Puc0BEDZGe2t9TyHwN85tQV1otSRZbxyhuECi3ZByM/in/qzg4yJ
wAPIRHN5Ue2NtgSfkFUeqHPkRIC1hFWDHgXIz2EoY8quW++t1T/9pr8+VkWic07+qLCPMxGAzxe+
iD4UnE2GRcdAXPiPru/zN3LkeEFIVKpJfV045mhluykHvaV6YI25udeetQQnK4KQcQjAMhzOU40B
u8Hgp++l3guC6uApL1PgSJhZe3clBYu85VF75NLvSwonySLLm/hh03Ka+kQLN+40OB+dH3xsPLso
vYsVdLpbd2UgZGbfr9g62PC0M4bk3PwL6qLJj9HiRJ/S+++c8X+76WpNWjCHG/uioIdvxvjGemrC
C7smv+Q5GXdi6We+y+OTZ49mUTK4y2YUeJvVjDr1vOBlUUehVRA+dxCe+UJTIzXdg1RW9ekUf/33
2kjsDimuBRfSswywtFCiT3BvtqnkX8CgdNPpSLyTN5FBP97Y8ptkUmmmpc4RdHJggv6O7xgFjYby
PlGAn0y51NsjWW2UmmeeAU9V9KBdVXVtmrEM5+0G5NnYoKHAFU5M1dqmwIAiJB965ecKEpBB7zJ8
XAYNm1JSdNR8KA1YoabZENzutMWq25GEXHDlzoo17y4URdiewMKYt9FczU8F2IrXoVsmllKtSNNL
eTCxzh1wrm0CFAkfjF5TZYMyMfP+bFQRLzdyuno7Yvfkoga87xK3rpxgzsV04tWpNBBMPm1ZnK8z
NI8wxvEj31sCf0KRgIU7AEY14UuuOOe6u2EA8Wbis+C+BV+lM7b5sMsWRqRfC4DoQDFaygcrePk/
GyVrE2V1Ysay5AZqlBdMzqyYGLNqwhtLjFT+OBnovaRlLWn5B8oQ8ojYFauf9RCieuobn2fch8Z4
lKXgZqkMjkEHgfSLq+044Gz2jXDYFjdK0qnR5/4nbvjugooYTcnqCjV63/vAoT1LtUsO2KToD8CY
ONNewWg9dtGg8If0Ui+3hQXMRLSl9jXTC6/vno62gK2LYku+z2jFjwEYqZcWR8E4q+C2ucaAAEMl
eiCN/GDCZvKROVXKzudKsxn+f1E5d2HrGLS2IIh/tuz/GRLi53boyivD8Kq9n1a8wRaHElr5DGCg
Nz9GYH2ckYGIjDUHkIbXwa/Sw87YhGKaxKv80AUCi0U3hNQoGTrcTCLJF1Iy4EtjAl+z24kN9KS4
nEPbgUCNGoQUlKteoz8frKSeIzheeOKe2xVA5rfj9sT3PKf7X76rlkF1xxdlUFP1a3Yy+jjg2RmI
pl2RdDq/HXK79GRr0PdzGAXAqKqCX/GPbtvieWxz8BdrlU6MD+z8VkpklYd8oCJTM/tPKgwPyH2L
OYK0dwpF9owRaF9DD2o5lUVkDv5bm95drbQkML6irq3qzA4VypHaaeXg2+DBJoB7i2POEAJpN1ED
3MjMKag2Oryn2atwFQIqWvwHlkStTn6zYn72EqDfi9IPcw0q/nf1xwm1shbvV7vhZ69XEfMZVEkW
pHAwkIGBVTUNa7xXNnSHzuGuzu9IZSb0iU8qMujCfgqtOqWybSwFGyng8OkcDKvDA0qT4bPoqUUi
Goygghr9dsKuuTVl+z57pstfTsEeA1zWtFZWlYC4MUstRJypxRfPq/qdPgmvda0DwO3vg9QJfGRA
QD5/El1alvdHpmDtQZZtJfIZJYmvHAk3ZNgaqE/uSp5OPnqC3vCMjcjz1KVk3Df6d86JAXyYJUfX
yBeCb4mjX9Tftnvx1+mvemBCM1iRYpI7tNUrch0fHy2HjOWMgw8LyIunigNd9PaBGQTqMmrZ17RY
Lf62EDvgBCFPPlRM1IfZEHO9IBXhaMbRcSO5XFgjr5R4yORWIcou8jM2SWcibs/HY14oFEQq1veR
Ya0d4AmrSgURTWOYzDyITB9jWzTZLXY5eonX9f4FewSklfc9q6rT6jygiOVWfNZcXqmWsm48DApW
EvqdNXqdUKxWsKP3cryBhX7/wMT3SOaK2JhP6O67LCr3fskAQ79b6kUEbklSmciyBHCF8FdYxuzF
w3bYYLe+hopOYw6gUOWS95MWrGbX3s7OtHqe+WyfLfEudEbH0sJu7KXjvLl5kmKLv746BY+KhkGE
GuNZ6eAUL6B6l4j0kNVy+pMz54E41fFSK2TAuBEr1URPeMc/6A1AtweSgTIR8Ttw8aeKHWA+kusg
LEg+UJWoEk6GqCF2YfGtAhL9OaO1oy0Lnmmjnc0UFZgANb/BfiZIB3SaJ2PwGqSYBvuPtvtuZqt4
RznUcwej2zt94NDprEMRx0u+w+9tVvoVZ76wbk33ASA0NxP+qOQP07gmu53ckmAp8Oj09Hl83dTY
3VKamSVCBKkwQxGdpuqXgRpm8c+Qq+5Q7cemD25aWsTcmasuI8+BZN2jtbwmwBKiZ6MB8N30GEkJ
dAHG+ptSJAAv+cU/3F0dSeIcgUkbq+9kyhTtwDDsOJeTY0+If/+CAZlmiqt+rONcjOyhZF4bHOE4
TqqKcAdrlDGYmyyV1rvGKsN+/4qds7+JbSenFb2ziRrBJZuDk6q+DCddR0cgybU9WfN/pO93LuAA
96p6wD3FcvGeRHYOrFcaG3UFsKl+Y1GIackcwhDr9UDJ0vSlHchRDKYAq0WtsvPInypHkcVEHSNS
b+ABlx+tWwaQMXH08wp80Zn+rcfpgjxldqXzYNBzCVMAc9GSbxWFXEh7LfuJauuUQeJ4DrgxEvU2
MErsYADQ1t3tzoTf1azRjddHms4HQ470ByUBs5xwUyJ8f/9Qw0+UTlmBt6CCtyktMW88JjK6wi2i
vAObVlwPX474h1ctTPvZib/Z8cLvg2ECrINSBvs3IYCqwc+4sJjNzfvv4l20H6zPO+uirPUoog+a
L7RJAHXsgikvp0wd5Knr5M5xgUYhf6kX3Q9UHnfrGglJIKWpUtRu3JYockAklRtXx0KTSgjcvb0n
NYZg1vU8nRKO/eUtt6XIp3l6SQ9OScnr7lk1bJoGBwxj8ZAToUh1o+cIkwxKPSipzNc4fLke5Qru
m/mPjkvbnyRDDN/uSeJsavtdpznJHr1hqJCYrR6f95cTKAbuvsNN5HgJi1Vpw9Z+W5ekm3dIsf8j
XNC2+KeZ+NlOa0FQbBU7+JjgA9x94oXN1U1lSlN+aohCs3IsLP2Y24QF4IydPT992nK7EoDxyMDq
+P9MnYyckbP7nSdcYtnkO/Z8wy3nMbCoS9hcBFVyhK9OWRN4BIeAgSazt4EB9883JDsbGThngxme
wbvn2Gxe3psRNER2QDDD0LF+Yz/QfS2EtpKEsQ7sYmi5QOHwGETxJKCbWWbWAH8Ha9e82h+VoX1l
FeKlcTe5haaNYGfwogPL9OnjVO4bisdA/heL4OalSdIKLWlBCy12RECVNcjuIu+9KQ+QX55HVPrN
7z3PvNIcrFfOfhKyRmSTi46tIZ5uQMxDQulgGc2lT7NxnGQRnw0KzjD+09peauDPAWZKI8qllbIb
JWLJ4mVw1anfO4Khi4iAfBWjMJMQUfgQXeAj+54ncPZOSD1oIJmS+15ZhYd2xV+OS4cLbp0xNWXp
l7aFgNSu1myaBTr/9ohm/COty/RSF1c37iM5LEZmommxz1kCNV/vPNQhHf+pFJhjaOSsXoJRTGPM
7g199oA1YWKQyBD2K2huWqrcV/eZLmjg6KFi2xq4a5dAluqFB8O2bHCCZ0uHmF4V57wFE29BF5xX
sPU5Ucd8Mz8bsZz+iWK366LzqXqhq1r3SAHs63kLWne6PFiwzmOFi/Cw05pAUSH3tDHlifu+i4ko
SzQNAY6NeUuf1MnGursIdmIPWtoeEGakLB5tEfN7dA7FD1wJd93eVFwREDW0ZqHqcYD4DOEL+KLl
XJZnzKI5JChZwUYGsfByjKkTxzU2M9I4dPhQLvgEviw4zts1KayCX2C6rdxJB7Jp+3Cs4hImwgH+
VnpU25JnxUpEGPZFdPuEcFZI0YM5p1VYM1Br/zH2Qt//ThXBP5eBlFrBkAZ2wanPsahjGcwzgSTK
h8eo+W4AC3TBtTWDeaZnXhYk15jbCzMLjOEQSMe2InOgEsBxJBhTQaYvJbHtz/5naQ2AAJjkBPr4
ktiOuET9ZM9QYIDHoXwMtRzPQT06khqkW9GNU4nYFvQtbzjcI4aVWapoe3hZrJpCJAUQUmc/UuVQ
ONod6k/kjRzWpcaUU1lKJ3VBvi2Glu6d9v7FpccIhahd/B7Ld5QwlLXo1DwC4t6zpbTHP16toS5n
xGim2FBoSWl3FRfgRYZfkbHwOJlxZBPHHSEBpHV216DpBfACMuHup3HoumsdI0mm4NvupwFiGvDG
1hjEbXQbJfmBQSPm+Poyaizk1NryajhjWcRI++XHSHVuRnAJ/zxhGmvjxJEscbc7GKeRjdeoD2hc
hHCScLwoBnqIcygN2zT4LXvz93lEwfEN1Odnv8hXZwh5+MJlMfS2qES9MwFPuHj5XrFNNLgBPFlv
BCLTIc+7nLyJFBhWiB3lkpPcC4NJyEr9r81l4htG1oYWb1k6dgwGK8iSi6CUys/dlud3hzJbsRJP
yYaGvtavgrsXiizU4dtKJSBGg9cObiuZrCbPxYhnmRQeo8h2W0BHD4XFnNPg4q729ZyVuxdxyv7e
jIDv1PoIuQnYqec9IcIQUpmJ9itqQu7gPNbOTefcNvU0zlgnGZCBZ/ICSkJ/cc0IiumD46LHWavP
9IfhF5PuKKie/qWuyoWfn2C33VvcQWfUddskIcjvu04dENRZw+mdpj1jAyGAaMPhJlWLe9q1nPV5
7JCWvkD144VKsKiPv+QGwe/jQezo3vE26rCffuYGSpPBEJP4DmszMNoo1wWV5U0Blh9YlQrC6o9a
GHA7saaU+miQWcu535FOLQpvzM71MV2QBifdTC4pELlyaRFZG/09rheN1HS1KTVPOuSfrQWt+lZc
850RPxqdmxm4Cd3JS4eQMs+o3EUTkl3jMKokI4pLpXnZ2qtJ2IPV068iHYMPLspktjQfMIsm6Kz4
BMUq4nLjrk6vxns2hERUMP3V8N9/Hsj6Hf0bOkk+lqO7/UP/EOiytO1jlIk4fBEUXJIPBu1EnunA
zTiM1dgf1WbktoxfF4ALpwRhmiv+8ISOrIwLPg6WUKrLxq7Rzn341DBrppE3ZO2M8pU1lbx3bsdu
OHiAq8gy5ZpUY6gzV2mTQwhSrCTwAZdg+iqV7ph8jOqbL298gS8n43jdfTxR9eVtiuZ9mc2X0PuK
b3sTElcINlkOcC2xu9kBexzC4aphNLevtVlXtJpIluJEbBNfNRgDqZbmIIai/h/+JIdwXr1fU3jJ
zQ4Kn5BNGPlx8hPmweSEuPuNvYhlBuTr8oT0He4+VC/bnx3LQfCs49fF6AbV6s3dhtUFhiElqtr2
8VuEXm2HVdU8mdRdDrmQvNgqTdc8pAyIRQV6f8DSlnt3uAXFrtcADZUjROlN+BGmvE+qWWszOiA3
72ouWjkQyb9c/2xrh/GrSUWtFaFKz2dUwqk+LlOjuMOoxoh0diMKzfjJVbSpGBTYqr1UviN3Ero/
7rJRgriMi+q76C74Dern+lH9lYEVvATORb/KoMs/5QdJf7EDFY/JwDn3A7D87cAViYGVijEXfNQE
4NYfTIQYXceITft0WCultqExr1TN2u/o2P775tOVFVnc7c8TarNfMYQTlG36OJX/UP2X7NURGKor
+R5omtFhsN5C+/JLL5GMuTk34eOTwlytZNsoZn19xrEbMNg7AJFhDiql5hr29VshQQUzyK7rBU7C
RzHs73AmlCOzHwQd+L9IBhNudNSFtrt6UXp5eGkWVbex/7WBrqEaoTKD3tBJgL9tP2cXAtiPUWbQ
RJce14YOPtC5a4v9e12SdkuiBbpyS6SXFzcEcyZ++h0CNQ/JrRGWn6BGRMq1MDo3CS4OL5tamLue
DkysPlhZZX8bz1XmMJwFLMYGjQXj6mTPU37PIKK0mGCz2jw3X7bi6zLZraRtYuBo44WCHlesWz7J
34acmPs1IpmjF0Z5sMnv5KIdMiMR+orHsB+KexkvxTiV2giGwScBlYmUWGtcs2lnpvKykfIqpazF
ddyukVFqSv9OHv79nDxMpNFQE3m3JgMJFOtz9+mI3IXYcjtSznHoeBLwNRDtIN/YsOqx/pGdxO5n
V2qmiPwz3Sk6BoLPUk1bc8RuDP1txNo17GOJmPZQeUKFGsWerhzYrivAXdCjSq066VqVgPUpxYjH
CSPA+WrrpZFjsdPznE1VijftKS+yfGV81slYjPmJZ6I0dLDurujnPJV7gmMX++wLLnM6hpVBuSxY
Zhkwer+i+v3HlI1GgLMG1rfeq2q3x6meLb0PI1Z2A9jacX8S6EooVMHm3oDCH3ICiClinqKI3UVl
NmY0twOd3szYXfMeg8Xv9bfWwCkI5JxsNgAVTULPQ1NcZbyeGfwm8ZKSp2BvpET+KV3irYFbyPYJ
GsGcvqwCFtzf9cCXAJ7pUEHsVFO01Ze5Ty+ZiZCuDR+/2clKtsA/z6pJAYD59Afd0QHwkW+Hl+RL
g32CiUjFoxExX0cG7ytiwYmJemI68YPBq2sWNwMo8IZJ6Hli2sLf4rXLkxAtEAJprr1xp0KMFIvA
u33zBV0Y2LPj+JMor8HghHooMCEqBZ3BQtwhSxZJUhN5qBGe0RvCefU+ulfB7tLnQC1Yu8ky/MND
8jjae/e3AaPiqhD/V6oz7qyBbiUFsAEi901Bdn3P8baUQps3HC2tl4PM9ck4g8XBRYIg4Cd2/6gi
KJ++TwPWH65pRSCPGuv925giGCY0hHE7joTtn7FDUfG0SRsrYzWKy4LGtVoBwAYlJYScFXEtPCvZ
+56GAhOc+Ov7tWDmW7cKNMxHav3Vl+KKbinTMMBekeEXZI6WmkiTVqT5EUxGFOqbXLD8HwK/GaWw
UZTB+Qa4GYjKdpAhX/2/mYtXIXiT4lAGuLThUVDl7x/HdWJR+OAo6RLWxrHkuwcFhCo518XkqNXu
1zuwqFyhIxtdQThZ/FejjYMTA71sEVKLvsKNiJejS8DDNspGqZ4r1ugU6IXNbpcjVJA/IuCDw5wG
adRANIvVqkfcvLqC8MOvUdPNbTUQQIKY2J9+jYqcXrIY2JhaRU3BhAwk3Xm9aVIVLxXqjVOsoeyz
qwAUF4cEW8iG34SwZ6I5GoKTe5qoRWbcgWqsTRPvxTJ+yslCbfo3pn0YRzxJ8TqhX3L33DIQCSr6
NXNRmuQmzM0jyoBdTU6u77lASA1RfNFeICB+UyrgRwS4gZzSG+AzbXwpH0RwmHcptVyIdFvq4iMI
dg0YEP/N2hZk4ruEBHimu8A4xMcT9XVjRUkFRvlesrKVLayyNu/UCHvWHLVIzmxRzmEsuvYOfxc+
heUe8vcDnL7QU+G13WRcPDw6ljBoyGWZX9TiEipYKUDQ70I91ISnFzGN9d7J0Yo5c9COK3ErmWk/
oIrw/HfBqVbOdDBBmjGA1BBuinM36GKX2XEX+dQakqMeSPLM3q5W2R5KQK1nSHbHCHfgbi6t5hT5
y5Gr4w8XEqTLJLlKWnGiXmLQcwYv2NCgEeSSam252yw5pzuU9J2+9pyMEKnI9BS5bKEBGpQUaWjo
mtql08TkMiObJDB411ICZTScs7kg2Iecm+oyIoUMFMlEyblrUKlFz8c/2Qld9djo8rrYPEhSRGFf
jaYT9AvLXyBvQh7xH8p/5Kos/PIUexhfwV9Dk4iRGlX1vT6OMDAgqssKkw/ikUE87m8BUEmpKMs0
oZ5vXk01GGv2NfmryqT604kJu0DlDSC4DVS4IViNjhzKMkQ0QPvmX33Y6sky1fJ66W0CcNd53Smo
1LZOE1itA6U8QZyJdn72NAMBiSuQTS0bqXOYKoRal7m00DtlD/fhyxIEhe6uYZaM3WrgEV2+yAJ0
ec0LnWGLL9/9gBrbPTgWm7G5H9yPTiryObbmy6RfW6UNLKlh8WhK+hcF42Bw7Ek0OR1ayhnvuJnB
6f0vtC1unR3r0bJGAYYYueThbqrRI6euDeo+U0ti1lyuAk8yhfW5mhTQKTPLVfhy+/LBYZfXj2W6
VW4rIm2vfSXfK0V9vcJZsRhzXOQ/yOjSFE92lNBLhNzLKbQHb3YIQIcgxpACKFlSeMoIPa9qqcQF
rDhamJkrvsaifqAEwlu+Q2EbBvc+JYzyLwoR51/1GAZikezmggPwHLqnQAjStYxrwXFIU5qOCIk5
OKLHECcIz4/9bqBD5ZqqdRYN06l9tSSzzx1IAH25gKH1ulG5IlPX6NCtCjvFzoswLekj/EJsMFYy
AGmHwFR3Dw7lENGGW0qBMbw1bbWDJD/yAwArUEsbdS/09/PSa75fLmX2cgbzZ/07ehuD9Ztzwpe6
yygV2WgUt+47j/O96rw7hBzV0QRrQFAAIT6TZfkoG/htQD76u/TUZwPqNGsz+ZhHo3eRhfFnnEm5
N1NGF48+1sUjfDQlFfi2iwSA8m9tQ8CbL0V8uvPo4OhB7NaNdDiZCnWeZHtrdnHz/w2htzTNy56w
zzihr2EpGYciDb7oGg153z0rWIX68WFrTQLzT/J9iQzI/AmuoI1v7jrw5H1AUkBEiQlpuGXF0oDr
t6PpwV5jJgKzHSP9J/s/61lkqinnWXMCYXISfHt5sWBlTX+5BE8aA2AfChz9zUO33x4HKh16GL9e
39BNrrnFdQ4ZevKL3A+4xxzRSm6WO5CnebdjVq5JK2hus97o08wuk4cYkxKrdlh0DBmwXyQICJht
iC5ph7wNBe+UkkxTC2heWkj44cOdK8Zvb0u9y7Cs8yRQ9aNmZ+tF9BXhqeFpVpKY+egcTT3YeuVB
z8wiXmX0+dvlep9LDn5H+utzM7Wk78xes+WHiEQmlHmB9rEKFEtIxmMkY8VOyt/f+Xjq2B0w0Xl9
2rsKvfC9LOUebI16wwf0TmBydkGLSzuHJUxCS9alh4A+I8hmCceZW4sW6DIr3d0o4qqweTmqLy4j
abrISmjh7Xdj+tK9w4YoyZRvJ6RvTJXO4VICcoLX5uEiZVh/oHB0peFY7fb3YnOalzi0dRGjCrQp
XOC2FDFvOMNqNrlp7WWu7TrUOYndLjJh3t/MgwhcSOJwAkwYQ9sYon/uiUHZF8DKJE6GiZw93ci9
J+RXjtTWyBrwp5S9sm5Z80IPRrNguKbjkrWcdTOHIsJmO/3UmZ95+9Mr/7kAa0usvZgNlp8+GAFB
5OJk8VVIryHQx0AVzkS3Igjrfi/mOmangkcHU5S9sIyHDfhg1Qtruw2OtsQkCVwUq+V5x9XBNN+/
LZzBxdIpnlG7n8DVCfSH/p2OHQEEZoQBSdf+hJfywEIMIo35ZCD95SG27cMOl/g8ovJUqzK779qQ
DWXXq+4A8PNE5qzIVb+zZrWW4whNnAbgcmCk+9/5mT4KsabEJy5zBg8GNHEmJccB+P9sh5JCkLGH
MtN7NhhtcLsAYEsAIQ+Whomw5mXEEat9UjPvwi8+uqhP9Pi2yJCI0+Q7icqQircXKfE2A5Gmvhvf
XcfEAmgHmk23ZHsPaxhZ+Y/EHiMW4bPTHjheunl+eM03wYCP2vznKeBGizDHHolUqChC0jG1yBhN
bilO+TPa19MbMOAD/iyuPi3X8scXZXp96DX8Ek0ZvKfCOpx4WFhSl5jSX1+zixvtKNn8Y3EfMgy7
ndQe4n7KSxP8p2zZqNiGLpRgCOWqRZAJSWcgRpeOSo3ckZp6lpd8tljqVXQMRSxHwu7lFnxojM+0
gJLzGa8OYs+CKFUV3ZayDya4IrvLIRgn/tKCkUSsD/PrQKVZunK6AMcj/aETJkiqluGA3GUQiR4u
aqp29SCHtX09Yu4OAFF5BWQNi09wxzMPjRruGSaRqfnv3ORl4h3OEYDtCmLB1lJq1l738++Jn0xE
RZ84UzT4oJvTEhrqC1rn7SNjx+4evFELoh34FC7D6D44Tr2lsNz0wiKsGRvUylS8qM1Bf/DQ5Npl
jvQs2okrU+tsL6InbaOCZlc9hGl0VcCrHxsqknO1r8xiMu27Ow75z9tcAnN+ESMSKrYvg5KIUo0Q
13eGMmMHiOclS7Ajbvcc+QXL99CIBKQ8ykkCkw1R+i6xajk8+uv6lxWoPssLbw/0lROWr/BnVtyO
8bvk/4/iVE2ABJIotZkgYNQqE+WovC9ccc43XQbz69l6Ihn84YVsrbYIkKlc63gkmTnef0hx/CeX
gXxXlYPueUM/o1Cz+xH1zJUqrXz7n0GRyJBr6UBp/+4Kts8BLquwUZcn4vckcdasOfQ5YnRmH8tU
Z7AqoL9D67aAPHnaZRYy4eZ0V6mnYNH/b+15pgzZ5COqn5S2ql1Gp8Oc3ONKv9UHiNaO6+YHAr88
bVq0jfH5ah6vYjstrVDXX2LfMaKWlGDbSJ0naPm3hp52YJM9hx9X59d4tAFLS/oZ1jcDj5n7ijbm
RNUlCEBoAKEpcnxOMIj6O5rF4dNavV7svJepiKdRO7sBkaHLsuRs5JcCQrc3WrTK1t+qQJJiRK1M
IUBcRXOdSw7n3bX9QMpbQ6Vo6Q7iWiMavYZs5z9mkeqqe4amJI8yPjdCh0MHDrhDBUpi6pgciAjG
uALrtlM42g6bT0ICYdAzmWi20FhemTaJHgE7SkkKnGtBNXit1Mb6tl+F/wQ+Uthdu8ymCmbR/7te
eapkDLwD1Y296vtLj40jZqcmqprnEvy5vkhx83hv0EofrumhPMGOdoo/1UqLqTbyEaWgivtCGdMi
YaFetl5rLt2ebAA+qx9CiIbMkWXt+1d5l3P+xAqeBm9xsViM+Xjar4VGbxzE7sRo1m66p+rWu7WX
SQZgxIcMdG/qUiwDPnc196/Dm517kKlZclZzb1sP2ODuO/DqchNsNI85ehGk3vErxI7icXAwxrI7
odhrxBl0gMVxlsMah7JRr3sXCywcGKDK0+J8KqYBpanRW+p2osA6t8WjJ3RwtWLXV+hzIO49O13t
5E1g31JeBMqWbKUKabkQTbu+I3fk8u5Dc+2WKOOicOHmaVDFf4HOeZaTROGLN4AuJt7nvabk4XVm
yZhrlDd6wnUeHKCGprzJWm+E9EeQd36NEY5VbURPS27dDu0ZmMZQ9btihrbRF01/HDankLUqqnda
egm24RJhOdQHjnmYs74YotRuIDAA9RTIsycAY8RE6y7PC2Abyx12Bpl+h+HiSB9SKmLqgIx88qLi
mUAAyCZ0HAd8SqdZytXPaCPYV8rLO0ydljMDzn7ZVs7pqbKwijWTQnUjbseqQmmgoO5kURWKtjUw
4D05yiw25gqgS1BT76ctY7mKZXUPuVKMKZNvK3XQ3VKfDn4PNpq7dnvZbmXyLR0xo0GJlgl1uovn
X7MeLLmI7389+UDJA4gcYdi0G97I9T9TWI7OHAzZfDKI7vv9pMWvg8KkVUjDmfhDteGJ7Jfkoht9
hvb/1z775dOUz92sjN8MNNYNmkcFkAXmrSRNCH6bpOpvE6iGJYV3EKAbBAO43KpsD0uGi7b+bE80
2js7zekYeIqI52BZfsKLbs7sMrxbBuD0XvGnrD7SNv3s8uf6dMYYjtz4kw0iFgc6AwmFl1hakz/i
xgDl4h4jBVAFa5F432eqV/d3MjEdW0c9ZgbjV56nHOXYvQx2oFw4Vuz1jRcJRSQtrv7tWYBkv0Yv
L03H8Bp51vuVrkn9jPHrQy9sTdwI1kA+p0WZAX1u0B06z3zMRBWIaxOZ/F96cwYsWkLT5K5rx6A+
/GNWIgIs+VwvZROYl3oKweSpXdAi+pgWeDc/0G/rNkBptKBebj1D5evy2uxqZoPk8TjQybx+03Wj
rzsGkQqfkJKHdUYi7foxOXqrkUGofsAev4P8RjhXnpwmJ+Rn9h/50Uvaim5hKoGRxtznN0Z4AIdI
owhnyqpN6P21EP9viJ0N8DKg4nB6S8xy16v8RYTPe9m3xK5S8AvtNWtV82LmleIgY7v3hbIn5oQr
K7v2WSaStx5/a/+B1fc6iven238zBsUyHoCik7f91ajGGyuyMRnUjIK+ujt3CeVLPa1lw0a/u5v+
nDhM1wwDVfCtlE2tbzbF1a4wVZYoggwzSWgkQqWkzgfLioBr/whE8RNKCBOlpC36YKUfQtzQpcdE
LzzKXkwK8XfXWx4Aup3RFkLYNf9EvNvMGdpWBdBqJ2Z6wxLedJBT87BXrBsXxqtnb0y+VOWASJfa
iTLxrqz1XTfbn83PKGeVfEnEAKOiXLQjwXV6AKHzyK8R/YYNBpmYz5c1mnmWw5CraUqwgLEoBF5x
WwArcqE6KwwfctphHE4nO2K4yVGMjSB7HqbKcmiQlf1x7Ukk3H2ttGKaE7iqalhDT9Srq9VbhMaw
EJBpaVJa6wvdEhj2ERFMXzOtEbrIeJDRakkthtab1N8lq+Z2Zm/gxD9UmzUIhTmpgSc7CMgRh73d
F2Ja2QSIgvFeWZC5AxsPxcLpWTS7Tttua7JJ2y0E65gdSf+DpVNDbHSJatHw6fshu7A1sItP+P4a
H/LrjDEpQ9FFPvL9e8gWfmF6TYN3ap6gp8YJLj4qUB6QPBdpNyDDDUOLNHZNemajMhXFHt7v+8yf
KQkeTVKYE8F8MhAZqyGluL4nckCaRuqVTLw2NBrlCBmSW1p/B7lLGh7zVqFoipsPoGXpyN9U8A3O
PzMHTa3WOpolDud7UCt5GRj+wd8yuaAD3+dW7RIfye5OEedcwLoSK+ZbunN4RMsucO/HrILkiqTU
wIPQgqCEl4EhyAVx+QG/c2pzFqtmgB0G2d/4ruEbjuOJjjb8Z7T0Kp/3MFI+0nX17SNVkhFsyREx
djwuJIFvbHCFizlAzJddvMWC4UYWh2q4BiXi25h1AAI8EUP12guJk0jKHbXKgt8//lzJf2xtA6YL
eJ0BGUiSMU9/7s7354rhU/yhxbb6QZz9E+0WbeLssfB8wEIZiT/aL92S5mSDKaQ02wDS3l9qT83a
Y9V9+a85FaCZRiSEHEP3gkfRsBrlleU18Axjti3JACxiXQSiJjNL69W9/pSOZJEYGR9tt/Oq0HnD
LOVV0pLBB7+tSm4/3VNgxiVvAez6XDbEWr0TNavwrL9mJzPP+4q6eamHh9w+Z95+A1VJ3mR2p5YU
LsqcU5IhDnY9K93YEkHgu4AnDLoRFr4Oda5A3Dbx6pVQzksap+X3eg5vpcdxXclsqhCI1lzO7st3
eId8gamAyAfm9yjS2x6bClZplN4bA0DEf3udKPnx1TWnuP/X5lGl6+lB4920Y7NsnRcHJQEjb339
yKXOVrBiQ+r/PsTJ0nOyBn+OqDBrKd/8q5rH2ydU71nhdacRIONaLsGCpEf+slN4sMmVh1PReqQW
PXPOT2jhWDQSkplTjjXMh9ay2cRpPwc2kSkD7/d8gwBVhR+Cz7JP+I5n7FOtrilVtKc/TF6GD8PI
FR1GOPUoH3yrQplBbvmPpVUXG/bsz3/V2k7Utn8y6wGeVY4qEUfQhvLNpFgBkYavKJvIujk8QRKq
ElPQzgRl69nM70CQ2kIetKW2gonEJ6zMPjXz7Tkib0NsQCmo++oVAHAcfZV/MxnmPB0PrxK7IJc1
lK4XnOhM+V+zdzfaSkTxa3BHWhffcMSF83RrKZWLvanAgwD3+BbnPR9dSsqHZMRsxlgD2nZzgQiH
C42ixKQ56OgZJvWE8Pm++MEB+5Tat6s8UAwfF6J5cbRv0DXm6/Nwy8gnkpdk0IS1WyrE519feIPF
4tV4+KcKgx12FmS7UhONwzGFwYzWY8peB/RUdTRIV9PqYQ5Wa8KENofM+rJfHZRXJkJIVepqGmOz
+nuI8GwiOkBI+dfK/tHC8UCFdUd4TCRdF6fd/5Nj4ulKVtJgPmkcn8e6YLt3qpWINuSNSuM141Y7
khelC0cdTXw8w+N3P4eoabOdRDAmCS5a1IVOOZUYZjT5x+Nsx29ynH3U7ov9c9RUU5y6Fu3LRefX
y143VgNpgtFA44RvwdrUgf7UNWvKC35Nk4oMU3BcP6z6I/+sA/7drV3OSYtrcOhUWhKdrwrfN9dN
pdPqA72JcXQf02YsMxcPJO2NhX0AIgXdsSQEvfqFpbAE2EoqaIGWarIO2WR/bHqOQJjpxYkysmsp
rlhf5fNFb3RpA5LfD49LMa4rk9kOEio/j/T+BZAZ5iL+2aDHCf8vmjQgpjPytbB61+V0I/pzbjKN
SsbHLpUV65kYDBq23hijbkagqTcTuANgZZdKvhrr76sveF/mbWAYgUxs13HjE8fq/CwU0PHKzw4Z
DO+scpoQqJuvqK2m8LGXarL54pDv0Uqn5ZhZZEbqQn9LzHo0DV5VWuQjJXO/SmktvWKIjtAKc1hH
ok9D91tGCz2oXjeyR3iW0gLh9Cq9DVcpszitWTrDZ+97ya+rIS2ebOi8Z+FQtv1AdyOSz4lUE43o
gUjdEwSBMYypGA82uTDfMMnF3XnQE4u6YHdRoFkzlYKLD4q06LAhV1jft+eeG++Hz4s6SFoOr+/u
m0pO+JshZug3kaKQks7rHotLFM0SbWmZ2YDUkDM4oyIJcyIY4Bn6VSrhk0R+4e9QPx7WeYMcj9H0
/57XgdnPPLK8Va/Nbi6ETmjzKa5ewLNkJXgoJH8eBVWq38AxHBeQHNsE0YGORbvSQCAFyjMitIkz
mLME1CaHUjVLwAdW43WsZsdvfBcDNt3JMZER8/irOuugpRm7USTwBa2Y8Fm4CTJkoEJ91/ftghiI
wJ7kGm1666cU5SHjPgqzu8H5BJDRR4idvvGmVT4eZror261BRkRCGeL27Yujre/lbs7ZrJ/KzTns
9nJ54yeYY6LuwyJpUYfplsmF2GXE7xwQ4yw0NxkeDFFGoFmOu02DKACPHbxBwMPwk9vKH1oUIJ1u
LUoLuOFZnB7rsBtPM/0NsKT1G4JPW6xadW2pWfwDDQWosA0EFuUYW1POlnUJu6Y7Ot5mVoWawYrB
GQjyirko9gids0scvp/C6vXdKDE3NYud/IePiWqXpMkRuqM9HSvlrKSqUsL+ihupOogMOlRf8qD9
lBoZKdlUNBm7qQxroXKxVOLWKvki2mxsJ5s9LQIlrMZGSblbDHI6yn27l39PKgG3XDss8nwT+j9J
3qBpMcmxDbxHbrjX15XONghMqP/P7E12bAADcHIJuNhghT/YoQOA+9DSuqaIkXfb+FUdqmceBjHS
aT60ije5Zs8SwVbQvVndh88DIseftPK7yzU4mg3pnF1cpj4A4MmQi8sMBgfucfRO0FCxScgctKer
ks7vto/B1al8NEb3zjWhhULu3/hMXJSFLLmQ4x3IDu1FWgghARVbdOd8mElv+2GFvKnTckDIzvtj
C6ZexNdXg/qYGRwo66GP2EvpZeOPbTaOe/jMLbMQ5nA7mj9tUHYvr8bSvTnjYESGRC/kKmT5HaT5
ARY+Rxd0YnjdLnFDUdXmN7w+o6ID6jErg1p6uTfONTPsEM4VY+fZWgGZNyNaPoIqUO1DB02dmnq1
U52hsDKB3lLWg0DVJSGrf1hKYqRnWZ48RBqCLMz6aQZKvSuaztoc/XMWEqXnSx84NprM7/6ckjam
XP8usxciKEuGa3nLCpNRyqIYS7yZw0VSHNjAp0K9iIsqgoyAz21Vuvy9B+RfPsvQa0SF1NSlHWMB
ZWINYB78G93qQIGypY+mezRx+OxE7GeBauF7BD9eju2iqMhaRulpQK0QyUdv/+omrjhqu6XhCKeG
gngg8w7nJaHdbYPxFmUeL9HNl4w5VibB0GeHSOkMfBIan+8lVQGm3MoVMomiX/gS8ZqZbsSLPPBE
4VrVButgt/Cmp1AW1Vto1uhGBE4ivmYzJbYq8tbaK2kSjA75Icwd584dvy7hXPQ05mfwfaarlpWE
S1NNVwUNrGNMAzMYsyTfy/9fIoz0qEKv8p7X+/DeaDtZrzNRhPIYc2INcXvhboPRxe3zBtLyPNNX
tscurjbVZihvMljy4laDybvfbmDo0bZTHn9+3KhQjGK2Nflj8QYNm99m4BsjbHp4Y2Ri8b6OjrQV
lNbSRDI6rkKGZiU0n79rMmH6VH/EfaiiiDKTtbtUEelxi4C/3K2kDV2wnp0d43wL40aZhJIcpCuN
3KU9CzFrf2Rs0nqdqVE+yiijXCzSht31CzyRPB7+QQ1ANGwUhvF5NymCUHrzIk7Y/Y43vTVdehZH
39bIOBzE1zyKqruIduS5OQb0pmzP7ynNpEOMjwX5sgKSxwO+qRqMYjaLrNGldMFbMvcxzR5b9lwN
58jzDHqcik01VNkoiwaGdpFqqyak62ix7T9zNjdfAgOkOSUwIafQFtFf8coUo49SPiFGZW5PfRY+
UwuWMnBKS19mjkjilsVIBtKrS3M3VrzwN1dq0fVPjDDGtQyaa+H42b/isOd71uDNYHXptYb2cVv5
YvT9Ex1d6d/UIVELnTsDSXoXDJ1tJ9tnd3d8BeUVpQaBUZNbY8b605lr1hPjHHUkp4pr9QkeDA2V
esbyP08O+NJj6qQNH2x1KOH0L0H6O8EgZEwr/hV0QdJOMp3KNXNBt+h6i75bVuFUR30iZG2mBK34
6Qn+ph9S0Hz09qLp5AEOkym9qn2hJ+jNTLj7rIeNDTh1QYAVzYotX0wf/uytSW1D6Yv9lGu0eCQ5
JpmuOdr1p87cw8n/4+rccIINgm0mJ154ZllH5YBTOlSNsVySDGVIa6OEtGdS6Pikn+9jCqjgoUIr
bc55Q8GK8EbPLVxTP3d+ikbKInPwpEL8hUBT4Ogd+ovQ4+gvoTCdA05u4bZhrnphcf8zi8Yyghtx
Zh/371OFJVaBhRReqtLYO1uHDHKsakNQXgXX2gPcr2fE8yf6CQGKbOXiedhFjFSGNaiFnnzrlHmb
noLiFIZPHYdsGZR067JqcvZjLgPQrGQfCmaulhH1X3qJFeu5RYsXTo1Z74jDn1CcCpBFr41Ixy0v
5jx483T8W2B8L6nkfsV02JUBA8p48AhoMtb7iBMVKFKoeLjaX+oq/GpD3FvJFMnq5/Ni6HCCtVn5
512iHBIrnW+1/po2Q/rlzVsJf5I8ONIT26vmE5mhSfikOa/upQQcL6j2orTjPeVv2kmZmuw/IxVC
4ttd0BBrgXTz4HPlG686DLWdwM1VCHwaUEB0k/uRxPVpEFNTisvAqXTz0zpjV8n/E0Jn/HlZQUtt
mmL1fNNlZ1L6q389DcNbYrxYa3jVMsBzDPOZgJ5J8EVQKGWQGCUgjN8X+h5sq1SHtLBad6cSyB/V
rrje0VTl1MvNAnzQd4+5TZj2KdJ6ZQ6A+S5o4pecrk/zVzbPf1hkAzFX5rqT5oIvdtKWciBhQhzy
aiutQlyX8+JhreLN23dw1xX5/u+Djrsu6HtKfRkLZW0D2HN5gJumoVSTyedTBNPiCCeegz9vtJhq
JxkxGxi4PoD39k3sLjcFnHsIqp/03hVtEGiV6CPyzU2qZTfbzTGLkJmol5Z4nj+56BBrXgJuTM70
zlWHM1fMuOytODoUHp3kNorXEi8pyAq/Os7kiXJRo8JhP7YsSeVsXo9RKhbhIROnK9Z68ErCXu+4
k+BDpBF4gwdDRJF7Enfda2qqtf9eSDaYtpijdgPmlWPesuCV8flKp2/DGuUj2ljm3USunkTKVhwj
9rHVAS69xMjbyRTC67siusrdX7nE5+tqn1+6TUxE1dv8WR1CUiTMz+iQgKkRJXtoJh+5bzU6FhWA
awNBzwtCjYQBT236+ST0bxBrB5+mGq0tJPDxm9tUfKoTgv49NgLMg1o9ssNPqQwy48l9PjCWbr+H
rmLRTy+gp+7DdBsxgsVG1Cs8hWi6gnKx2bsYkFOlzyUjqk6GurEOcSMpJuM/kkhPkcq+XQDhAqkr
IGbkX/GaSEInFhnGYPzwSzHxP41MLc7NXOa2RZHIZxpwEaDKQHr633ZGBT2I+6PuZ75PhcfkhYSJ
LS2pSkMmiS3CiM6jcx+L2W9bAEfttqqP3uaX/lhfrXPO0I4IMul2IFkLoJ678uNztWyKpgIktylI
FPS4vC60WMyDVc1jQlQDEWl846Mh45ok/lk+A4LW71HXONX2C9JlJtyxc8umWDU5GkRW/mcfYpHb
NauAu6x7ahvqqbnOlMYzdai+mlb4Q0sbuNnvJtf1kwp9Rvps4piv4vJVVaMT4pl0GeZ0mYDFchb+
343thxKyI8PYLYLtgkUyWa9yJNt1+e508CwHMIJ+AA4/La4v5MJLHwj/o8Uc2LuiLPBw+/MdhM1+
QN0iNoDb5sd+7bmoBn+kPHc91rVExcViSuY4/WPkyUMyvrC/V6WULhjb8w985MSTR8gnS6iL3kKG
Ii94Y349Cm3PI2bxyAk4pBYqRFEe9rQkjMzHd2MVU3EXPVRTMvcNK6kVo98l9wMOUpd1t6sO5wW+
g8ElX/v3ChyniqYlFNaflAtkZh2Gwz4GtjUhG4N016Ugu7TXDOi34EfsrCtz1Ky8UUfmfOASwbrF
584nSQonzkasxTe1lKdW0atZkmFoR5nDEPZZKH92KoSdLFSLds8U1SQJ+b6owiluZQYxxpM6NHM6
C9GKTi8LXnbEIq97GVM5NpxaZBjbIud0EOLpD4/x+98Zzy0KOw8RV2U+HrtquFdP/vgxCQKBb1tw
GvzaKq8Pb40fnQRWvvsrSUyIdWH3gHc/ieJa8A42HI2UYvoeXM2mU9DDjOSQ0LYh616NMmrCi6Ka
z8z7OMFFEbEouFhZ2BVZp76WG8271OzHHdKZnJn4U7Fg2+bEN+6CqvrLH+sng43KUZ7bIvAeDdp5
3koiPPgs8oPWpe7HBn35YjDfPhB9nIEhtZtwftPWvzkaH+0qohA9atKRxZrXavufeVVBQBnUyBNJ
e9ev6S06jbigxivikDsDmyIJc7cVR7yK8efzIPCBZxmUleXeTYPA2HVKAlNLb/CPsT+Dqg51UbzM
+k7KSuFnnJgWgKZdr61dj+o6al1TS2E2m/jWmlpSD2zLNJY/dmWFdr24OsWlWislEKUA/iWYhPTG
28+HAiv0MHY832xvJt/3U7/cQDZfBsbmpWJzALWntYttAWPOXSMJTqTRXU3bEr3tfo8bnSzrCOSd
3jaP2lPvJjqy7kD5s97VO3shJKgS4c1Fflcl/qDb5tTNPcDlbKGsCuJRglnPB2kwYWl/PDVe0V/w
hVmZv0LCvUQMmo9WNHM7m3glVO4gTT72euRMNuInWQjK5bqMe4ZV96up6btNjhCo6vdin/MeW7R5
Cy2Edb4ez6J6AL+Zn0KSfVFp02QFA2EM8nQMyt/I0WAdi1z8OXn9Loeev3Q8r0ZcYSyo1RYnf2HK
5h+nz3Rp15LAEsSW+LF6i4VYTbBfjQqmobay3iszPaenwWIRgkfLeH5g5v6yA1e/n2CfoGZySyBj
VsdsCGvb4MEtVAe5+fLVqh1wo+prxgbE6Gg84SHScaN3oBmdfy9HEkOhaSA/1AOTWU9wHlJof5FJ
jrwI++syIWY2q3piH53ctoNf/RqCDkNMKg/42B6o3+/02eFc9wAcoHBpkR/iaxPNkRSCn4AX92Uq
1o+6VAOBqeEeVlWmFzM1RdlA69VcfoudSgpd0udiyBN1tEMOpME7HKd96nFtLYjLowMa9TxjQuge
VH5m0SfDHvZ7IRBlKpyX+0Y6uBssTwXdRR76ek2sFS5c2+t0WhIzfJTISqjc30Ka3nXSz37ZPj7R
x8YwKjMnZ8P8dYD369ErOrUzFT/JVOVDBzVfh4td2kLaxu15hBK8hrIgjPrRUu3o8k2LsieXrFYe
kEBNxJxZnvwLauvkPNiZCTuMrwPXlgunPlnXprz7GIdYJdY8BdZQS4sOmvzbfPmHiOavhKUF6Qds
SIxuXwh3Mlkl8Z3X52URdVZSQkH98/Q7GV+dLKN7ikcgqHWBtX91zDVMAO2c8qArpSmEqXwhOs3T
n80NYbArfgHtlApBdD1ZHqeNYRcGGXLet43+NEpajg9FHlciFXMlisCt/6ktFYnA0K0LQSwiCUmh
pFInHsYHi059bIojqvF6K9eyV42O0shgc9FfWk1juHrNPGZVozJCklodduGpdhC8uCzSGXTK7OQD
UtdBQXY3UQjL9W1xD3TLFssn95T5aV2J82Nwy51bX1DIRNsyDtwW1Yx2cXuZ2D1vLuKifyOeNYLg
wa1fDEfOpDgPPosOlbv+Ldf1WwgDFog4VHbjyLOPoRKO7exvV4xlovNIPac/EiyZ6S4uyTlY2Aaw
ulOoLv//EXcNtidK+FgWopulhgoklsklGYzOyO/b6dDZ4qsalAmH3OJqbiM7eOs47KnktNRglA5a
j6HaDTrhsYXKglyRhJ5KgKjT8POvlgG8oyu3YVhS719wI/RxemXQSg2O7AlT37TToNXwMc4AfiQl
SWFLicgham0JhBVovoOUVstC7ZUFV1srlDK9oyaD95pjPOdppzXYeGokGX+IIN6+chgluivLZulr
7cFAW+l76HF1Gcj55QLEAHCap1Ir9VyyROwXQzSt5UT+SuU+M8WQLVnAZV1/ndQ97iYXZEKKujb6
cxeBopicxAr9M/U8432NALesAU4yuOp1wi4KuKcewXRrO/arfLVtr4JQKhnFncZFVR6lgBBYGy6d
sfTSAik9Cqw9h1544P9kn+kogjsr/mUgfRiuXBYHD8AZW2aczxsT6Gc150pvbFoLIKyIPzUoNRGc
IkO2LsxN6UyhN0emHSzilmwEULg+eiKWXm7/VnVPDURQRUwmJ6GPgh/y95KRSbFzAJfOmvsdYbPZ
+xo5noUpKXZjvXEJdVMkqSW92BOw2F1TDIKUc3H1r391x6ylEZeb3Ym68UqGeJds8Ic3TudtG0U6
jcdRtcNuhWduNw7UmKo888wmYQkJ3gHyEcPlcNCSQhH+6dyqwN8rGbkxy4A1QDvTnl64XL7r1vTb
Opmn0hCFYpAVXA1aG4F4FkuQh9HGbyDxod3m2ETSm/LYMZouRkusW/qFf+yn2AoiILjwO0sl9jy/
d5Ojs+KWvT2V2jB+6x2+7K+c21vlR7HX3WERNXnHXyvQ5gN4FHGzeivypLcaCP4tVS8OMm8ymq63
h0GBO72EBOlMSYBZ5Uw8qIMLuOP49xwsMqgLMYmmZ3BVgrAM3NzvZDyUaySMENZg18fCOJnOeFFQ
51yiCXTjopTSfmVdw1nhVQ4+WV0bbgraStl6Lnazyfcy/pr8eUlZzx8CMh5ybGUz0fwTw6/pV1oW
aZUa12hbMVkK1ahiFqbI6j6halm4pRIjFUhPNtBHiPwND67JEApgIdki6ZyfawlSf9KXlAvU3vyG
sDTZR/Mq20iOf3e22oAv2sw/qLo8KwLv660S2MP0JhsXtzUHoktUR01xCHpS5vgCAPmHQiVlDTj9
qkKMO/GznQGl8Phx9eGjVp+vLlGz+h60lyyqxWAmd/beWpBCFq8kfvzIWB2AWaZi0VMno1kxC9pJ
Fakrf6CXxNlFcxDa10dIQwVOBcZoRPGADkGHyPLsBXB2XF/JlCjWDGi9vutDg4mPQxrivOySNvLW
Lw0YwqUYWKi0Bqv8UZNXD7IUuE92S6qTNosdIpdzywo5Q0JzJ++Xg++XOU/GWpAUV9EIocbnsqiW
1ipzvLGSJ6UxbSMfAorpihrZuavACDZXOKl/hA1PvQ7JKy1TKhjrDcMaKAlqFCloDWTXg0BnFAyY
mvWlGJkx1tTJsTTRkswjz7x7hSQcqcjh2jyUa8Eoj+Ig7/9+Ud4DkO7Hv7H2uHU+u3eISKGzWM+X
kPjBi58A7YKDAwJdCiG5of691+2uM4halPnfWnq6KRJYR710prF5I5A4LEge09D2HVLvLVfAJzsz
qu41hov6Vrv5KZvMJz0EEC8CKgT0Vh1+nGMwxoFmwZ9+Wq8I6OPNnSsPhXqHit67YDi1e9XBTO7B
stVvLd4TioxwjdS0RNYDm2Mk3K8sUmCZGiOGx5vRocVOUJsmmTywHvljoNE3s8QZTG+UXyt69Ys3
7MfbEtBHeCYrxJymTl0+ipZ8xFFbYuK3C7GfoOXW/tj4L7Q1nJtZey36WG3UGKYqXSDvOK0+rDut
LiUgsjvT44PlnxCt2+Glvlz2tC4jOls60nHl8Eib8UG8vse/uorYtKLI+q2dy7tgcKDt+HtD8Bjb
4g+NMefTHKwvjlRnEECh5nMQOHbaf7l0ZOZf+LOF0hjE2Pe1DJISkDSmYhyZIKx6iHl1Ck++SEV3
xx6e1Yki1R3eCxYSFonIDEEbxNAsQajRImSchGJB8avoiyOMBPhwbNtTZuls9Fo3/oMJzx2GovKP
8Bb0y0qTWF7nhpLUL3KOtdUd9jKG7Qnn4f7KYaoY/L91cPB5DzUxaOHAGWDERMvBJX5NYRcuGK7T
Zd3VXZP2okFqHe/Zk76sTYAVNcapHzx7wBYxKbuIugwHUfAT4Dvmt2+JAlQO9rmHwy6umGN4l3wP
4ht4lnzkSfCy3QWndrsqKn8LxGUvzAYauVgnXqPsFXxAPj4YWbY3l9rdluGr+aOuwGgyPlNYf5mV
3l+OOeeEzFQ+B7xBvJ94J7OTekeZMmlsGzXzozZw5XygY+C7GNTvN4Wotw84aB5CH3thT3ecg+9l
yxXTSY4o/QMDQsj63ul0yX4cjG4HabPykGS6A9xIcTOsJAKK+sC4Yv/npYPnHsPdJto3okoB1Bz9
TFcCexVdi9yB0lyy1A7vfN2N83N3pCtnAK3g/6dFRw/ZSF5Bty70Fvp+JECCh2Wv2q+ovP/3Jo4+
YWnXefNyYFi2J/YOPYQE5g+NQXCjaqMK1W1r7sygeItTW6eXVCxQwJt6krMz8tu+2jsWnxgqOXvS
Amh0Qc/hcCW77HpbbjrcL1qL7mxwQ1jJSMr24e+N/eW7CX+8BXZNTkVElwbDRMVo6G8SRwWufiwk
X4UjgiFvzVFGHL8TLEnthYfYLeFEDC8+nb+/XsaqC1u9nOODc+Acdh/+CRlna9YBU80VNpoZ5Yvp
5UhjoTqivO+dTxAQaUISe0P/8sG5hMOmm5IMF737PuBw89UjJR3SxSgTj5r4JKMkoH5tGUt7EvZu
DfSXkHpmm78v+6E5PYXKh6KNI7Bxo8OAlBQ/VnFk05mt5ecRicZ4bZKINiKpKoMoEhbE33bvXeE4
GLACDbR+LlbAthgoTZ5BHXqmyIeGkC7bOLcdKlgtTtzwJ0Ng9Yi1cX9iao09Vbpey3zfE5QlBlnr
4LrF0LAVNtzwy1948bpoarOhWdrFXbWohYo5Ihwm78N6WYY/518OVgRXic0NlXIMzeGigiszNcEJ
Cmni4+HCB+kWJsKLsm4x87UrJ5iPY2dKY0j+Y8Wn6ns+/66sK5Y7qbYlNnlCyJqEka859Cmxj/qa
NyXh5t9MX6A+aju8BhlmwTO23UePk48pIIwfumpKM/nxJ8OdXGoO5yDNuokF5tqfKGuGuuPS/M/m
eOVfPjBAgNOJJQLAO+gx5q7tKKRF5W6d/QmxbUmfrcZM0Pbs64Gu8JpyTqz7a/DftSVKwN0OWk8W
ZHjomwDplyE/2k8S85vCKH+q2ed4RUeIjixxo54h1DFQUxiltqmuICqLhcF/JoHv4p49Sap+faI2
jpaKcAVAAto0z6cpyeD+y6dSdFipQAlnm4FFISQYcAFB/aQB9Wu6qJ2V6kepZSmnnTSB67mrc1P+
QNq3roLcRndy6L0RibABY6o+sMbNhFtaVrY8BWO3D/XzJpqN+vPVtRA3aRmWF8cadkJmAxQ0nHb5
NCHI60fsr4YqCq+KdjB+Jrc2zQH3CalvC/6NYa8LkbOD8MD2odA/4jxfYuxmKYZzXUM7THa6eehv
/8w0e7uBICdptVSDtIwBdyajXG7zQLTxiSFrKc6xP2yCJrfNf/H2Sd8+dLxP4JVcG5VMjggBW4UO
LHOTRaCwa13anuI0oCEClst1Dcz/qnWJe4ubRkTYrjj1JULOcMPzb//LGqiOsQY643q0hdjj+SrB
8/gsSWQeTFM6NrkfSKpXhXi7C71jQU+wQmgumb80yBdUY4XKWRwdNv2Qg0Mv0RZ2ZCvwj/nKVGqS
ZMeZMkzpYZ8H7zQzJ7ukvCKAqTej/CssMkTeofhNf3VdxxVhl6gsRA9lW4+qa2S/c7y7tx+INezG
ptow1zD1kuHU60665qss6m0orkcH2KSaRTNAdXWgtJ/aey2l9gDd56IUE4bI3ygTrXRWs7Ntzv02
b9+O+6zP9dzWFSltog3so6RZaQr+bph+LvQrfg1GO2Pux2G0Tx1k/6TTr1GQh39mhE2zwI4HqGCr
7p+eWnN2ULoE1xBK/g6aJnNfZPApZVlJeCVJOTGljtY3JGgqL/NMaOqfZ/W76CSZjSJ4310M66e7
uMNnrHaxZl8LJ0IhZf6l2T3vpGIT5yq6Cwpe9aGJUPl/uTbXu+Ak1jWeZV+4PHiBuWBXUKv5Xzp/
HJedv9wTbjCALQdjHq8u+0lVzoQenrzdamVVrRX4VTIRvPml+8RI9H9ECSxAYjezRJwmWz6qwUNs
dUbrHdP4OJZ8nPb81k5SK2YJy+0q55hyMqQ68lr6d4ZBs4xsh8fsEfEPm5ewm12+wgXD490I9cYT
37siTcsvMGyxXAbVJAxt3rA3A2yL3S+tNCGbfA0LMG29EA3yqx8knU1QQzveYM9NxW0vN7ACOorf
tfsP0X7bFuyOv6R+zBgewoS8r8fbNzbitOoDbe+UcM501UqTSGMDz/D8kHHueWJ/4OO1irhb3/nk
ZFjbodqJoZ4tfC5BFbxJdzTelikeTyNe30cJjYFcRuNS2fJpszBLK+9OC9spqJYiIfBIJR+fwJyQ
ZHMrAuipdafX2zT+h41xtxMkGX3TUqmkYcADAJbGy4eR0L7L7NCIK6KgTW329WfV7HsrRtZahDWe
ToXGTeeaI0RS6Lpz+oeHr+Em5kPsnJOKKrku3EJ76glP2skRLi6EH9TdgCtJHhV1P/qmJKx1U3VD
uUb/E6UTCXQ2tIMnw918FzkXku0TXthS04oYN6xxXJVSzj9OCkHNjVKmejhDtavkXsXNaZQO7jnB
sG0/hw5umW+C9bhomEOUwWT5uUMZtl0uMu9pEQ/EGJFwdED67QqvWGAeEQeL7aDVQ6VWeWDgRtMY
D9gYPd12Ep0ZY5txDFR86JaBy9sIOJVxOwAVS8DEyg7S1iKxtQURReGeTLy/JrN6YBF0HbjI49dB
7QyylKfE/6nazHJQjdDQfZVgwtvmGod7KO9belKmFOra/NKFyLD3T7AJNYmhLBas6CVsfgXSatzL
j/LKC3mSfGj7IZcibcgeNioZbRP7UzUuJatpEZT9mSPSAmwXbPq4bvYh4mYXN8ks1iE0DdjQLsaj
lVcpfAQnuFSZi0gvxho92jO/C+//7hWTdJI/bZNj/cEIvm5YIdjjmWjDJjyyJ6MTZzZKhUd/9p6s
6Q4//K5JJwgOfmYNoyBd4/W05yMfJhMOikBKaK5xit+GIDro6NC9hZfF4ru9UWO0niWb5LhwC1Fe
YdZaEm+BarROR7N2ErRlc30kjbURty7zLVfMOWmG1WP+/mkxrk35CQkM6JcaRcLeF187FvGdMe2R
nRT6WPZrNKlgDHSzsSvMXyeGTJ2Ltw2g/gg6Qeb0DEJx0VsipGlmvdGMdHVLIhy5D0lGh+/KOzOg
pecpWHVB3iz4HPG0czbTVEINOaBjkCTId5xTut1sXv180+lerN2Jeapzazq6bVD3HOnggELVSPRj
4fDXy019hGfeTka5pKSLBqp1y5YEIoogzuXFNv6vWcVEp/p0q9ELGmA98m6CGZAcDfLxvd1DUd2W
ifnuSmFp0tVqVrFuiKXdFqsvayc9mDXH6D/kMFwucQgHOA6lHB1BYMBJr+ceY24WkAs5dE7HZBUF
JIT52OvEYRJZeh005S/v+blb4/KcoBoOaORbqRt+aG467LdNPx70l/gybGPo2dBDwQed8EZQkxb2
sFHSS2DgRo7YcwyDXQNCDfJdeYizxyt/yeuRjFXFUuYQthMCKOc+UxpFDk3qJaocS8wa4v/yMRl4
Rl9zv0QZCVQLnj18r5doO/1hwexd5L+5bLj5SJOO4x47r/S/hT+nGsd5SthHvVDEmecdEAGJIT/l
6nb+c6HRn0PpCT7uGiAb2pJmJJyZtZpcvpxENRsmSrRU+TY5Yc6NMNdorpjIUUhssrfhvZ+/pHbK
wQg1zjNxyUy2yIUZOJihGneG7seJhUyQZbUv9sm+p5OQhtLFDU8iQDeu9hJqD/VJdm52fE2ynmeK
2AB8Qghku8yxuXxP0rUZDkfaEMqpDgECJAinfnxWyG+5VGd/fjMjvpquKRyRWKdQQYXN2E18eQTy
4c8N12w9y235OxadScQQYNiCrEfEw4G4CXC1ec0Ilbh6Jd9dGCBB/5ZFzPEZqS0+QFAEh39PnW19
RlJver1SeXMTHKoOQdEXFYASQkqwXoQnCSprd1OtwhR5ynuclq8GB9BOuH5HPp5CrANOHpjj+5WT
b/WvYwazhOlBFQ4U4e6Bw1HGRdCGGVh2ldlAEK0sUQQCsGK5Wo6tJ76Yq/NIWE+ppdZ192QHdOKW
CSvfrBOhhafe449u51cRX8EIMraeP8pVZPIUFPln7rOvcCBO5nUpkXHM1MG8J6waswcmyaaLmV8R
mmeA4Ahi1szv3VpiDqUMGRlc6IbfOM28Uvcl2nh3YebuFXX9J0XxwRSRyyjhoHVByZKB/zTnxQ9m
IT5Xs1B2NiYHnI8UgmgiuT6VrwAiP8DsGJd0ud1kcZS3ONOm+A7XbXzoEbnnH1sCTBeXfwwJr5bG
c18xk1yNC2gITKVqHQCZHWHmZP3+QPX/VweXSJIk2uIJYRhyTwFTXakRYkNCB5Xql5ncZ953a8rK
Vj1W0WoRGSjv5Vc1gpNC4ze3cBDtkoueHGMD5TidDK6PLZTB8gk9adbUE8Dv/wTsfuk+CrmiOzmI
AMr0xd1lt2n+Ru/5Xulk+70DhjveMQ4gFOZhNvbhSW0vcSWoGbR5n1bEIxxMZb9Rj0CoNyVMTyif
H3+BLbMxJXU5ZAGMmNWuO0yUvMDZRYZH4LkKJWKPEPR6uIbdV4CqradtomUwAo95nsyrzqnjHoKe
T5UId4muBYv05tOVRNMrFg4c7b/C+/f8mCh6ogosfktoAfUXFYQsM0YrkKj8Gptzs98rG2vNsCGI
JmhzANnI2z6gZ9NWFad7U2tYlJ848w2TVkwVk7m1XGQ5f6DA6PrZQvgzQ/iEqEfJAEEd0jaMT+YG
apXMm5Titl35PyFIAbsgWFTtHm+zG9cH1uqhnlM1J7zOEh15EFBFXBodIIK62BOPxY5A41xwTtlz
nq77hPFO8Cvizym8+djNVazs4Q5u4u52GSKLycRROJ1gnF7hj0IMsrcl+NHzC7xv9AECQjdZtldy
719oVW/wMdFEmrbYvF9FBdXSuy+Xni2Cp2Ze5ufb5bctjg8j32/xIZBTjJDJtox85QGUA6iNxE5k
3hKHwYVHY4u73qN74nsx/1aMt04jBabe40Hz5RChAEGCPoXHs7jPgqVb5HWTUvxqm8rhFfjVbKIw
W3tjRN1Ib7BLFITR1omNeAKcdWMp1Yb9zadGoeHAQ09D7l0Ab4EYUha+RPHD+eH5xsiwL72WWOzC
/ffnlZyv//92t4Yu+BPiyLbLv/O1KY0Pnrp1DSQ6cH8N4WZluPOa6fv68LZobapDRKWKPWQKB+D8
Bpj/ravo6cJu0W3S7prDJOPPwEwTiG5e5DbqUpr4ktoJfA3h7c1SCNyKdTLBSN4Y7tE2PFTutNyz
qRhRs6MJ+gRc1kvjMs+fHZTQc5TM53T2t6vx7/R7YUMT1ijYyRfMugWN1jNDVzyJysnc8s5KAIsE
I6a3+3baNZGkp6OL4rDDiU/kDG3IPi0nirnacg5a9tyEieRoRLHV5yV6WmnhPAdRG2wCKEpABwSZ
LUmTRe7v+2TZ2YJMlLKyuZoGZinBOCrCiF1ZZ2UeFul4MgFJ35IJFRFm+pOR2Q1b7hZugDZxrvmf
Z3HfXAY3XV/H8Xi4OTAK0EDofKzL9KiUM8wkMQzkgn5vQ0N4NNqeq5oOE338pSYG5I60bKIpsu/R
TTxGVayCuM9y0WuzV6rpADmc1KfQRDPgZk8pChgliiWBbaIfwsOrLKbVAGfDwJl+mKhHTqU4WeLb
Gahl8+iptM/ghkoawnhceZDGIiREVbhg4JHCWF51/NZSvRZxWobckBExkLO5D4cRzpe+FngRk0Br
wZiCAE5X52sCL5xihgWSm4+PDv+S590nwohCdVyiRJrBN0U5pp2RnKuQCFIi6QVOmd8D9BUY3oXr
dqUdVUbVRzYAJRSc+Y0QxCYpCgsI/cxfX/h6/tdiuhOnX4e6kcPDVPjRyz5b47Gw12wnh0KYbeMS
VChbDT7PuTX97Hm5m7IsstQdzthb107SgNN64rTSL/AiSSjHL2uYPoq+LIBAls3A8BuGxAltZGRr
zTLkE1jt7bh4VzBFz1ecIdpVFrHji1p4rd56kstwDfiyqxgwdmkWbkXvRjZWEByHXADSYd3cr0MZ
zBPyhb0Ool6wzHtJUiwzfYowWhGa2Ql+Rg8q7CK97Cqhi7GNKw3X75DfadYpz+ud2Fxue6a9iz9V
OGXvmw+IgFCvmxazrA54JCeXfM3i5kYb5F2MNydpEcEAX4+UeTo8N/cxf2KrBffeoCrTsHZyYlCS
fSOkwhfCKq2Pd8vSrvL3JQS3VVbu5G8yMkjVYN5ZVhAQViJ2DW5rZrXYzAoTgknvwKjNWVMMD9Ej
3In7WWeoeVVJaxehnBu76CuQG/GXY331lq8zys2wazpv0Zv/83QabBZ2E+ms6E4oWvuBCHUAMzE4
KsTPuCE7+dEF3TNfgJjWnNv3L6f9iyxf7QpFWI/zkQr/hLEeynqDAqp2XxDjUZnYm2squUPTvcVM
80c9YNpgucqevJWm4o8atraCAKNXtau3Wxt1HmvqKQiZD3LBO/bRCNdZoNtIAtXh0Iw5vl7j0ljx
tNp68nbWEpF3HHqwsEl3y49AhIOYs5duUjPp9h4/XUglSqWr6MCUMxW/epl/3wDn99dANFCNGuvr
EFYKGif3kN2jev/gVH6+HTwsAZcz8MWxDtbO7xJjyIOFgKxo7LQiifB2qn0ntc8gTsWAJVeeZ5xA
v8sKnce3h9ZWEWaauFYS8jNhGXVFTTMooSCbX1a/P2ClbK3/d3lQFnct8GG5yveEF+yxnnGDW0mL
aT3jygCgEaQzxrqEsBS6fx6e5Gt4nUuW2CRb01qTMUmLoRs62KLmCFHkajqHf7NHNOqJP4Ib73FD
+1NYPBrGfPWJBfk0tlWDxudJSRuxZIIGxtTa2x9dmz3w1VhR4Kxv32jcwog7pQW6JXuG1nQ6CsPt
jsO/OZPvWeLts4i6dRChMf4giDlfnyjmZJylOcBN0OFCZWo/f/ryqz+lcH0UXBPds6GAPzCViZpP
fQVViXx0sCjrctaNLn3yvFDp3L5HJf51a56esD9uN0rN2LZeQVpUsbbKiExBDRWIqv+HaGbCdmAR
aOPsPNf3V4x6aZ8Jq30JhpobzppGtAQ+6qYpOgwFGvH1rvHMb5oBeWV7mJXIPKn597mAAvaKTud7
vIi8rL+3t7FkTIolNvITuqGECmkQi9bZMa04IAJCIiYsVpP9ykXYZeamD5c0IIhAG4YLhc9aCYw2
GyxcCbPyclu2wQgur1IlYtG2p/2URMecjNfHlYoV0Szu5SCAOx/PBKUK3YsLT0zIhH27MP9UzU2m
k51Lgnmi9XzQ/X5qDPBxwVNGWfDdUJlwdb7k9nbiTkq6wVpMdrmkR/4zQo58MQqIiOp/IoBObiSo
1MHq8eDxwqAOjGXay0QjXlMA5ul+76eMywEWbDnGgNNfZZBmeQWtynWk6VCJadnkJnZqcJx3I2cO
4LJK/U/QB/Dqpv8iOq4ydr3mYKzwaXaIOdK6cfOuixoWQtCLMwPDA7QEaX0XUQwFmK2Sot8D9Fjb
EZ7pYY8PTqb9BRh6dyjE4c1woDg01KivzoRacJayGdgu9vm5A73lzti6i3Ae2jagagLUKULhzXhJ
cDD4yrY9chk0NSY4O9ATiVBRXcF5XfAAjt0yrzkAat8U+ApOpm+lcruMMn3GUD0moYTnl5R/8K+i
CaPtPHwQnJl4kvH8aBn8l7IHJMV6TMJrMdqBVHf8YcMXVgoqibS/CclZNSpfPcXc5qhpqItxrGYm
u3BC7G7N/qAjihsult1UFKsAOX3OaXnqd/aMVIMtAdMe55m3zJ1W0adN8znpWWY3ogPTZmZhqgLw
6uIZ0Q6IjoF9r1E0Yo/hiKNpxnAtaJaDeRGTQ03yRPVya1wPLEZtUcR24YwRZDpbabZQLIV01Ow8
3q/pURp2IsGVL0kIuRlrMZnhyMn5R6i3mkxsNGXARCTLljVxrR4EHNyJpefO+/AAt/QJLUZP4sZy
O4+OzUj4C1deZr9QHz0PylphFk3AT21G1ltX8kpVxj3maAtYjzIpzuU9xEhvCQ5qb/Xg0y+n8JVH
fOmgSAW7jI1AGCIfc0yCX9tOw/pdbKhaD0witGMqtgNtrOoWp8WgrZIQb/zUC79/pYILOh7JrxbE
4GkveK9cUpMBUSL1Z2xZuXtH/9imQinN4oKIfhQxNI2h+b532EEXco/lLuhtGsvRSNQ0njVXZHXK
goJxmloFAB7LGw8UamiaGpANzbhTPVPF1vqSV7OVsGCcb8953ru/ruJ61DEN9jzVY3iN5Mygdkfd
/TsK7zCm/oGGo/dZRaaxIi4NB4vy17JGbZ5m815v9FyRqUDGu8LE32CM0n4EjRmkVB1xZgDL5pB5
q7pmONTBZrvfkTBvFOG81Bdf1+NyRaAedpuPxygMJUGBRyOiNazAgckmPNAwoXu8YngJ/ZBPo2ZM
g0nGk5iL4JAnoeCijEHUyLrjYXgPKVG8OM789nM5u539oUjYP9x533y4Se2ay/tyYpjPLQ35zBiH
vtQasu+PxrrkKJVbc5HktirUGmtLvqNcumPReDiH1wOdRIBll1MCJlQfbVGjLmdHmUEr521XgE4o
3+MFje33aPQp17bsG6478AXlGt5c/7Aqkp0GlHe8OXZRjogXmkEc3dDVEIcUZbenCKr+vhHqR0nE
l9RReXDrRFiryMPQAWxJwPlzWy+s2WRswNXn6fm62elJ3ig1bMN/PYhly67dRBNGrAauGTZ9QCuD
nFAGfwVRPw9iZiwOtg8dgsv9qM3d9CPcOcexHFszH9Fvk963/IuyLnmP2Gy87SiJaCImF/FhH90M
1TaR5si6JHR6j5qAZbVWDFf788oWb2ifhTEVFQCBktxVH/ZYfOA8z1hcNfuaalAFg6sKSOCnUCMO
V7Z89QmAwwUN2p72wj8NYh7TtKV8fO+41voDU0mQTttRoOYzLZb3frGl16eHeKZ34IxGgs+LoMi2
5fXzJGH3RPzL0Wedm3BO4TEC1ifKCmTySuBVVomttWKYs7JonIG02Mg+yJ39xZXd1wQO2nwaLVOh
Ngk7dp+A1/rt7TROSMW1I8ZNX66+UjDrcGXknARZ3/vwrlmp+O+N+gtRISjtjnIDMaOp59rS5wBh
4LZQoelU3fyNUKtS9ppWWZdkMZ2X+ZQpjFmcCyYcV2Oiwq5+Vnii8jWGq1Qy55koxumNpMuXonll
CJ/Q7x9gMfCSknnm2MX/vd3IRILKi93LVeNtdb83nvrEotsmd5PxveovPXE6bvA8xamKPvvo7f0G
BG7ZnXiCF/agckOdXwP7y4j+txTe6dbqgYD1of/MsxAwGclecFVN6IKV4eIPx6bcb1nAkIUSqr4e
02xCdhNGX2uhyOVvk8ABTYZmW3b2A1vwb5HpImf3fdExyjkEYH5qlmIv/XvgwM9VP10vAjVuIJRA
k6rLhQRZ78k/AclSHBgoXEEwuVIWK5MPGi/ysIlI2oTn/YCC5E+gvPoXBQxJjNNM7aIoRPuhWXUR
RguCcUPBAoCSCVEUCFjz/EhqReWEaE0W0eWH8T7uLXpMuov78iPcdUlulNEXhA0kUKsjWJyqNCgh
5/iBpOsfGjXFR4D3BpfOsCgLJ+RwvxLrlOibq6GS4reCeGZ0IkFOfZmtopjHYRqJUeMQCXSorfN1
nx9h7QekFe+NZms9NVspRicjFhazWpYTKXIai1asllh0nBdb32rYulyz9JvA5ICsa1hbyNS3KDI1
hIyGC9CAEe1XFQ25X5oO9hw1mPGSK3xt+huwIn9mzqZSicdsWLWRJVL4YBpJgbC7Ybie0+RyCPgY
GyVjaS5jEo2rY6x2msHB22sWg8GrbRFB7C81g6ectMtU04Hi77W1/g/dl1eFk0IO5GjiKMIfRo60
EtgQmkgTNlYWdXzwDT9cQ5SCo0m5odzXs4XGLGM21Gd1c0sdfO8AcRLDsoWzQN9pxWutOMJ0Ye3i
NeYFaSl9EJu1gd39mPzSYSBjmZ7/df6lwSSx+mdoOTlWb4Qyi1QPu1QQYUTet/BrWlC8kkYGWl+O
QvzmL4O+x1YnhfddP57AEbEMqFwsFy9CryKSevLFn6ma4k+KPBaxp5VXEbb5GfCGwfei+kbs0iye
b2vTZxTFKh0FAse6QtEBa+YahxYARIZS8tV1bxEBmfe28rh6/AcvHNduDAH0gcL9dGo5nKD3smuI
OkVr3OFQDmagYA5rB8xVqbIV1e4NhQGKzQZ4prqyNAfYaG0j0o7FljuhnD1gD9b11SxHpvXJINMS
gv/H9WqYRBMBWNO60/sMvAmApBGQse9myltebhh579A/hVT2OJbqgmaXcoU5kakm4qJ871J0W7cc
+7cUJ/PU7vvXQhd/HUUedsaGmuJfOuplgGG06cDI2kWEt8So557/y5HELP4cPob7LUhiAD/XHzP7
AVOm0d22xhOQ37rKZIgLjTS0lYSRLvEvwTl60StrYQvCju7LSeeaLQcVqRKCviX641LSYMxPwgwk
vOmNsYopcreeb+pFigIQxWgoUkTq2ZEnCqhNHH6tnFEvpBR0vyBxmaep0ESKQbG0ruEaoqVpj4Pa
NL0G5MfD0aRri5fPb3Y4sJKAyoWDa+VHCLm7gRHR5TtwfAtfCu/QUoawgwFd+3674mTaS3eK76vH
FlAonqb+8L+lGZ1UZEXnritGDVMKaJy+meILqQ3UAU6bpz2KxEkiYEFhNvEnz2St33Exd9Vtc3/o
+ku0IoRzHXX5Ytccdk97iy0DT+04avboNQ9lV4KNUCGqqa7BShzJh9IpvihQjmL4YmaCCi+srGcX
u+luUvORHE1U3BO3sn+mSDrWAEQ/6ODTmb870rZxdX9cxVPWsSxekcjeSX5Nfc+h9GtV4b/nVSgL
7nPlBaXxKQ4yRMXrLkAlDxJhtonKIOqelnz39cTr+ut2HsvW/oMeI4IpUVEkSUKMO2y+bbSMUVmy
+jtua9RA4XJb18GmB+tgRPEYgdaK4dDvYRdA0Fti3C6uEG/Vi6iDhBLV/l+riJ73G1MIhW8MxJ3H
hHfzU1a2AsxIoVkOvTDEWSKms9UmpScSXIdY9VRjOsIRYDY1a+6d7SVADKBVUz6POFdYynSEOYlC
3Ih0d5fCKM3ZDI9fuZkxWPN69uYxP8w/DtVG7Vez5ys29IyugyMEmUxl2YpcBlGt2OiE81C3y8mo
c8scsk03c6uLLEQgldjz241u3vnZ4YeR67mj91xTUJjeYPJXos/i7liSZSJIUIj5fUbwl03PtoRy
byRttZhTJcICMFAYy9HjWtAg8uo+zA/p/Hr1oFtnegs7Ducy4nB4RwV8/F9XLoOVU5WR/NbM2GCU
t1bua4KI/i2ZF8p8W6pn5Az5ugqPKg6xVIfUFC3a6mEzN6fe2aljvvGq4k8v74HzHwlA3iF8KbCq
qeJj05xEduieK5RCFRIi7jNbN9Ow+picQFGZj35CgNT3bM8mDa1j6WDsOgLyQqxDn0CymM2s/qKv
Gu/cB8scjvSHImndB5bhVYGO8KpTJe9nO2XncyTubM1c7u3F23EpNsvjasN4rKx7lDDfoGnXTaNb
yVCieiXtN0x1qQGXtvDce4JUf8nMCWfGs4vhg6ON9pdk/hiyKgE9KLc5jcoRUfYDXy7CnoykWQEP
YfUbt4jCzfBrkQ9SKlGW9zHjhSMjmleliGP9jGlzQuTtkzSNRsVGF48nSTOb0PoXI9qweWcuO0jq
PSKnuPLz/2y77MO8DqmuGSUurmJWtB2GxIRaA3pjQ3UjW9qvRe6cd5JAFFRItzrct7sDRreTI4el
w0Ychg1J22xqbOUUJtMOIsLD5PgV+lKV66Ixd9o5FdfCOgeD3+g/ISJ/RCVnWsdedsKN4/Q5A5a0
gIIRRMCxWZLObHdECs5BjX1hueOVhLtPq0wl8TngV2Sz1XGNHfBLS6KrqXQiY/gwAXSI25eu5v68
IzmDmxQoJFg8Yow0K+9a7xWV+krIzuZwjMMVv5frZ5E8yD/5EgsdumlmOCyrsFdJYf4Lw8pJiLFi
0znjhNC9czDwmkelz92eOi2xlaoJVNrjQMHR0MBAoPxQ5Asnm1m6qRRBkeTxIBt2+FBgebqjHF8p
M6uhyTzidx44gutUL60RHr8IGG6hbkPZUrpjQKxUq7PaVSGz2sAlCmy7FQcDqx7fYWvswX+mQoww
t56BOVuARTjWtZj3pwUZt7gq/iRyleK9KPzDfdpZtiIFUe1pCZ354zNiVi2LK+neWdpclpCT6+B9
Z3rql8bs17KIojsLr5ZJRnIO5CMX2AeBj8fW75GqL1+hN3mjdyAksmUc0VAmyTlWhP4QLwHx/682
mVgtYGG4kLRe0+uoqVt6nn1XN2e6OArg/fml+khoyL/Our7ypiZ/PwTImD9i2DyydQPdK+o6vlUf
bLT0HmjrdSSrFVQ70hS89RzQJwICCdm1d4YdZykhiq+cO2ZyNFJI9+qvRo9FuHe9yEfSiiFzujRA
dTYxLxrkA+3W/SOvMXTcCUzhIlXRiQamfd4fVX+hs2gWXLkFoB8dCLFQ9299NUKgkuJXH7Mf9Z33
mWX+e/rYvbdiCulc5cY4kQCjX0TSXvxZ0EEroWZ6FjDUZmo7BopuQGE2IJSvPo3p6ynfu7iixTLW
46BHU+8+3QCPOouWQgxy7lfymDo9SG2xfF+uhtNCShWeVkcY8T1wrpSewG71OEDAosb+QGGBauhT
UJGl+1rH+rRCw1h7G16NivXRdy+J/sREWZuE/sZBS5io4C5uSjVpng6H+j5kGraTb6D3L+7DnJT+
CQzkww358guDbMtfM1S0C7r/ukruYw+D5K+mRlG7+LcyF5wmUlDnXpAaB01NITjK2nqGmOhlC6JM
wn+qaJY+8VpRbAogG/THqi5wpmjUP7O+pTsSnvUwgH9XMqqkbHL/g30AYdr2El+HFSbdbHszrq3Q
4a/QO3ItZh7qc6als/ZO8Bi9H6oF4j9HdMzsJVyL9nTWUquWJRAKM45Icp4bWjORyzce8z+aSEhD
TsUwZErKUWv82DLcjMwiVXQFLwY3mJ+nksZxN41KTTElW0SM5JOnDMGEoNw9AXFB5zumRWueqlgQ
cQE7HazOwwUKfmu7K+AbivzquqbRmN9Q1Ytn/AaeQMK5OfmEoI+QOzaYvcI1WzTjS/ksNIQu/EAm
gT8dImy2S8IdjoLrKmCPhir/j/4fpFbobRp1z7CAJmghr8OD/nBfhSyYgrja3igKVfd8jLGmUs3u
2Iz9icjEgFiaMJa0RONbVbR7pr736dvbJF+jYjvd2Ge7lbMF8FVBs+nVqYYA8X1MwB7ZjQfOARaM
vIItleVg2H970NBXnI6tCodPhnOdXyRxZAc0kaYhGyDqMw4UUN6YCFPs/A8wBamh0mXxCwLJ+EFZ
QvmoG2RAYTMilxEnyro3vQwZ/whfwIX6SjhVvs5INLX8KMbOGXMWKvCV5WS/ps6+LXnyLzJmh156
qjjk0RbA5QeacnMMR/+EhsrfbK9QtVbRvNKZ2jr+0KDYu+e3wlHAZyhzZXKKc/lSY5kxsrmprxMe
vM1XqYrHQUYSQ7yLmUObuaSovtm68ecpaDkpXpzPbghmLO5j6RP7wYG6jG59O+5c9DmgJOYloV4k
wp+VrHUqKByUWIiXHOtRcCsf3tWdwC9Y42sAvhQE2D0hR5fmwlWwwMGrRm9p4XSBm/t9Gx4qJXh0
ECSonTR8Cn0VG/J3WElh/3eAo9VKYBuQ3zvfN4wzah5xZRm0RcXOu7lUS3MzJWNriZi0lpjf0e3v
5EyLIG1iPa0cw06Zhe4o10C9I/rSDnlMpqeWF914vzVrm0Tpz6nYlQvhVXTxweVeljtOHz+BjK6Q
TJKE2fqs9XuvniL1toi9ytz755kl6y5s4aX1L3Lf1bjh2AE05sUPYIFfCpaCkVk/sgjewWHwDJGW
T4oY5HXfwz1p5sAGOkoa5v5OJgCW/hO0tZGzZUMlPRm9Fq2vCloyOz4JJ02drLG/ZMYXwwXjekDP
7F0cP9HPMtFBVzO7UFrDTSSWRvtHj4GTc1dOOOCp4S/+t0i1FblVxD1rHluj9FxBUGc1t4Ny9FMf
kAYNQeyMBfr4f2u8cgqrRNpZrwSFRXG/oQO/krbVpL6XAVQrRjfXdyJFoBweCXYGelKrl0b/G/u4
I26IgsxwmM1Kzs8ij89R/QR+InXdWhNG9yZXV/6wldSrXWA+tx1dX+EmriXZeW75D3u+LPYRk6s9
/Bouubsls5q7M7FoSWuWofy0nQ4xfuM4jYJG+epCnqwdQp+0EcL81R7xtt2Cf2wuq/jlXo+kOFpP
OFtasAhkiviUlOSbWqYHoVwWJklhk539cEdvnzsQ3GfVOZai3psCXfyw0t/RYgl2vu2Td95C6p9X
OL6t4IgJDoLhvLklVOk7MsPatqSjxeDCCTnkol46azR6IzV9/L7IM9CWwzPO9/6yGWTdWgNaGUHx
75zAMntWsbXsAQqUaCUHNXt7jitq8hdZMgOvXXJsOrT1+Y9M40fCJ+tJ8AT27l8HFdef1nKhOQUI
/D75F+XMu7z2a+1nTVCBhvt5r/d+HXuCZVIL4QNAUFJbDubh6fBX0eaO5i+1OypJHRQ1n3f1dzvw
7Pior4JhhGRPK8NANRqDdEoee4JEbdfzEKC8GPlNvSDsF9QsD1eIiF0C5Aao9xCjGYckqHqzQbV5
0MXKAEFuFkV9V9IdPm+UQ1xxZIXZnkgHSJaams4XreNC6+J2SzT3KkoHcn5FA0sf1iH6DBOrFug4
iLml6iyeIyOrcy0SXmXPUJGh4pIbDnzL+Xj+k1d2PrPWyJWKWiEIrYbNf6FJM7SZB3pML+EOGDUU
rDX6d+LrNg7QKvgFFrMUpDEpryTzpWK90VT9ngF/VbGyfbrTt+pmhA3vsR9QRhxDLh9sXxcrET9u
NVnQj+bLHrw9WQ+1Y1GVQI4QuDpx9/M/jqlm9klya/pU3WwBl8lNRbgldrHlHriSnDX+wvoAeLfz
J0o3rYN87tY3eiwTYYWUBvUz9t8BA4uW1hzXK59+3Qvsw3cTo7TpMfEwxwpyO7gyQ5s+UVYJfn8K
1k1pxRQRns5AkEdKg6aauMSU7KBYaH+KspnIRxDsFIO5FIJ8cetbV8dJ5Wjj1ENWV6SvQWDlKJ9J
w0djObaRG+GC+PKqbmRWtkqfBl6nxBYBo46OauijJnu3N21rWDJbVPmpcKexGxWDpjU/Blyd0zLq
XmOKhzcHtI2ro37a15NmT7dlROQaUlT1198uqeiO76JabfQM9tYoqtEIp8yom99Sgn3Ky/3Lh2sC
f3+hhfMv3FHfR5R9oMgoB7R0eV/ey1/LEBOcOwW1sfIWWMEitotrlJdUnXZDIA5lyk/9j2bEojiF
Hz1xwhAYpEXW7bPpJhMLV9KwiGYSIPEwVkICFptJ83iEMEBuMPgb3OCdjU0JuCdnGDxnphhhru/c
RBedDs/k0i3M/DDQkGg5v+OXGEXE7LayJ2oQS83S5rbKE7Z4686RTbHkyCb/hkh+dEVXQ8JL9V5q
nRM02O4PVFvAoohyuaoIcG21FmHLB4ypZ7mHRW4qJNvSgyUeAnbHJ1wqGLjpdhNQ5Yq5B2234NUM
mEGL0nSKDKre5Laj5cCWG44CotSJus8Kp2uuBDl08FJDmB/yPWABTAGRm3s/AYa8G9XVrFCXsV0/
I4bcWJtgiXs4Gmc0oHMbZRUUBHtM26fWwJhtlVXF6EpVhKwQbqpxhwhCtJfSXESDGZgHUSnn+32Y
tn75gNP7G//oAeYEiIpdF3rg/AkeP9y+7aWQ5kv8u9V1RShrD18P82Zy3bOa6gbaambuQ6hdJhrk
aYqdyOvjdZNsyrm+necpJ0H1EvQwwHDQKV8DYfXv/yH/G+M0gnvUYvrzpBpEaJKV8koBJOUriR84
Q6Zqni3o2A9kx6/HxCJHeuHH6nvRYljlrheHNoVZD5P0SBuiuXRy/V1XW+tV9WBOjmfgQnNLR0EM
SksNRcSZ3z6YWGqfZDrGCL4NLBdc3fJFQWy8cAsL+kkKSscgWkZ8EwVyQ5pAOcOXkPsipyJfhnZN
iUZzX0meduU+AC4+P4iHH/K8jv2iLurSDod5P5kNz54/bvaZs8linrKjlEz01nJnOJI7A/hIKbBS
z+GzBNtAQZBmfgI9eH7fOzqL4V6Oa2/WnZUtKYxVPS67YpYnlxoq7eyH3eFk+oIdyi4PDn9/5ZdE
rE7HPwwYsIYwjzN1dGR/LOr66VMw15b1N4j/Ya24z+Qpaqaxr38GtMOG2P7TWrzE5rLWPhmOZYpz
/MvSI/9dFQesXGJHHIujZzRw9/Cjm8PG0U3y0IXWS0HTCUVvNFq9+NbG/CJELshHKxEcN5hys/PE
uT4zaolU5SxnFuS5CAM5GeZqPDI5AMMliqYJXPK7qvdhFlH+/ktdM+a3J0bAIwbRuPDSHAaLj3u7
KgBlslX4y5Gd5ZAw1TtXoVDzI2MFgf580xCgQbg7nSgvCnGsgVROTs5OilKlT0n3mwD/zNYaxXM7
pv1k2ZcklU+g2GAy3Akz8wJ6hbNWlxIX5zcNoBUwPLZjJkhBJFOMhjg9Pr3LCCpkxRoi8MEKseXY
8ubwImgIbnyWDWxNclHuyf3S5WYDe/T5BBSsDwH3w7cyoflWcjCRTpFDVKLFwQSxec6BLwY4Rp/p
fRwjB5xikI7t7/DwkYdL+rPA6se0Q7Ls00+X07SgMPbUBOwSJGBgdgGrIPTQ3720bFOIYqOl3qpK
nu/cZAFt2yuFSI0O0aRf0XYygXwc4Rb0XiNSysyzldmE7LrHmZtmxWBCuchI0ETGfaZwEtqfRsWd
TWvV5pJLIEgn1tcfCE14f7PbPQPydis1KEATkMGtgEac51GikM7zbcuLYvDCe0bchg2QjHOrFTbV
nILZ+tZlDmqBI5QeWFm21qc6uxu8mzN7bKHGqrv0iqUgZJkfy0K0Bwt6HssBq7TvVHQaIg5pZjhv
Nu/fXkKE2wF26MRMpU0S5Mss1NlWVYp/rChTy4UjUd54bHZ3HuY8i7RN9BipGKqqmASPBYnT/jQC
FBrHGubvXF6ZNQPAF1LudwqjbFkIjYqV9jNOYc/b+XsZNjEnD2UAWA8Ke0atCuqV878D9PnVeolK
Us2D9620BTaDTDBC2n47Ab/jVnR/m+UQVIwRBtl9UbF0VExvYsXyZfS30aOQn2mfcWvaROmfTXi1
Wl1Pka+VKkom1tRiG3TPQrnfIgNcdDRq1Z7zmFP53VtZR+otCL1eD5aHgB8wTtL/PU0jmq9J0aFf
WX8RT//cTdi9Fo2s6cUoHj5rFEkHVW1dJbGACkEokAp1vPxAvBpXMuisr8Yb5oftkGSW9VOBlhS5
wTHcIHpuLbk4M4H+QhQVonYyBUzspibK+NAfBJgx6zfxdhAB2+3P5zbo/AmDLSWnDLLGV/kzNWtg
36QGsWrzym5vaPhNnE71EMHcddaWPN8lavrfp0IIiACsmaDRu8vaSeZEfj1KusFbUKmHXjMbxSxz
KR0kIiMzJBRO+ydNIdxTX1jn9Vccpf5rMykT2k1ncIvbUiZiSH+XD2cndmSUik9uACE4OBGhXGnv
P76z30qwgoKX6/7mOvCLj/Z4jFh8DuwWX3ji4UqWx1gguC3/hbKgyb9XhEQ3ENpedL37V13dNeq0
ztdxUJ5mZL6xNIyD0nEEMosM+cGj78KJueRdmnPcjIN2NsGAe/1x0G89crL0ur2Iiu+nAxAHjGzP
nehOD0zhm/+P5fodDl2lMB08gFF2mWb/GoMfFdk7E9vSAwKPRI+gEsuMrhIZJdMZJUK8BbNTMzLj
3A/7eju9ID6hmr5yBtRhLnWKjHJ5pcKr80Kl8uz0AEfzpVtqcJ+Q7g/PB58e1Qgki7gsxRctNL6n
IoQTiQ0lx/RgvTRhZUGiD3Sy6rmOhZqN1unjKlXizYUxM/P5KRmA7Hup7e1/TPpX88C30Jr5VAnA
3YMkqOAWtVLbBr9NNmTz+pY6ErSWlE8j9Q2q6rpMnNXFSETC15XxNlKaNYvjZuF8fgeSSrlMTSO+
ugseaHIvHCD7WmPEjYYi0Lm+5b9t7eP3y8jzAs201oRlXXxnb+JmHVKgv2TNGEaf0LG4Nvq5Rg2A
SF2kcV5ASt5uBnKEgGqx+ZDadeoCLmq9aKj2ao4Wum29oul7m5bbBd0euG2uuhVmdW+QmsORxQF9
ngW6PH4rbYP/swy1IhZp7xJgmpt/zUNl41E9l/A/Qf9gG1RZwsJExiK3/SKn127qCgrJA4G5TP8q
zMxCyCHZb4jDWDTclq4fqA87Ex855FlQk/TtfQ9DrSbR3yl1qNv8Pid5vxc0prQ8EF3uOARM6P5H
iD3FvZRitx13mQ9lOk0wFI5TqEk8en0dR6Q+CkSFsvgJGLmOkDJFMJhKYPUl6B0OhUiSHH+uJCyM
qpmg+/looaSse1UDYCPQTBTg34Dh1HvNkJDFM18xUFdrSAY3J41/j0P9K5uyYuMHN114qSLX1ITB
KUoEh6G/xLwWM92STOE9+Hu0xL+h7IwP3Qd+pj9AFlXzpxC4WCVF4j9FFkmoZDLhNzcauEUwwj5m
ymQrk1Qe+22H6nMc/D3mfM8bQNrgz57MwqVFdsInuGzGIDfBsCBt3wD5aizuH0/5aO+JZ1DktHzv
3dGRa4BEDYwgofX2mBEt/5PFCAzWMobN5/fAwvmtETVoQE19GW0SbRh2VPlXDuBm+pK01iqHRjeA
qh/7ezKUDwT7wXYeF+9Er5gQn3nO6Ax1onmWeCmby3rsauQ/FxFmLhie82rsaj26k9Lk6vnEn94P
+DUB3RvmFsqBvoDUEbCAZ5moCkvbPGmmT/gwcfMUSK1/oj75XOtNUwqNCmqO+kYJm8mdk39LrhQa
J89IJJHSFCXmDs4y7I3/OWA1GK3mZAdPj+agI5O++w80jsDlceYzybiV9StrxtQfTRxYTzKcqhb+
QiKCeRTUaXNMFtKHI49baWAI5911pDrhkS/RlrNw6aGsY8V6HnBk5KyBUvn2VoGyBkSyly6tt/a3
CPKR28EXssLrzZU5yC3iOuP3kJDaG+42mfu82ArpUa5FITQunRjVpEBn1NOTcPtAOIw7Bx81kDfy
RQRHCUZTh0+JknyDzwh+/yq1tYVBpw6mGL8VKaAZHtGux9+MGCGc8vFVfiWpe7cRSSaUeUbk/pKq
X6ET01fOC8dARZ6ct98DfK11RVgpD8JX0Q1ZBWFLbm51qvvQXnf5vE90OUrIr3xfPvpvxlVa73z3
KNKc331XG15hF5tnMzmpfXq5rgm0ggxR5frtApoXKAguiTUPEBRSIjOO5jbj79Rv/6PfaItUv6/u
tJMrIZ0MgX850gQXJgbaxGM8blu873GooDNUnuLIzEtLZ9MCeF0aa173LehvAz3jFr5Xy26ieHUR
8Kwrg8JAya0LVcAm6bkGZXCYTc3XeGKeywHaRQjmJP9Xt/Y26hVpxn42vACadc7Guhl15ps01KWg
JYn/Iui/rFrPBU1SxR0+LA60VuvJCLEFGi6O2oyHJEwFvYqQLAMAQXHjs7O5LSx+9zOdlfewUZ2U
ZcdrXXWBqEXv0WTREBZEXl1CFfJV38KK70QmDnLeJ0WZnBKpipIoY6K94b3n8v9wHyjWOzJqCpzW
dOGIvIU9CB71NYPyAw+Ev/tFFZsQ2Lwp41jz3AbDLAPdrSAsWhaR78uo1qr/Me6EyejI68hZZWvk
IsbcDkJ8ubta96CsOgCzrVLlCgoiBUCx3lmXClPboCxHBF3dCurcwxCSNQ4RaGOR7tI+slbmoafK
hCHFPNBue+YNiafL8KgWgBJL/xvj11qwoUtzud12P6+iRQSlVAFOiJTuCqFg5QGEJc+a3Fge/mQz
5XvtZqhianafhR5I42qz5Qo6b9qdn1eIjTOwe7t6RhtQ9pbiAJY2pweglpVAPXReTwwWZxxS3kjg
VSORHzEl2aPel+YPziPUShv1A3Td40XiJXBO6gFwMgDfvXH4XI6nfCX2/yV37FODdCYTLVC/RJel
N8/r5z2FIO0m3E9RV3l8UNITRHAHECJozCLSrUFgiF1LMwltzdGUzKL7WTH0/mB0G5HKz3vC1O9K
7N0d7L4G/p67YHOSeMxaG3uBm6KowSTSMfNVIO4sVDb32cnKsaD/wZO5ifl/SyLapfQKIj3e3O59
ihZV3SDTDx9YVjL0tyIBX8RrPLq+kI8k0SDUxrAax9sYEQ6Zulhgu/mAlqtwqH1b7Uytc8kR+8/S
rfD8mGWTWWs4X5VM2I1wDwCKdUvHDkA8XwJP2ibxktfauKAWmna3/4771wy6EiFLRg/5u6kU5z2j
2OIAgYKcDbgGb4jDX8Pu1URkeM+2eVlCFY/q51OQe59dP0lYkJ+g4wOe2DjsHbOiAFbfPPdpWtJ4
QEiVd0hvrPc8rSRG02IKr1ATQg+a2QAc77FhhuYSZnbHUYzfaFYKXlsFK2VafEEdst9PJrAYMkcU
JhxmjWDrVWGzRiiMDzqXzZgb7aGQpz7rfH+Erce4OA2mZx4i363qQYFjTBOJ9KusQGX2XnFQ4XJM
TYmavIu75GUC9s4peo1ewfDYypbuzBcbxCmlAv3+/lwQ7Iq1P7x7qiBr9SOaZZ323/TrefyNpJEt
ly+bn+AsGeP/mec4jTsNV2qDrWFVlA1GD/sivi/pzpTUY1k0QY/jkqXxTp+J4VGcUwXwqNA12HB5
EAStLfBDALKZEUiG2F9FOYO4kyrtpRev1xywaJuQJLNbfZqjNVEJh3tQSo5hxYv4Z+2bo7i8xs4m
JZ3Akqyezc63JEVTNVWmlcN668xXwXk1ceUpHP1lh1bHU/Mzi1AToMg85k0D+TdgNN4UwlomFIEo
tdAdsi5r8vFt/09nUWR/l1MmLHDUnFbF3E2bbrnbfQfhOypQC/DB0Wm/xxSP3k2ivITvGbwYQCK6
eOujuW1+LrorSeaVMJQamIS8pFd5v+GB+4PcJJbg1vodetLNBrqTYI46DGCS8zHpNPhU13Ofa/pN
F5aiId0BIlUeiJuR9onxlhTrxSG2Yb74Kb0HxYxeG9L/z7r2IEUY2ycUxHaXc2Vq27fMGdxV3HH1
cW4JFfVYC/YquoIxu+Misc+ICj0OOmsxqK9svZLXzReCAfX9OBYi8B4V0FlM/IFKLm1LwSJh9JZ9
3in01ijrHj66IBkSu3375z/XznGL4hC1yte6pXJn/jxOJpZcnAc+bVY9w1cgifSQjtMp1XEm2j2Z
miPpaeUN7mSfPJryZRqbaT/5FSTI7b8MEl8+dc+gI1YLvrJr8v2p1UnE+kdlMoizcoTQnWeY9kjy
Dq2FTHYFV7V9Xq69YcsYb2fa5JG5NvgtGphHRpgDs4eyryOFnx1bRBT+PKVfOczYXfWXo/d+hOX2
oBLlkXNVcG0jC/02LJssvbZp9e8DLQVLJtked51Fkup6g/s/Eaub8cfsfQ9X0S0wVzZZGyCP2QtZ
X5psau9p8zMfPXAD6iyhcHjtIhuXv/T5OjlFX23YrDnKNxEiEHamlJk8RCADgDJ77EQLQBTGXBEL
rF4mYQJSV1OmLiqGlnTEffpsJQxuOyT6vHnT4CbgNWzcBqGvR27HmqRXMVnE2vX8odW9XsiGTXA5
QoMV8uBNZSX8DRFxrKBZ8Brtmd7OvlwFDVEE6NANdWE/nsJmj2TPWfS9zv8XLwdkODjjAzfXEUNa
IexivbcMh8tWiMd4cwNkFCJCYiXJ0jBxLSvbGt4VeqIXKzRk8j/kdclumqlnHjEQVIP9T5LPPETW
fHplYjnepu9pPpKUUccVjMzTMvC/FfhE+zFiOJNPB+4FdPfdBlVJwy/tbreXJELcvxSW5vlNrvg3
nWbD5sU8Hrq+2y8/k61mQZcYHIQto4ZHq+VTcNbEDye7aOZa6/lx7aUQwHZAAJJu9G4w0/qckh0Q
g04lkxCvvF1Fo26iNoebDuOODW9MjPdppvetVToSE10Pj+yHupFiFmHEl49xK5A4ATmCX1k1Xorn
t4m3PG7CKtsiXNpc7wyFq37K4GPjanONlijFImHSy9brEiKN7k76bSDCf+oN/Srdl79+7AzQPhYk
FpF3ByB5Tg5g6sSnzaEOFAI4oh920D8YOKcsf3pxgGt7Of+ASMr4UHnLrubSymY1/2IASS+7D0u2
M6xuVUxGHHCIx4N20m7QHmnadtql6+Zb8aaM1dh6Xt1yQuCGRSKBi2jmP9uGozEFQc8Km4kPDAJO
eX93oZNxWEitkEicXIyp/k/uuGv9titcytIhC+0JAI7s9fWO2aoJoGn/c/q1/kpuGKMdqZLwzbBp
3N32Q+bLCWxgV3Xx49jOfnMHuRm8gemwMiYSsfCcv4PLa+6aoURKflBR+zYk6mP3sZRKrsHkJ/ga
e2XoZEM8EPysRRl1owmubjlY1uCPZJoJAdc26LdGG+gnfN7VUmVzDHkhUdmZM6raz65K/BnwC2OX
eJmClsxENkLPoi2z61dBdsAZ8phyqlvoe/q+UYHeWmW+srZgpRjO8Uu4PvZiK+cZ0M6gw3ZRTHst
Ncjr8Nxa1LzruOOMHXFP7kvs7PRAwe7dlagSyzEshSspCLzMABkZDXZ6dHTy/L0iKe0dnK3jILEj
01M8dehuf4IUf4xw0xxP8AIURcLrJg1efOYjPn9fKGQm8tRq38JLpy3Qvc4gyIjmkj5nGOISnOF2
zIUQaWJ1Px/Y+yYj1o3y24BBJUsEjdBzlozn8OC/vkOyvXp6K65ODvsleDVtPYMec/+mBIrDHziT
BlnDlLRBYhYcOgEvtsNu/2WSk4BvOz7Fk3c9SVg6K5/eW5d29acGSYEIEWnjHSFXdaAp/sXaBx+o
5COjmbYeXoZObUL+8yN/Asn4P5Mi61WYwojjHOXmHAQaXyloW0g21X02htyQN+EIi8uUZ7pCHexh
S5vNqqkEYwHPzVcofdlIUPcPXV13sw0eDmOPqumARACG+8DSla/AOF7v9D/NjR+K/DlCqBDotOut
ily/1m1KhxmrRd3qQUEt+JKmSyt8HRdj5h/oh/XTptNLmYYANoczIf/tga3AO2RfMkUwtVGMerZ+
RbSqs11VrE7TBxwEptlibjOxFEOVHtt5jEaPljDXiiX23p5iWfxEXuk8HO/k/MJ4txAi9BwXMY7P
n8pmYI46NbEKfFJn2DZeRC8xmPIM02Ivh2NgjharRI6tNrA/FqQv/y6Iu9eV98d0FCZX3qUI9Up+
hQB/NxPkoZBn2yGwGdyMYP8FBq1/IO0Ef46BBJtFmgc/oFqracSFJZq07NAJq2n0bf5svJr5JQrV
jLht0G4AjDN1vI2JaoJyl5yVJkLDBLGCN2JXZ7IQXvA+AxWvS0mzhU/WI1c9SqCqsxO8C/uXlFCK
9+sN18p9BTLJlz65B9abtHy/4ynrfcux2r+6HV9jbUPJGtklMLPRL+Svm404ZHiVEYTpoBr7TX3c
LefId9fwGFspLlLqoFOMFre6z0fXkoXLHe9t+gC0cxWsNqH5MJ6/bXnFkfHC6fu3hvcABNjZGeRz
ev/aIdvZZ7IDtCAP3zXUwaaQiPl0dhq+AqNdqjfTCggHSAwOXc0VLundI+Q3obSKV2z1VgE6BNgP
e8QXuw1a4eRH2KtVEtydgWVB7ohknqGdwSMOhdqp15PVbu9V2dTIgP4iXCuHdkAA0Oe2+dwZt/HX
gH9OLY+I9WsmoMIufX1LC80sx8Q22SYu2SZWr3HWdl78SRaRxeSLT9Ta3dBiQztRXnkc0RK/f4NK
abciicLkHmuvfte27BcgXqNDd5fVrbZ7osZIloPRHyTURy8cmDQ3XBVndgP1X2hr1glZtxByvVtF
gw9a7VcQnNvphNypX+HaQFCJtehSgRkoUC7P37nyMD7lkpWijKigeegErrj6Wprg2O7IuQveU6NM
eglPk5k7xHAnmNXt80teX/V/LcMlLlNJdjSK+SK1bNLKwQbQt943+J7SBfdN6K1gJfCuKKGlkipn
skjKQIg0TzoteAFGKtXr60azDH5tF3Lry89Eyy9GHdiVpyplq0spAv49UhmJ7f1cX++UN9DTRpC2
4EZbs1nOIL61AAq9NjU8R/EbREX2sW9yjIvq8CEChVOPE89dsO7ggQ2FQrdxrAGZoHYW1ilKs2bX
qnGhJxf4dLiKo4lkPZtzIldBlCHzGy6dhzIvBoksk63oAPjPo3wPXtruOvC6TVQMwW1cMjkDQKZ4
ZEEtclox2y5OjOAEwpnI2ig2kKXdjfM8fPpeP9nuZojsRSlXHhj05tu333khwdOa+E1tHlU/N2kD
rdpW/zVM2gaB/n761auzgHeIDhTzBg5KqXOXS36hGr0js+/+YsCUOCHE7Rm6tR4CJgJMyXw1Jh7f
Cb1y0gIuRH/z72KpxD7x3rixpfP31BuY4vKzEa1DDI5owAXjypKZ/jUUtsrpizbO8mSMgZTnzr+n
uXILU6BbwlBqW1j7QFwe0a1JK2wgPfzqOEznpu3O4uMcD+WKJZtJhZGGcJXBXKbjqQsWkv6cU978
wnN22cq4GS+4hVhO0ofmZfDzk9sV1XBBHQ7YHy6ZkB0h2Vgb61VVgfI5vwJ6BcxB+EuRpBksyjAk
MIcKUqUiRZMKxTPVUOBGjbkE/0YNGl5JS8k+XBN50DWk15ldm14CU3ryYAHYGLRvf8KLRAmbbbSw
CpiLT+2/aLrHL9CaNZDKLMy1t2Ut5x1Id7I8j4M9n9g/2gMpHtOKohgcTcQ1U50BzIXZvjHPNF/6
8+HLBC+pmvHJDQlImWqnFfvu+7nsvf0L25ZoneMoIrMar0WLW1gzGnEpXUUrCv3cJHY0FVb4lUqj
557tKPwbZ0ATmKPTQAvLxrrV8/U6keAwEVgvh8W8QENAuAGE4sYK7bWn0SkDj912aRT5ILpSrdms
t4PhmV4LkqAQ5mxEMvjQZYZpMYKPBVR9MPtJ8Wf9Rl9cBwL8J82Hk+rUIuP8+Kbph0rq+OXv1E76
nxsmveuwt148fqNqwiqNzEX+vcf5+DLfW+xceYMaHHePJ/Abs57t3SBgX6N5OKXXPLRL3e3IXXmz
zJaCoJ60rVNoIv8cRCJ/3YTruR6j6M2EPqzFwayCvEEPWByYZQeaCQ1dHtIaGps4Y2YIsKOltIUo
Ji5aAMft06aESd8CyrhDorAXbwei8KamH7PGHG2BUyIpqMNTqeaa5qIsjH7NLpoXGIOWocgJK0bH
kUWyfRXK2G0JYguYt2hsY1ZcJkUSsFpbYJ4LVzKvfadxKdPY1Xv8ipDqpbyheFQcHUJFovisHqX6
VC3hzNRgAMEBtujW4wCt+n6nG5zYeSpVLyaO3VME6DVQM4YIsWdm5NCmfCPD5pSeNHRIHRqgV3ya
yuvVbwWigbNXeVMIIMFQvBSRaCeZoVcjzwaYeTuav4lHwR2AosK7PcKEcFrnZ2YbZ5nUHtm6NMkS
CVaYiX/yXgOgqWuijsYsOh3df7LNjnsYOlrpLQSRfZ1tRD38HTRtjTJgAmYPIDT9gP7wSNq2FYDH
+6vs+wjAsOjGlZN8QKCbOVHL7IJgspuYcodsYjZjYowrqZnILliLMMUqWZU07kInqZ8cPcew/141
oX1Wf5V5twESr+I+VXEUoibiwVXdoEOd30iNGPAc6p50XdMhumyDmEt5uIYdzRNebmyvKGWBq4Z3
HK0DETh+nap6FlKiOipUfDycivKzYdkC1GMt1vSglSH/iL59V9NLsI0GWK6Yh5jdEPgLspt0/hVD
4W/vFfXPx7eKt2A5Ue5StZLQ1dm9IuqJf+j9AxLQ8r6+k5d+7GMU1v9UWN8+EYIgPBWa4aJttTY0
6pyyLLxCWykU2C4Pwv6tgdMax9mkjpc9Kao9VhxcDsYOHJ21eu6kB316PBN9SFylBzcVvtGKQCVg
DI/2+ylBE+wN+AgJHcuaFG6/cT8HVUOGdNIQYSSmZubVUA8EZlZCinOBAHDPT6wUyJba1aMFtztX
HbGDvaO/1fKRkA9uoUFiRM1yr0fTt+gBSwEY1yc0Kz2L0JqyNDj/8ZJKSNIVIJqkxKwHmbD/ToKy
JvSCdjZsjXmmaP0DR3DjbwC8BycpsAKqmGmbMPgiHyUusvusEmhmv9PUHipbYjI1jm7aXiYgjUEv
ODjh1BvteFi+SvQwPNJyU4B3OxsHJxtJgKVi8Yl9VuWOlwFBRp283Gz52FQiJ19ecRqmHWwJ83iv
Avzx6eeHS2uV5hXM0MiW40GsnlZTlqRjDpXqUjjARF4pe3dj6qbyqAPQxiSkjNwFfPRO0O4W+i0S
38syxsmwi1OQifJXkmLq1XMYFpmtghe5ohybPmJUF+8Qz7m/1j8BAg7V7fATILvpQFjfgXvau+ID
sxmyDpADSS1ZSFeY44iPAblO+8MoqXQ5YKzX42jr6vt+LrHWB39sXi34Sbr+1fBibzxMgKqieEuh
45qW5ic6iaUu0gkCoL/N24JtARSVL/ZpBE4f6qBwB2OSa4WE4mvFhDjudKykqjqnnp10bkCIAsGI
zl0kIv0wZJEiajrP8UcWlDZcOM9JHN+NksTX2gnLq+GMrhn4vRl8Kn0fyorJYJLMyXc63eVaNyEB
JygLK81BvKgvve5XkfFk8m0K3EmHZdErtweb3CuhYdzlDO/lGO9YVE7QEt4yyKmG6wZ+UbXjO6Kn
Hpb8DH4AfidAs0sEbakqE2Xrh7N981babH1tDd5F8Wga8MqAXxR+T027c2I1W+R2+6BZv1AcQIBm
Y1RtyBV9fhu5gKowutY3iNKFFzzF3u92dAZ/OZUJmeWIFdPobKrrngJDiXbKcDnnl7cU1nd8fqbR
HmqtD6UZeK/osj4anucbwnXy/58jjypF+8vRJPBn6UygK4UESQSv58CQiSZWnpHIBruUc3X1u4/D
T5llc4l2tBpUwU4d/zljzN3f7xLcRqZI7lTnIbDcekKCbZEDlPbweK/7c3VwG//t/M20MkbJjYc7
MMQGl0D9/WMRfj61CSDMFdH9wkPTTErqYVizkD3/hpYnQRBhVVWoxnjN95cHpj7C1kNddQ/aHjWg
+umfORbDMbQy/BnKzjMmxjAWEY2XYPs4Ep+lKp6rkfokfc4DE+uBiEGubW1cn/Y+I1yjrDyLaRn1
owS3ghJkJc1ZXL93udMUGuvGStTLyIYwi9pdVIOa6iH6CrZSr1skC1Xd9+OE2eI17fOdnub4EAbg
eWK+w0lPxdi82FQ2mKGmmHbq3sLRTjJegHVTlRW0gU+Z3pGnvIayFg3RusqkT/y89wojRU1lfTRw
6iLYg//rLy2u4W100T9JzdGwmRtx+oEpaRMlC4/sfu4KBDUGCk+8V7xBwCwhqEOk4QzQ5xnru1IM
nvjscKCF4txrJrGtplT3MWXnHY65WjE5OQshgG7lwYqnBU4bxrfk4nXnbc6GTASN+aXOUSQE2wJa
NkioEM5s7j/hrsJF4+00KkDdDeQMtUtgjY50fCODqejIgbATbtBDdj1M5H5a7sP0GvDANYp91yyY
KtwvOojomYdN2dg5/YpNxfIPk3f/U9YU5ZY8RSpkgZTWLBHShmv+qinLa4nTrhBngirpOiuxSJ4S
kcqqsfs6FUIIy9B0+11jKSYD39GkAotEXyVyCn9+Yg3a3r8WYTIGz5hVXK63luB51ypk1ZDrX0GN
GDrnSv/D/pqLyAxq5tFxLi9TMjbO6+7ZZTq/Hr0oFSEDA+2yTX6unOG1Xz2fcsW3XtUL2sqZI8nQ
Qa1/IzAKFhtKKHNIePvLXGwazzEa65pmyRR0s+l17fzTBQnfk8fjz1K5P9yQ14vHtcbwLySUAK6A
vMxpaZKoFTz7ONJOeDEamp9gpdID4WPoel1Ep3YllAkI0g7F681kLFYxqt8jpOtO6lHLiiXh49QO
xVyodXdrVZE7IcMcGit+RkOzeRFnyMZvqjYOXSJSPxb1eUvH/QOWoNgkHTmkdtGm9AwXj9R0e6Ft
USsRBKdShfPSprfBCOtrEgEJENyDdFG8p9B647OLW/LUvEyXrmjf0dIeOGeuEeHmMeZRWAbXF+9z
FCHLXCxoaTDZuSlvXacDTcxfuFNkn7LwdiqY15vntGpsw+FmdxzK8EH4xrP0vUAfWMVYeZvaGBUR
RKn/hgmrCvGjwdmM8t36EasV2njOe11/dXxImnpL9aWFIpEO3/tFXpMxzGKCbcaC8OeCUmxr2AeM
WS+cCWIAfSv8JkBPgZu6LXsoTjvdJCnFCYJBMrUM7oeS/qPbOS/dTVsaw5oU0YanA3y7Q8PtrJpX
r93dFMZyYj41KpPYX5FBY1twkyeeAaVNFc1QZ5VQUWYTnUi0RmzQAY/e34LonFumtqFY/dGGjISP
EEivFGeP1+RoUvebItZTBAlKnLyCif6A7u21GDXIo1m0qjDUS86MdRWuJZP0PDKf4Dplp3HrwK4R
y3KH/cwD0XBQr32AJa22PhlqwEywD6WMcDUCQNpRtAXlXmcRKv2QbEnzMrvtjUktipG+k0LeWVIP
eTZuVR5gXhVZlEd53pYVIAxPXFcR8XrabtDSmTcdis+GO3SK/osYlE2+Z4yfC2jHLZdsHdOJZKPK
suLiAyx3fUlMGnAOdTGexOc3fiLN8zX3g3EtKhN8/52560MVc/1RCfwJBAxbp4tfDJ6IfxD6b7Yj
5MrfxZFn/OWb5dQkyhuJIsGnmXhZyD/vfJNWrz4p1RwKRRLBR2+qA0jHNX9P7CwT5Yyvr/RBGEQP
lWTcrKW0vKgjTRTXcLVQNrXGc6y4EHJShI7GsBuDQsbx7zF6+mKfbTyylVDOC60Xb9hrkq65BFwz
8CFokLXP/ibsZyCVEaD5jpVS99vrybEnOFJP8DXbQqhgq/GgMrbFePQQtoj9Suvy52+dck5KTJyT
7lPlfq6TPKsWYn9jY3MG3WHmnXVJtaKyofC3RjZ1t84VuarLbDDrp17BE+9r63rKyuATZOh5IqTY
FXmEWyRwVER3NSGjabIH5OHhnV4CO0ZJK3MWLZ/WR7e2TFY7bTblyyc1THUfqIFyUvX/oK1AiPw0
rG+bS8xfLhpMCwHssyrJ6lV2Bxk6SGEhua0rlWvQyG0X3ouE0/sW1azzkFXwe8Iju9KYbcFZWyYH
e+tlkVjGMM+s9DVq8cNTrN0VZzus94oIDLWBzNu8EOZCzA9E7J6GDitHHpIFya851/nlRBmNckbL
tB476oQnMs9+/btSsLgEsqtNSw49VvZ7lUdQjAz9pNla9h8lFMxZq/ejeKEPow4i1oyoBnJgHHy2
GI2pTNcsW6OEd4Bw2tB6ckMvXlKNo69v3FyNryU5bOKDX34xW7UuIqtP0ILMuaY5p67PU4KpZ9m9
ZMXM/xwGTYgPExwFkRvGlBFUvAkA1XwKS+rlgx7/t72TtD1OyNczxqi9VIRvZPfFduRzbgVDAGu3
l6IPZoLwr/qk5up6mnL2DjkKFPoEOMZJZrWx0j/nV2YDTRiDA68LyKwAFgNXH35mz8HHT2oThxXg
W88Sy2sMMX69TVc0b72RZwQvir4979+rQblwrx2FPZHia8b4ZTjrJSQk9F2sZIEE+GC8XvUldKPT
5Ca735Ifp/HG6EVf8pYJzbwcCBSLCaTWDzkum1jN4+7qRbiZ7eBWMU29RsDW1/Er2ZeF04rMsZuD
TaL1PSCcrttDcu9qeju3J8ns9lvvcebIhjRREBdF22hESbxoyEAPT73kyIJMvuKlICGrLbAl7DHD
IAKk6b+UCpHK08T15xWvXgGInnzY9Mf2owwzcc/TECICEv6vROWHJOZdO/K0Gdfh2ru6/3zlfCnd
cLG8xMncYJNB7F3fSyEPm22nn2Va4XU3JwJMMPEIi86q2WsaLQ39hU0XIOhkRvlJACITVekTYQzN
GpXIX0ZGuw17gUABMPP1dvQcddtoPwiOxBUFCKVKDe4ERd8CgiXZxnfrtDV1J4I4rq00cufgjrXf
4RY+Fe99UqkkhRfri3RtdhOYLI8T/UIu4vZ9lnGn/XflOwuXUUZeHVldri+oRB372BOyrend42aU
54oHydnr0AoNATXRcuCEALfZaTW2vYlTjizqigS+5m6LHuR7b2A2avwkLMNjbb9arKH6TWQ+0SCk
k8uo3WqKzPMNhzZHomim02AOUROMQuK9Glxt8ScF5k6hxhUnKnLtaKLy8mjBZUeL0FTibnk48TjE
oYMeMeafxkdsQe7XLxPvtOcBSZfuE5P11Hw/6F5Bn9eKVbzBI8RXvI3PnWPBZ5ruackCGNttWvLN
aFALUJZmmZ4T4zUPXVvGNAmosIlNNS9PF6Od2FrwE82Mrx4W23io/H3xrVIUlwxkE1s3MdNoFQ0k
sShQOIqITgZ+IyKF3ndw5YxSppYWbZyXl/ZATdBqojtDnTFCEXcI8c8EMWHLZkZ1xe7XFqC+IojK
RYLVDnYgKgqNFutHlSwvPREnPb3copk8roLpm+2vVsGjXKwg+GiRC4GquFkmNo3cnsGs+EQDPHnR
lmOX1F9DeLdKnp1igqemoSZDWkGbSUIuvwrEUu6v9Q96Fd2Xmp4tJdg3x7ajz6yC9c2iZLNolseK
tsoqzWcZYb687sCgzBatjQTOtikDXgrLwSY+yQgzlON5wLUEuMsYqbfW8O0t8DoUsuNe8QQui9C1
SloXvwZBJur+8V5BG1CxDxlqEZ1YVoT5PFlv+EWp/V5Ux/ibWUCKBLTtGYfDDjlyN+4ea8kie3Y/
dq5KIFn2af2Yawy3Zh5JMoezbSpZundKTOolm4BVR/U/MWdC+oI8OJOnoIEbeGeetpqRIN3/dxe/
yibsqNjG/5aRPywIx77iOxp9Ip/QN9S9q8sGwL47TR7AZVwZzCrzIx/GYMIOLz7oIoGfOfgQG9aC
3ZyDm+kij8/eZHitXWWCPCsyjpxKtdIX5iEegzKOdpmGvaFRPmgHterLb2eLR3TBMXft+UBgKWAu
utEOb2TGqF15ojBMgbQJdHOCEdm+n+mv0hqyYpkOsNz19+qJxbB82nlZdt3sMsx2qYln+4mUiWu6
Ny+SVBanr0nureEEqhBjiQPZMOVLBU1FYBECKsQLgBHxMvzOB9PD62NUNtwHdOo9J/pBN5qIxERa
LYfXYwGdrqeWT1XJr039ODcbdpMSTUCJ7Omd/RjVIPWzpT9g8HIghUvakbia9nya+M+ADoJAwEQr
5ulWSaFlGrBTIFcq7kEPR102pRxFYfu1H8YoCnwAeBWRH8BoALLHJhhx4qOIS5mw2RKULY8oka4K
w+fSwufTfKQpO+x0/PP7tt/SIL+5+L5cdWTqvp8ZNBtOuTWD49XZnvat9s0yGBBoAsUzaScxcFqn
/JuDUW7Zp7GZVllrJim5ty79I/O2aTojHE6qDR3KUVNs3nQxStH9UFGH2NFeMWvM3yKN+hHotQTF
CItV8UAB6guO8pdJ7fz70TWaKdxT/lwi/RPDJLB84z+nqAL8XAMkqTWaKT163ogVXJwWQgQ91sKD
1ZvOH2qMceWzBORWRUlfsib9WlcdbhxKqY3B7FZFdiR0/A/6CIAv270AHGkdE2h/baQScdR2aroT
mK5ULbF5Fz9YVZV2C0Z1/CWo5K00ZXj3dIsPHOM3a4i7Fvjkx5NAGQ/BVy7X7B2FifgHXdv2K5hk
t5TN/wsu9DBE/NePcg58KPsn6xcGMOQPa013m/95E8P8Q41F7uKZl3IfQp6JdT3N2Nq5eSWNbF7m
X8hhHOfkW1MEBaADk7eW9w9B/XOPwgx1pMzUbb9R4R+M42BItvhrvBuGWmiSFb1hkTmUSMYvtwG1
aqYtB7NWo6ZCJwups74B8CJbUcdl/cz2fouabTxHnEDmBWHHHpSTJ3oj6GRTg7gfGAdchJxE9N6s
6tVipY4I5fJPHY2j0tt093TN7Qlg6jM86UIA7CJsgRFDIRLIui3JuLDYNPQ+DRVgVYUKyaR7bMeb
XTiFJrYmkMjHIik35SgD3HBqY0QKCtukgDgT9SpLq87ByZbg8XjuNP7Eig8M3UgeTeyz4gJVvdL8
b+r29AXydiRyUByB9x7CqE8muvxBo8ah3qQGMINH87o2G5JzcOX+SPhll4mTKPLuc3A7/dXjJrqA
emU4/x2BfZIDZiGnRhh3vWydrJ0xACh+ZiPUop1M2mSjxRXv0Bgl4Cb7z8IqlEnLBHqewYc1vWBV
RQH1S3u1Ema4xpbWZasxzueB9c0RBiPZe2bkAjrn8VZmJanPM3rS8GZbytw8hDj3XmokIbekZJm5
dwMIBLLbbQjaUuNBj/ptT+xKIJL2ibqUKmeo26ONgIo1TeknpFPu3aKGcWXSb9Ee7GYdGey93T2/
poY1bpSJZVlElzEyCK9HxhIxWvbuzU70xgYUVb4nKRC0m+l3Nl7cYaAfLmcZaWZlW/rsBrHalHjF
UWi2HNmvRp3Sn2W9L0qSeZazFgfPxw0BZ5bKjEr4w8CRvvn5h1BwpXloC+uf5eSFYiWRkHbSCpiZ
QyDMXuXlPIejvug96ibdnEehcuE99ijyJp+Ue1BSwOoZy2XXdkl6vD3aGBkX0y6mCM80y+eoM7E+
lP/JcutmWGxT6hdgPxT1QoJo1NNSq0ra5a0bnOEMlnBfZSPK6xoFvq7/5mmJvHvx8kLx7cLBwRFk
bSEvv15N8vdvwiXh5XNM7Kf+verVy1rGkvqZtYY29ITUbji6+/uqMMwlIU+yxN6FXA+55EXPDjBl
/UwIBj8QXKU2OuU0uFPrMHBJz9okOwOenQx1lWiOufLn22bLVx3VoCvUUFCgfSRu8FlFo9Wy7LBT
mSoeYHW8oWH+YZ43J4YG25fpXdkha90bo863JPwi5rbOFo80VPmiq5WU2aZKFpKEpy8jSAmJUOe/
b2H8DxakqfWsYjlB2rriK2KVEID19TROJEEq4bvo+cGqIcohX1sWZqHjkNUgNQolgtTbL1DyAkyN
hFB6LxyvGPz98CFT8Nn11Vmk1So3fUmhKU/LOLNazKX2Stpxd087g5WL3Fx0ZWuPLxkwiUb0OCFB
oe/abVz976qGXMPYgBJjDrSY+B2L7ks0J5AjRzjEl26SSGTuPgo46dpYRth/9RcVcu4Lia5rEXIb
3uBeqLQcOJV5uOOqQTA1hCY8Dlps/pMMYoZH0IceapEVCg9nr7v93w4DqYc8mCtKyHcdKyscUB4F
6LXwVgI5nlDoH6b/o8R3GOUTUSlW8Rir6a9uq3+rEZkwR0IWYqPBPOrHhV+WemjxRkqvoFATQhYK
RtWgIcje6dfm7iIW9aSSltJyvr9Hjo8IWUUAjosXLpxA+qJu+9CyPq3LZLZ/davW/ySyl7Uy+XUL
/gGkfoCzK/oNmjQ6lH96ULkJKN9JACOQRWPh9sUVhXCxh0KVYWHGh8XMJYcSuA0pn1DCVLAiNfix
ZG2xWe8QSeuYe/KRa3XsnUkx3sLvGhollmY2fMIQ6LSL67dWDHPoKer2y2QSWIfNhUMqgh4rV0NW
TmAFOFwcHNAKe3Bwjlmu2hpYxIw/2f2DVY3fvXrumkAGZQldDb6hwINMUs7GzvsuNXxcJ6ANeEVf
c22jDoFSCeXrfLJt6MLmCsDxNdaRZuxoJa9wOL2p4L6SrXHKEMVx1Istisj8A2WwB1LCrosdN7YN
LvcZ2ZajvdY7hhXU4gVAG1SurSZ27NTyD0J551kQGGDRcgyKJXHakT6HVD6QMe8N0uX2Ukki8BDv
HmD6NALxGKEGWyGbTvbDehjT0KSflO3zgWssMHr1xN+QHasqxiv2V3eZgVGzhug0mR8fbwpCmznr
bUWIHKorCsmJ4aHDAp5YRqGUWkzgyiUNg6OB5RAGKIA1dxa6bi7qycCuuZ840GfAyhotBupR0l61
/1ptjdCdvEC1FRIMCf/Z/enHiPULdL3wGYnmOr+j91thLQl04Kvjdx+pm4uhDAI6HiVKKB6ETpj+
+AsPLvUj6M/fPq2mRdvgewHUW1VkThje7LXZGa5AC6QOhTViAHA6VnnruTnaPKtrDyv82e+qHXWb
TXuWq9hVY5JHiYHioqBW5V3Spv/tcz1nazu5YLfIDa0HJ5wp5iw6ZdniL2GLfAd4kW4xQ7ebJRJi
PiA8iusAI50pSbm5+AciftkULKJYV/27yu0nHGRyRZu3C2jpGBlcNpCdpvFGPR2B4De8YTOq4Zjn
Ja3QykyDHCu2HwoREdH28XHfv9LZqbeRqHNHBXBPWnB3uINgoc6kb86NA93uQcyh86/SyF6tGNh6
TURr+jtekMQgcU0knug06F1c/8y2L/RzJsN8PbQ6gMIJAf1IkQRlJRQi8fwgp3VMoFrDGbI7JB++
KSPL3dlUM4hQgUvnfmP4ph9ootdgBHu+dnVdmx22ZZhYij4G0ZG0nVdhUkJN4kVKY1qjAXvlNDGN
z0XMHS7vOM5pjFNujYIUyOdG7R+O5jr7xsdWDFMWeNcyKmNp13ffokB132Hh0Kdux8HP/Sj+vDqJ
geot28MCa31TNPogUQIE1b9xGDxZ0pSgWlAELjSZ3pxBlics7h73dFeEcMcbT4zCUcjfWsak/yA5
jmHK5yCMMArfUJHNtewZWYrofYFj+53dTuT3CEy1ONIvryYfMOO4vViidCBEo0i5pDxApHCXEUyv
2/nyPfVDiEa2pYhde76wIYASgZUH5qPMTyCdtB53Ve7W+RUvsU/xuZ+zV2E8LMIHUNsnSSf/1fml
niKT0x/c9ArnfqhZYaqw20goFdtfHBcvAqYGJKeF7I83QMJvh51kozE0HN1+2WuZKco3hrTViK/f
22rh4OUrD25vlbOWqOJ/JlNe3NUYhu1JspGuGN8BI8wODF7N9sDUa/vYy95ziC49KW50Xn8EVAzZ
YNeLMnRSWObYlImSl520DH7yfv+phXNodCEnBy74uVZUEk58KDg+FdSr/9BXccha5JY5BBP+UNvH
ntt3Vnn3TFs/LDaMLqwRJl4cla0GZTXN1PlBOFxPGjOm24Ih9+Wyx7vo19ku8FfVveBawERDR3kw
ucNuHgw9aILWJ8IL4LKFod6El8Eb4nJK4LrhXQPfu8MrgbJX055LMShjsQ0ft5YqGRWDNwQxGfpA
t8eKnzFZTmVAo0TQEk9gKTaP51mSnkIfyYqthHtCHQFXUEDtVSqX6IAFoYh+JeNUMpp8Mv5apwQg
xxevbg6Xrl10O/PbBqgPzZU1Cpv2h1nYlTfa+BezkGSmE4Jwe3dsJoZKeqfPUTY7InlbbUbdKrhz
CCi+CefJuIzx1D8kK1jkubMlFVxV2rZoPZosRSGOReFhLwcJ7qA0gMLSHCVTRIvfUMUVoa9O6HKL
snqSxXZkSdKwdvgiXq5RWnAGO3u+Qfq2axuQ38FDqxrh16JAhM8Lz5ElFgEN1UIxU7eiP3i296u1
/LmGqzV4hN1BbvkSvSQYM8pcpaQWuyN8QtDq8EmbGE6SysRqLQ7bYhZiCVlvcFsX+SvkW73nH8/y
9azRqpHMbwP1B2+hfOUv1aTv5/7GsSa3po3EkymRib3BkIxbAyo0hRiOs/9PjE/9XcXHVS4DhCKr
HeMRcrian6GbgSa2S4H6N+4YERWou6DlNmd63t1103slBqiFiJDbYPuHoKJCeiNz9y+Jy0jRYjDw
HI3LvjOilO4WiJegVa6Eut4tOxcdHMfRizVXR4/jH8LYRgPm+1uIkLh3Sh8UTDS/7V1FAj0mmbvh
kxWjHcL/vmFO1kjJsFxh6wJfRQd9IbQR8aoc+Mn9GX+sE6Dz27dpHws73JNQSq4Q8sX9AMCdv+69
GRBH2UPmX6uAO1Cdwg7YY/0ew6JT+fp2Tsc6BlbPk+FQVCs402DDAFVYtR1e2uyFRvqqUJEbXSui
qKdsSeowC+dq+eL6P11EXLeDrBL2UVZoIO+EL267pr1SPqWLedc7XcVl8b4FFAuZ7ULaCq1HIq/F
6l9/t2gMP0sJnGwtfFNSj1RsDDv5o8Rt9N/qaokKaf+O815d/zvPo0BBHiA6PgmTPl+I9JsH/Hdw
1rwl3J+jxn324Wk6nYSkMQtncAZO7Q7k17+vpfvIW9osFWi8Z+V1XB8XkUwIsx8BE82J/REP2Tqt
lpCfTr6O1imLVdF/19q+o+HlhBgkmLqx/6tjAaXvnRlzU+sNyA/MFL+uUdsOJm1ICE8USzW0/GSp
mVjxZhQbtIDo/Xe5et6sYZwhhLATwIKVWQtADBKIEPwDcldnJc+SdtJgFwFCfsScbAVW3NgxMuO2
LybN2VTrdgLzjqTt/B3JOlvn2Kg4uLi6lY0fHlwT+40+SXRF3w3SY2gbYyPC6xAXiJiKnxfXzq7O
b0ORS2mDuPM3+M0Xvd6QiXG3dBLZ40JI8JCHr6bwM+XtkHE3tG70kPIbTOssXmMQ0+vl1ikDcNh4
SmugAIj4zUUUF314KJTgbB7sqOP6OF7pi2mUzOO8AG6r9cJFqhjT3t9BUJyJwN50wEqbhIYi5Scd
nmkgl/dDegPUl8pXlv4yXdLb0ZbEgvhiXw4C/ZDaJt8uTeqSUGxPUU5/lq21zM9ibMgSlzA9uacN
Gyk7KVNcqALlnH/N023NCM2HgQlIc7n0mm3k87RxcBzEXOk8iXbjsZRCCeIShPjBj/tSI4FrYBjW
3KLOVMYpVL6k3m1qo5DFIwl1WQrPFkiMayvunLI/L8wK+wEjadvGi4H452xqxn6UcI+/bJ76wJ+4
jAfQQR4uMiuC9YS/ZgOi7mhQT6RTjxbVjgqtzbtk5+Ml1HYS6LgSijw+SuSQs6MKK8KjGr64UX8C
fVoV3FYSLN3EPYGnOMrkxQsQV+cSXAEDAmAbn5l2hNVQWkQeW8PcYR7J9gllHXrWrmmdVeK4a13o
PWSW4+MO4YtNtQ/Di+rq33jaCvGyz/xxOtlrAuYEOMh7ct5Ix9AcTzNzeXaUum4X+jXtXzH2XEFA
rftEVwSe3R9UhU0ZqjIAVDie+Paq5DzT8ZSSgoLmdYzj3VMDH0MWplee92KNNkwgaz04uUQdGQ/X
zKdlAJHelOoNb5SrWG0YT8RbNXeN+nkLf5iCPL81AD8agHE1zLEw+UEyEAk4ys2vlYqhQkkWYGME
FIRUkr7Vcv93mjrGOr+luYdVESVdxApAsyFsPkBzZY0+6cJrJTWZwJp7WPyNCoOe7ddtR/46voQs
sde9K/vw9PxWu74bTZrjUXcvvKR64ywG1N+FBH/gztTmbjzsw6CWS0KsbqJmqOFoGgtQ1GObM8Zo
BhjIlfhH3WifHZo5PmuGVBnW7SQeQlE3snbvblbbrwORfzeYDzP2K+B8vV4Y8sVjW/bQ/tDGOqRE
1WQnNkGTRaz2DNiT4r67sxECITS/77QPV2gfhx7c+TDGs5YaO94TxCrT4iGy3nKDR7undlQrIwgX
oMh0b1SWWHr7qFAmpIICPQdV4c794zIsd1CXhKFd63ASqJx2GoehQfrE077zz3uAZRE6WSilM3ZC
AFeKeIy0OO3ztOnfs4HJfSLiYa2wVeIYfwx64KkX2pexn5q11ODtgEqio9Z3Amc9a95ki4xZHHYG
3h7ZzzLRLjVV1a7DAhjksCQZHkNs7hGaNrsS5gmjQXIYGepXrqoBm2GyBe1hoOx+IPTTSw+whWp7
rMLAxtQI5WlbD12aOhMSbUah3es5udigFpvUli2NTqReXRBYgSA4J/rcKI3zsn6zyayqeiPyiZg5
jckAStYWtpOY41bXTk4/nvEC+GTtlVJqDb52x63ui8Atbd9JmMBThvR8Ic1d/jrKTC37jkaBU9pE
8SNNb2chnId0o68AxR0rLWtqWCK1enIzPepcUdaz26zoqEmhjMJi8SHIqTBewJ4ZLn+WeYhW2FHj
zdCZkROyRETjly3hBAYGevQRF+xJtd4lgkRAfLd7rfxOaZ5PF1/DurU+8a0saelDpC3NubWwC6E8
4tP+lzBEQWhRMaOVXpov/4RRMbaIS5qPJIsu1szGxB64VH+F9pN7FXZv1MeDBQ+KPRPmZ+siyE40
/AX9wmXEiyOAd//nX52cCMp9sunnPid+s9pDYD2MA7Z7HLGkp52bUHhDOcHBNZ5jT0nfAYT4mh4c
jqinF+59v2fzOeZYIHiY2mzDK9Pxp4xP0WjmghBCGJwuSEAOBb5UYRp/zTZuuFbmzBa39bBrRbDl
Zg/yFALtmoct6/I04HR2gBucz9gIKmZPBLpMgJ7sReVoSf3nW7IiqXoaxRnJeZRwFIhK0ntR8e0b
ptQ0h1v4+ANt5VDplVzOzdWypsIohL7u5BsKzSLl9xaQCjrLO9Roe0GZFQbQal0ew0rGHpXcRcf1
wk+deagWEs3wCSG8SrTvfje6ly4sCLr1A48g22nlmvhGnCdFAIxyQ6KdNQYtuUVuRhuBGFU3G9DJ
arZg0+YWzhxtGKeaKNipAdO0Rae3XfljkBx31sbwQdYYEYMrG7BpTm/NRhI7hKumX4IG6ZI8isXw
ZTbAvRKwck4KSW+R14TFUrTKxyRBKnW27M8zsYMh5R3wIzL5wJIYGS7YEEcohyXc+xHWaAjK3G1p
GUNb2+PHWie4pFzz2VMsoF3WJm/gEPCfUFf1I8XsrYXKO9UKLqe7zBbvPF3J2VXqReX8aVeApUf7
fEwK+8/Dml/0gdnLGUMkfhqV6xW5Q4N0g2SMYxGjSQcOXGzoustRiBMerABte8V5KM+iYjlLXZDC
7f0juRMqH33WfSGv3fWXytg+dcIZeaPlneHVridxFHfDwTGBYzJOjJ9613co7z2Dfk/yWYEpQLoH
Vd25eAxk3kPU67BLCMOhnIxObokCGYA59G33LfCRvDWz3dgxskpjnGC9Z9x4kETThxkNuO2fzssJ
XyZ+f8JZHFik5ZZZTM0GdeptGmbxx3EnBx4YxHTBNWhjWwQR1dc+miTbCA0kPcnVDY+4b4poxiZZ
cz7GfMvYgFfy/dDbGIJKXurC9lQGmcpMNk+Mtq9869mI/xh/vmzlPieithoHfEp+iLZF0aTfQXnK
M2wa6x8UPucxLMAV7uq8rj2IuojAJKamWMCaEDC3ypyhTDFhNBX948uIWG134VenJiqzRWwIag/P
F9OKj0/3+BLXYU8DIA0mkeas5KGxfGW1ZMb8w44hn69vjXkjupWQG1cMhuDSPyg/1howxf9dppKE
EsX8t5XygdU8TOv8MEb03IQHLtE8NApkyh6a8mxCm020xqdlyVy12+Zupo7PksqwjB//0i8/SWYN
svWYAzDxlGxAjMEEwspcskWyTuApTStxa3gKBGXzS15TovxyZPNzmV/mqPSBzU6fVEUvaT7eNASL
F4u9+IAFe7TIm6V4M1a6dK2nXSKbCjk1pp7utaE0A6Equ5apefvRu7psvJoxjI6tHBXyEKn7VzMy
3y94r/lwbupWEkn85EottosUCcaNZcdZDJy8RXbCKkh8+V3Lirk1aVWbVFBl/7uaPB1TjOF933/u
jBYeDoHNDy3YQ0MBCJNRKXr/bK3p/annsTwqIbignZ9HX9Y++vD31WE02sPSU+i8pZzL3d4KPA6k
uFHl9NRfdY3UfMa9ErT0MbYSGXBScnNmnFb7FGAdzcpjmho4p7U15oQ2bFC3vMhDVXnSI+K3m+Og
qDiTekMkxXUeryc7BaxWDDLYzc9xutLrEqnMzh3lUtlyTxYCqg9ex8XPZXsA+q2LFOjsat2pyuXy
Dl/7jLWaiXa6xWJHLTkOgW9wI1+mCRbTjFHGby0+/hDhJTNs5H4sKsZC37MwE3nLlFa4SraJO0Qz
bJkCmESesyKaiaeUKrkv7oWIEPa1dXcZDYVo89/V9j1IjR2vPCM2lAX2PbiKs491bt3t16i2YWtO
IhJiYLQynKGv9HkUrboKeCEUw6JoSgQ5dnQQVBra4DBRyO/bEfh52S9Dz+Yzk3nvd25MaD8A158B
eoDRUr+jYWn908qWSAU0Oh9/aVAVbMLzsQgZ5D4r09X5IPu3M/iA/IvVWowzL6P8+iUswGylmMoE
joD7kedP8ORwhiN4yA/HVn0madlJiP+Zdd7yEj7+XPIfxwRO/E0RudVbd9mNndDcONzJFhCcCmNP
P9RQKioSqTN9oHk7EDhhyIx5BFXUpzlHMqwn42Zt+KuC4djyg6HOu/DfleiW0rn2wZOobU0SDoW2
Mw3DQ9PIC4FZp6WMgaMMPNaR6WRmyEOPpks6Kx1DiiIYub3NijDw+p9VtyrkIt0gfNFgItk7CnRp
2jndl0gwc9iIwUEmNRpciQnFXOyfjpsjV7JZaTOdjFIX2YLIJtrXL8DlH50OZ+5iJuuMM47vjGfe
Q2c/zZeJadifqJfxbESi0kLEQghdXoCtbdIB/l/QYNw6G7cqyY0VmazlCgk61ebChpEboV/ssWPl
OTgPvqPMkI1NrA2V7qPTy9QEMfKuGL9XjAmGcEaOy3nGyVUtJtKAwkr9g7LRk37f/2x1kG+renwi
8UlkJS77EwoaOpyS5YOuha/TI5td0iewCpSfZOIV3DiAbxRTLPsh7EuL9MMFiLyd49oI7YE0sfN9
JxGt1OlCusY9qGg8vLeNsiOhytRrTlNBH8K2azYulMxZ3zwBW5gD5W2FGwJ9xCzMgWx7wpr22Rhz
N1MtvZYE5kjfpZzH/7IgT3h920fns7FSK+p/V/DuyQlpEshrI3lG+qh9MTXm3EgEcPF0aE/SZd8c
J2IwkF4vX3naSQclSu3SGYuL/lxs1JzFdBP1eMS8EzyoVGFdViJg+6w2sA2OOMx0gALDVfzpDq/w
G8ip/51eJOZ8rQU8IUlXvcO9Uh0W9ot6YJP9Leo6AgOvZBBwgjljjALc4bmXArsYAJfXxoYQWe+s
0YlaAJJpySk76l2CLeAoOlC9MspPqC69dIHEb5KRwLfPpDwyrdr2hs6G1bz1Fdr5nMJ+YKFK+B98
UlLZjOZE98xlnXAJ3OaivUThfeSYJZUAeB2fzBPQZ8n7L/BeEjKPqP8NWwG/k9YD/u1z1cyUv41b
//ug60vpaYeYUlEVCA5wCJn2y947+WM3K2wpVqEc8ZPr6J5MiNkEHipCKdk842M/l4niYDsHTHon
qPE93HmNCcuYqptUi1C/fY5QNQVmiKc4AeSTH53eb73WOp4WlrmPj4Sa09dYM7zFGA/o2zt1lWSI
bsZEhdNPaODtWt0KWEcplgT+QaV+RJd7WrWjDwSR+D7e1vmRCVhEZ8LIjYwiKoiXPZRREUpUxZuB
S/XbJTQzhfax1C8GuWmINYa5tX/d0jIHs5rkOQRnm4u6QezJoOkrtqHTecwvCRmqI/Kbu4f/uj7i
ql0papGx2+vw7om1r+6UgjCfKhe+LbO7HKyGMld4pV1UN6cUgRrMp1cpNz6eaAdl8qnnYeTgwgCa
DZADyrGOQqldwukzupUe/BhTf+A+R0A7RO5GgbEfWn50k8TO+sYNZ5RdBADJ8Z5oX1kouy0MBch1
l7ahit/O8122XhQCSqRPJf9q/YpmVY73t3nCY+YelWuPjEsLX5IItpuprgvG1GXJaaXU7Au7B72/
HUSlNm3NOguXvdGnWZd4e8z3Sy4J482eb/7tuI6wKJfTUqdgtcKRrQvtCtyK1TByQGMS8qmVj261
2tiV1pfOFd/NL7SJY7Yc+zG0zMi0Z/BzxkSDMd0WcW0XkmSskZe23+4tkPswpNvjs+DQuFXsAYee
0fcDvm8+bVwYCXUWLcSPu+DuOG3vIgB+Elycwn4cP8axiDe148k9s3V2pQMlHLjfRIezW7uZ5gRM
BdxdPPJkL5qY88UyApTxHSKBgaZP0tlDSdIAgefwYSpMZZMbW0CytIR81kqgNWm/3ma0ISLbr92h
tPGRStWVwi7F3CqrJE6fFZ8NCNBt1KptpRwFRwJvPsu1WOA4B8ejSmp3hXEtCrUYNNZBidE079GR
DBzxPgjLUp6zxvkzDeg5ku8pCaGaEEos34GhUujO3oFqkbSfGPy3Tq6nP2j0+Q57Vo4vTIlBbQcC
DfXY0eVN+02IfMX58PBo1M67xmh4MH0HtLVKRX6lTURkyGcH8vOX3a1AEMk8ozDGzyyi8Dm2Kct+
dCpfOk9rIMkUmU/HTQBKxFu6WaENPf1/tz5W1NWJ0Htzo2XM0zAsopLX+Yw+sEWq+X9wm7l24od1
GccZYYTaNpMwcQyHvWzoj6c2T5L0Ao3wMW3lTXkqZ0ULLqV3TgvbNTIVtMHXR7wa3FqM9p1/3xub
fHO+CModolWuOCgWclZCWXr4D0N0wfBuvK6ykw3X69vu40mnLe15F7Lmyqy2SlomCu7LxurI/OfV
XKbaC9Jd0H2Y4AnQjqyeqVGj7/++PWVwVW7brwb5f1Dw94CI0kzrZcJpI2Teo6k0mOUVqwo2cHQS
WkJm90vmr+oCPDTBJBLLe/1DOsUOnRNYyf3psJmOUCMRxSb60vwQx5ox0MhRNvFINazbkgvrLPCY
pcx/X6ReeKl8jgrLWdutKOFSYN/loWA4b6W8p/bcEXv/1o/oImkp6nm/lJIlAvq/cwHPy78tCSyJ
0tWeliqZB541azRzPe2imJMg8eS/UxBcrvuxbykeO/ywmkllm8oLNkS/Ma8e6j0bzDqAo282nup0
ZJwg7Yj3HuGzR8QtKEwVD6sKUSS0JDJWFxUMozonFZSurSDY8aQjnx5UFkJjfosKehj4NxTStWvB
gZ1fnvHWIwR3AnbUXEYfaafTU4yGfzddBVrXBrpiF6LOjLwZFE0rw/hhi7vOJgjf3JVgCw0td1rz
nMPdSTP7fsxOSV5zHt48pco8PAOkR0Z34P3VK56txozfCxq1sZ2T3oNhCy+wxI+p2A9YHi46cUoo
vrk0mx9LJgxgNEw++cdSNGYXDRS07TmY6iic72jWCmiUnR5aSO/0FkEXGT/iQVKOQBXW1l/2hcJh
YyPRptO3XkZ5LHfE/AmocMtWX5wiAHnTZMI89WqzUAt9aGJUIaEtAlsPUs3HKlehl9J5rliqWWOP
Lm4UxBzutRla/1H5LPbYi8grigLO8dQjx5eH8d+LSkSVI+dd8vHEGPGxuLNN54EmcB0UnUF/jc3C
qYSwekxepeZ4b+maPVFPQGdRrbL4VzHP7+96RedB3LxT+U3ZSu2WmLxHR565fIYw6RHVi+6cv6gI
vUJ1S8bCpzEL9xWz6EcVaoSgh1Nx2myfVD0hFEMrmwJro17MgogTkEw5j7V88E4uZJ6Yi7IOQ8JG
nFPUObTEeVCz0WapM+VVQSwXwREARqPeEnbjDasc1KrQ5vBfsc6GZRMIY822Tk6AHpfXuGv0bN9a
ylDlw1eu06zss/Bxn0u0nk8x0Gca2M3GGFn7hSf5PVwYg8TfsomZ+N+b+oh3LncjLMvFerKm7D6y
dUdT7pOAiLJ5h8VFYTe6PBZfebBu54lqgUm6VaFGWIPfGKAAZK2iKeRV3ZJ7muH4K4JeZzODskSq
IklKUMH+YyFciMxyICrXEba74KI2cs6kRA8easK/ztO2dclWCo1vYiLIuJywzPdCdyAwFDiGMwaN
lARmYn/oGIU5V/ny5NufSxE8mvRs8SNYLEr5lI9sEqYR/7ToRSJRYJVeuJqT5JCJBIBlHXUs5Tni
A8cWWg2f2r6qnnoYNWMPITDr9WFAcP5YgagRXpEOib2QcgRy04wY52yXfN8/vtsAqNCJF8sYZsn/
XajVpA6sKvpi2g3S8VKj35NxO+EwFX3BwKyvlMtsnkLpN5UDcmYhAh12irtamdNtO8EnnesWitPf
VSij4EwO9zdhaSHg4VR60YL0va0/g2wMw4Q8Q+xVC4Lfo23XFVi1rGyx0ORYDW3rDTpXU8EyqPBR
LHJI4c6Q4zbaEdLuJ7YiNtpZb++r411zS1gK4i0Lmw5kTVEWTcVxJ/uYwEZhpzaPN5b/zTrr15/c
EnTUKEusuZenhYTW0U0LDZRa1aoH94bUiO6UcTEwrotMW1zUhgl+YE8rWg0Cj8uo3UN/B6kc1pJv
BSRoa6Lv8xDxfQIv1SSnp5tM29W/U7kxfXNDajTo8Hc561To6aB+/ausUzZtYK1nGEQcY7SCTUOp
rAKATy/eLBKrWbx9rVfCQdex3J04ibixTxIHaU+zh2Q8wDCrQB6Rx1ze8Gt0tmoxdeIwkXjoNrHx
yfPc2Y6kOAJBZLmbMyFgz2I+D4XqtGq3CE30KKEAZVHZg93/QiNWr12xiK5DXrS5M+rm7BwicjVS
nk4bIvSTaL9BGEvre2sAttu0L86JqWEU1EK1IUZ+G8ky+cTc7zM4i/ChCYyj9rSd8e3claEXz6aU
D70wi5OvzUNlxWwqlIkoRPSt8hGnBe3rHvJccF67kzx2EQMqwSpgt5US2HB0Cbw1X9ugl0jG6CFM
cPsdusrnjSdDhL+O2qcKMAmijpeGBtEMFLeSw0iAiF1VZHhofsAAUOjH3RfZqxCCG7DREBsPjJ8c
ubXvFFX5LGkapXfEjazLK6ajiwCY8tfArnU6BXXMe43B/JT6BMAg5KOXsYMkptfq28kejeQUtuP9
fFbCVsI0IMMJWTHbIF3OM/aSdZlX77Iobz8+b18K+HoOMy1Qsa7lsd80/mLNqYdBS21nAlEm5qWJ
I70KwngQU7FY5uL+oEF/tJRlReVSDmnEpzbLH/2k/jiic+DHEFMN72EzpT40ycClaeQt6dMaTmBv
B6efbErEQoWNTpb2Xqx4e9o2fuCDp5ypD/1Yb3aIFMVXNtjOzvQ1hJWf3e+2B/iRJ3pQ8UaVj8Us
YPr0xLBi4gmnEwJBayFxUAuhgCMPCt7Zud303upVkaZyG6t8kv0aQLCLLyQLgex7NEAFZXefhs5r
vvvopBGls84FM1mp9vqkfq0wPK6nFtp1akzqLv6wjZDIHX9NQYHWtZR4+5Sb3ItxsC4NO8PiPdAu
1yVTeEQqvj9vXqUISkAM51k+QmzDlyEfQyMsWLeeCWRQJzztK6mGoYm0eFPnGDeYFmZoj2toLDhs
LcD240/vHaXZyK1DeAdD+nk5cLJn0cZQdGHuQaYo6W1GspmAA3YFHBTq746how6k7wg6r/Y6Cr8x
S0Tyrms/hD4Ko5M40nzhZM4KatHF2LtpgihMdS0sx4HQk54O0hHN25fuYFeLPkPOwdkNOi0IVjXN
OK0A5hSUfk8pV44hL/eJ1elvAI1af2D13edu51gi2swYU7ZmkSbgOe8K2oL8Gy9gTKFsiD2Ar0/Z
BHNe6G/Kbt48U6jOuG8Qt/0TNWyGz/kalxzoy6FIbPqCac+muN3zZcfZKN7metOyX6ZaxPm3HiVh
3xuwjuxD9RNnqZrUwNPKRTIyvFjAAUgP2NCJIubsRv2BRRWj0Dw1NnHdVSBwKIQLmSk6oJNeIKc/
lYp5+ZtF3PPc3UWu47qLt9JUJRMCZDchPhrOzI/riGHSHXP6wPI/YbZ+DaeSDl1m0+0zzcfiem7L
UEOf+XnUr4Ld5B/aQB1+t6edFJ7MAvUDEB1ULfGLnwioLNC8I7AP4H+5Pi7hCOHoA8h2V0Q6BuaE
meRMT3w/Eu46lxGHqTRBi7kslObN1rieedKHeTtPb1BxzdByXRiYoDILXJlJROjukWFEuaRW7Fkh
xEILtCC4pJnhbn06BuvBtYwxAI+0g0DORV1ic67Eg5GIc9Gcc6BRgzVt5qOhzJtRO3rgJziYhvCu
sGfbhKtXwXrRceDbXm0j1XF5KBIlJOilJxrsePy3KInyqF/vayKwGq3bdrKjNMdYLSz9ZMWjoqvq
qhOkHfG5zwRDynifUuagaNOuH/GL3SI7R05IjyeQYVtJTgy8WylR9lYiO8I72GP1vD0Ctgu/ptdf
aJ+Yf7hk8eV1l7s5EbD9UbbiQeVSqDhRSHaTyFcHVbAwinkHwUcPkqTbfEXNI9qKE3Unj6jL5pmA
GtuncU5nck0Cbo+vtPaLgIU4qQI0hGn8l09e7+V41yQjbxu1MbF1G6Odt3NVnj+lwdeE/p0gbuSQ
ekKlr7ulcroi59TqJkdF2ABsnTGDxcId+f3lAhM2DCZC9CEHFigm9pNaxslsh5I5Zt4G31K8DOgL
PCXGuzW+HTq1dxKgaNhQViJ64aSYqTpTdUW+KJDaHzisUtvQjpmgv3Izz8GC69IjxHezCZgwpU7Z
gyKAHFJvEUGg1mXlBW9eTs28m8/AGJfAqzB/r5oK9t/dFVVuXo2E97AA0tzJKm2Odylg9YfV6fh6
yrl+8X8d7ESCo5mKzTPuizttiNIvSc1d//pmf27szrbmtmswJ1XIKgTG0bloX8hcMcTRLj1dNlq5
Bo3zzK1JxHNOnsI2A76aUEmlkqqIGoa3aLGl9lLz09kgkc2Xql6cVX68qh0ylMTjRSgLfGWxtR4Z
7uiBYlc7GkQ/dIcMvHIzVv4ncpB5zCwAIZuLk9QGHLLVtMkPr8dyk/PcuPCu1VMAitKgtSpwz4lp
/ZO2yeWmb3035U9QQnx37lZ0QVf5cBzJCxVr2F8BRcfQudpviTEhQxRgmEexgfQKd87hZdPhYy8C
q+JBH91vB1ePjsfFWSH1w0EKo3kh1USXRQOVXzni3nxQPCnsknIo8z/4cJ8dx3rFWUQMQSLnmg+3
BnfQGCumXjkAGNJLFwPKktC5oJRXxNuBWkVAY0BKL2lboPKOk/6LH2u8jO+lOy1HhlaN09eTpy8f
J4T9vNDLIe/A3GwTlgIGreO86HrpcReBRZ5Gq94Of5DuwDqX84et1TwLNPywBBNJJjO1yB25bL3Y
lbPuWIFOWzZ6Cr6SSWqEo5tGvbYly75AbiD2E5D8+SJeYE6DUZMP+z9OxKfqcDB3VHtvFAdvF61l
hx5055ZUojC4igzisXDz1F+KFu78uvykAadIuZ3jBgn2/gNykEW+PQgKf1+snWlpvbBN0UzbGwE5
YPaQYI59jgdvUQKeFfaC3JuG6KEAkTDTxqRPPBQtFqhIWQc7k6g88K3nkbIIxvW1cgNaWbdRwjF0
Njb7mtAWQKuwDDYfFF0WvPNQ3n8QOgi9mApTeuu+FpYRNoUKiWJrxpKMe6bzXny1MoiMi7DECa/K
KGTBgiKIpyp7g1nfrWBnLg0p90gIyrItR4AniXjGBsJrE+iVbO5/bAvunG4eGC0Fn7hG1U752UMN
WSdab6hXvB9FLbhBZJWFLGU65yX9VBpLjJCavF/ZfH1lE0NPNqwTc/bwMC7TIjKpH0QnOnLRygTk
LJ1hJcBvrNFmrgYATvKuZyEy/LrCIykgG3jnUCyZsY6WS3fbl4ovTSg3ZaR09+eHieKEA9B2gd9p
anxbT5OZaUU7C5QVZDhS4r+HkZEt3JL3BnhZ6SqBZEXNzejJSA/4tKppKWo19067vSfnK9rmzC31
B08gm7naeI1iK0EJiSeXWM/XF4v3htIe+A7hQuaIVDA+0Aiq6wJQt855KcWfhIdZ/F2IBrpxPqLN
k9zN1pc5YzwGB2JSGbyLf7dp9y6vqaj/42SAMNvhlbszJBs+Hv8gOuHNoiAX6tDmGTgLbdOkbbT+
Uh9FLkEpE8JN2wwdaBDGTRJlWx5wAz8Re7GBxMcJjdfyizhxhgtDI87bEXSSSUCbmhM8j4AVpV6M
rF4IgInx5tl+hM9DuVRKc1PL+wZxg3W1f/DyLXabVrFL2WdWCuAfNuIIsxw7yBctLtj05p157F3R
5Oc+ea9K1o3HImA0Lp1BtXNJWdbLjCGSTlxrU/pAHgthwG6hcqeygHuZL3S6kH68Vgf8/u5JEdnt
oa7bVUvxyqx1IhqtkQ4ujGLxHvrt5ughsw7O9mQROT6U6TIezh+1FxKIMgfTIxPqmUP8/HS+Ju3H
UKSGhgyD+TgCNclpsPz1LPMWGYJ4tSpGxVYXpkw/4Q6f01jP+J9TfNSJxP2k/5ZRildL3dD2WSF5
5qeZf44B/rPrDMb3M+977A2jR4gR2rpoL9FIKt1N9x/JHgvZsHdJWFJLPer8j5vwRcbtZxh4qoxL
B7+K+gt50m030XoY0VQoeoeuGzNYNsxBFsxvfRYeBMpBo+o0dubrD1e6XvFOcZ5YZOhIi7iaRG7/
TviyOzFHM2yqe02d6YKfLTYla3N0Kvk7j4IGSQGOsXQ0M7fc8iAHKjgo4d19Ny52I04vGBvtjZl9
LdyHIWx4jwTnwFJXFdSuCw6xtuqFlzevMgPX2p/rKmgL3SRjpr2ZoxtnuhF7tCahEhao5cjl7ODf
0GJP4HXr408mJ8Rgcw4gdOIu5GAFsn6AlEOpC4CRukmONNPqe+ueCBMphlRtzKVeNGgEX6WKru4t
HoHb0pphYqvcuDKI3RToO12IdWt8WT58en3OCoFF5yKn/4Kzp5huy+KpAUE8xvzmW+3lafQM2Kr1
BoNCuWN/JAvfy4cgxbl6vQ1NBQGQoLtqwCltW8jC7nYjNbkq3rsSsjGHF36SywEbL+glgl4bzGlC
Pb16OlWZ3ttPMQiHttnlhw8YhBtmvj4YLp6FnP/T7eniUKiTmsJgyApgnHHaUBaYxvn7TuUVSCt/
1UVrruhvPSGKir7VpaupNsWgVGRGDD3qCUPY7rxzNgqJqbTfe/EYqoeEum3SL247OItXUaAzuqaY
SmvWFr3TOns/eUZb/4C+bbcHarV+EnTWPcu7VGhJam4yTOx3SuUD/dR3iPKCw9kFJl0AozyF4xsF
gxFB7+1Ack7C05cT5H2fZQSnrdLJ6t+wv7sEM8Pt4YkQnudajstVAtqkODJyFwlAaNev1p/BjoTn
CvcoPZ3tdFGOLZ30DCVhQ5URovvewD3RPntqFwPAigquDcgBJ2iiUH247zSNV6a2f3YewxXeb9+q
ladRpYS/qrokOonF5dT/1qWSKCrnsr9IKVN1fnP3JgFNpC9xuJa7L9LlO+dU40OFjqLiU3vZ2yzp
Xk6hY8GtkI1VESCJtX0+yj0MLceeU7MB6uzLOM96oPxh5f+PZ5x3mYMmACwb5g9+lKGDPt9gRn7b
EHyqNgMv7DVHnY/gWvT282/cBU22xvHHqTgT8HzGyRWvT6gf5sw2Mmvvkj9lo/AhGUczQvwRCGSt
5xnm28zIGzF3kvqIhaOF7M6VhItHjaqUC2o1u0TLaufrAsXzGh0kGogRQMqOPhn5IcZ+YciSzytJ
S4naSoSMUTlxNPd+Cr1KAUeX6MCaF581d3qydnPRMtG0ZL9Pf93IJnCW02QaTnPigZOrFQgh5b95
o2ebkzNv4rZuu4HMwVgPFWh4jfrpFlr+MUfsqbrgU1Mp5AflDeaiuch1awDz+CPVW/msXFhuP4Pe
Imfs9xNa4Fv4u4DDmCST9c4909jDX7Gl9Vo3KUoiXInusfLp2iO6ji+DxNbUH6Dusbsxgwm3II9N
h/XyMQlX/4AOQTExdywxZx7dgTxcBQTtXeNBvZCsxE4tMqX7ZCd5M5BmjPV33VfD7NUt04aoCbDI
RR3jtzSLDKkinsmIMYpkVb6sh93q0RDMLF/ygUqFzNnJm3ox5aVdgXfREXlpCMlmxYBD3L03yIGv
4JiC0B/Um1ADPxckQNoYy/SWoK76Hw2gKbgbBcf3rU3wFuBhCN89qWRrE35K4YrWZd6IXYSeEAQP
vhNKxc+nrFVg1mlJfZR9+yLg31cxwGubCoL0+jJMoosr1h69EnQHmBPU2+ECfUVZNcCR9TXfSKo0
U3s5Cw7xCLb40HkDO05LjicbZi1UGCkUb+fwZpKBQuMo9gXQgaY5r5C80CclVmAGztoCJVxgDy9Q
A37PVj8qNlq7Aqeu6UhR5HwvUFipvIAUXAOVQ2BTpG3dgwHfbgvrKtZgN/pymCbpMYenpDlaV/OZ
v3PBGYwhIjSY5Z/+JM3lE1xpU/fDCDUlBYXsYKg1YtpPNVuFJRFGLjzS46EBHk4o1olE0qvk0u4P
T+2cF8qw7Zd5Mms3/6uNmiTfRLx4W3DsPHRQDvnE2qTMHe9HV8Gh/1M7S8VP6sdXFPxxetukyAjk
6I0nEmry978dHma8EkUgzYZeFWY6bgtvllUIIUWUKWii12VAIa4SfQJ3l9ulW8HTIbwxk52/+WbM
r3kERg6Vj2ovjY2jdNpFrCUY9q3eoRFzBBsAymGPCRKsLkXu7nkRBCAxj8W3vfi023Ex9Ko8JtRE
fDaVf+SaYiQOqPvZ6WmnyBYcyK7/Y1RRlsRUhVgZ1PyXMwxvKHAufGRAlxeQbgzPGY8yZ3gGQgUm
4YBgCxO6NpPympXqtlxnH4zpLYnnL1WfdjSht2BCjzgXFMI8alwhuDeEwiQ8sdkBQAo8EkURkE2I
HD/LDxxhoCHMHvn9j9MOHnrthDLhcOeGB4NaJUCWp5MrVBwl+0gtyzYqIzCfVLDI6IXtr8kR6vqt
IEEsoqM978B2DB10FyToVVgEOHINiSWf4HCjINSSmzrXl+PAO4RyO6iND5O/mTIslwnYuC8ahP4V
yb5ftCZR0O7ONj/b7KW9vmOp60BRLrQ6CJG0Yp4B5YOmYVZ9vJGzLnQbFmJUOlmqx4DMS8yD2mIC
4Nj9+v1PuTs8J3VhrYoSZIr+uTd3M4jQA3RwjDSsIEFz4H0XHbDhIu1FpgQouR/aJNpJhGn3j1oQ
/G71cxpQykobZrEBQEN5PuErk5KS1tRTZJnL8HCgqUl5D/6cS4bP8h981Nnjh76s77Jo6OmOjxbk
i0puHHsKhZgjN1JFSoUIY8kCLE7NuemZv6ckr3kC7jDn8Xh+Rr7272pvevB9cOH5boMevTEUyhGn
uuJELfKgspqjJhaKLhx9VDbh7ZMBfbha0a6kq96MbSM4J77f06JpugNCA1RvhgOXASpu8/yy2wLw
rNjjpMoQ1u3GW2rgLHuKMTJzksPxg1KxEGJY6VJuldGIEFgapwObB8QN8T/lUu6I2Gy19juf6zQN
UwZ1qwR0CxPc5nRZwidLQO7jSGkZgcCXk2k1bHx9U40kyRXcHF1JhH1kAAQxHbtRnXDDIvFpGrP4
vlFkL7PtXtVryrPaJLeQQf68K++bXQXRzoAwlHtyEodmbaNLJD4me8+pDd6jI0ZmTvzeevK/96oe
Nj51OR3V+6JVEZlH57saqR6oral3tDDM31OlK7MuCNslm0sA09Csvlai14iPcdZo11aFMX/q/LQB
DXqvnvw0u53vhDkO/I0iydxIqq3kNM9vE7kNCCj6xbxt60sHMl+A8IGpFCnP9l9rd3UyAms3qGjZ
/uBWu6hPpimqQrvCzVME5PRxU37SJHl0vII8FVfUQtDkf6pF0JaTkh/rv0uxXAwBWhjobh/Nz7yP
rFwxmGpHjHNlpiTgivgCGz2BsIuBr/jUltc9boHweXH7clUhmPxN3jl9Q3mhQD8TDUWFkzlQawoW
IiCUiLvGfCP1cnhtGvMlKs6111qMp71AsACoGl/XQ0pZMG/cgqDHCo5S+7zfv0n7CyOtSRN1wVbE
3A5jQBtbllgtlK44rnbY2aUGfkU7Nn+lBi6O7+aorJoJnIi/mVYqRVKCGZO44AyIHqz21ByM0fwT
3rxspgv1kSDYbX+O5hQtVqRclaWr4BTlHXU/smis4QQMebr/on0e5v2GC58ydIZN9Xg21d84Ickp
8q0rQ9p3tngzfaHEAzbQifF/Gl1TfsJUF9nahqKn/mtGHUJFcgXct3qk/qm5QJUN4gVtoSlBD2gN
Oi6ucxaAhOFNWPaC/S8qJGcGW/PtPjtunr0YFIrgagduxwda9ptkMQtZsG4m7Svl9Altc+Wk1pkv
9xe81my5w7Q4mByzeBNlAKjOabK5B1V9WfHzq9nKgTI76NTQowqqtihCYdv2e4IPMB0wF1gWnNB0
iHlGJbku3b5JMNnDVQo08ZbQtCOkhr1SByDmq13mOPM10NPBAEKoJl2W8aWPyYDYDfxiKu5LViso
8mT14ZPEGo/sdL0tZimZo/5HJlAO6BvPhecGe/2+7qJk9Pf475RTQXMNFDYDbZ6xcr0BSxsy6HZY
aNK0Wgw7qEiMo8TM00YVGfRbhDrfzaJgNqIRKwLt6mvhfepulygyFcVjSEkJoCITo3UvpXBLgpQP
OdnKVGHtTaQU1+xSBY3nwDyYSu8Tevnk5yGyo1eV62oq3sekS7GGfETFVE/DugZVMbiyjO+xuzav
+tmlSFYW20V187h1tdKbfyCH1iXwFBjPOyFIdXML5dLparnY/He/C52CZLp2LsmlYlz2Am7EGml0
yYeIsJOgwNqmsk142ooLxbv4/WLL3DTL17o/uVbmO14cqhlvwh7OjqozY8kcIORi2JxGf9L1LnLK
22gSSphQCLMOFEgvX9M9MmyUIi6fToGq5W0jNkN1h1GX0/6D6IVjdV4l3j6Mz1DwYAoi1Ri5fY0w
+MbXMd7HSuoy1Q6cOgep/KDFw7hTin58SEMUrNTEmgyS0tZiljPmzrT9iJ+ipuSoP+oKRA+Ftjwm
zq9sZniwqJp4CXFW2A3pErgwo5Ru6pgrMv4i1JON3fTs3P5lxBcLzAZTd6sePa3iXnFySaOttH0+
lmMaNyndS5Sp/82aC/dY/whMI7bm3EAtA+PQRg/3HUC7zEmmA4nmvNlm8eeBZWokWl0K9q30/hst
T0Az8Wf7S5NmutkswGV+UY73GLqHATutpPCY/lAKZwGsCFjA4H8D/cNu9Z7kQYsBopxIbAy2YBM/
Nm6MOMk1t5sMbl62CX9SBxPSaJyp7ZrCJ2K94FDasvjbI2OFs73e+g6sIFU2JFTQu8v+f2LQqwbE
ue9FiwC0LxOCJBuTWHd3bWYS1eHKbfxjN17YigkwQ5nhai2gFZgBhh58xDp8m20/+neCbBivmQbD
dAbl3rzkTqTRfE7FbjKZBl+qaIEG2o7fWdQcAkzYYGM4JequmPS69uYQ5cFzMnz+wKY7wsg8u1YK
fiaB810Jo6fFDOVIv/cI9v5EFJCafYI5FbIEZoso5rfvU7TBOcdVvW0SS3x9NTyNhTn2qyNXeZuo
V5MPnsEZ0dHiJWQKMRT7jMlYEiBxfAYmghFXoelYw8f3qbGn7jFFlZl4xKIv038eUWD8DEdIRRUz
SNRo52eFOwbE6IaFIWf0p5vmFWzVqRQkbXfX68IsrznaXxJfbjoKphFfb2DbKYAympo0JjFfyKdA
PVXjlz8f+0f/2r2kADSkw0nvhqPm+jsjA4xAiVYO6NyjRFlzymMyLCBAPS70iV9JEn4s0t6ScFXm
C8VpfNynMYxEx14OB2LUuaNjghMJaqKvxFY+x+FKEGwgAhZxrJ3/HTNXplm5av60jZKxb5E8Ixt8
dRWehAl0HdRmXIXlkMtjfjW8naYHKCQGMAGHRTGAEmcGjSTlfzwx/dKCFr8lHf5FXFpTUCJHQKSg
ube+IGaj4Q+OOa9Pv9pZlfKAKNq9MiZtJtBoKNnp+3u5KXeX30U/LvMR6ltWdqfvUzYTA0Movd6F
G3qujr7qVEwKLKSBrdY9zJoOkKNKhWl1pwkppBQ3mDxYFqOHedGD0eVYlDiiX/juru0VZlpkhL09
q2yqaLtanxNFoxmUHRNlFVzYI3V8hjT9auLQlTWSBJ7jUb8hAX2bIvGLgXWHF41q+BsQyItiy7th
c3IQ9LPL2hm5c0W/IWwdn9JpEc0Xxeb7SUYfXpMAp3wEj4YmHNSvP+myZ+KZsmZNuUlDk2d3+rSj
KUgDYVdRKQ8/sLylKiQE2dt9icCEex7+Btgk28m55kHzVQTFUJFNqo5LId4UUMOvvAIvRgMzDd1q
38j7l5Jil21WsqJ1balg8GiLjigWKLmFxQEv/JBQg6ADqAR8mXfT5wZEf7xIyaarTfrla41Af4qN
EUR9VBTkBURcCPBQipeC836miUAMR8v5dEhfaf2CNWbmjaRMgj36+TLrWc2h7KGUIBDbPom3Y9u8
W4Z35VHgIALQyXncNiTqTvSymuI73O+7u4dCKIuWP81mHheYX/hPBn2F3gkPv3XKA2Lo9SV8xyzG
i3vXuLtYdG0uzPWO9twAke6HRQGy2QOSTZCpqG5I0yhRupmMEHB8SClk0UAmgG2siYKWOm/zJeBr
47B5htei6eV8EO2t4SKT/cmesSzUd95cmstGOcC7BUMbxMFoPOfJ35z4BumFxNpAd6wKmLZtiwgY
FjBVsWQ1dlV+ueCLno/fxf/0Zqav86eqNsyOulQ/n6NyoECLs8naqGiXi/UoUwHHaEWJFFqECgCz
Dacp2uZU2NSEfUpV5veYebczWSSZ8OZQS0t5B3iEQxLd6v22fyQDwcsuUv4A/FubEcbnR7VpgrS9
dJE58UqsgNjAvjf3xoF8augMdjGMEotC0zlSsj3wx2jYgvOLOpWV5phVv1pSu8nrBZuqoMB7LKOd
KqPUXJR1pDv5N1EEUx6cxBtsSVAukYtzz/kJZJha2gqYamrA2b8uyuUrWJ4Sgv5B4RbSlv6NtW8t
+nV+MLVNNewze+5F7M2vtETcQSS01F6QVQXeZQaXqaIzO0ndXrZsTXskq+7VepoB2eknroW+zNuU
UDWSm9t+cxkAS3FJJSuOsj4E3eiFUKVb/41t9WLCZUMluJ0DQgkI7Jf8mRjlLGe96gqu+zk4n4rQ
2cgQygdswUNtGZhXoidEJyDlFMPr4fXQs/rwTyCvIjYMexR2nWImk1nlWdWx/akAE8wS5OUijwPw
FNT0OwEHkwlhLjSuYneW3cNqFOAuFOzhaGaWv50BNZs53x8+YbwjL/O/fz+428cnp5RAlUgwetnT
0+2l3A0KpVHiqkwxWGDSvE+6UuFcLS4GMkWHP3tA/rlVYow9tsD3MIJnrAK7ypHtuuDsOFYP+3w2
hgNlhuSt0HG8OuvNTP9DhPkB30t5kmrhOlO8PRhv2uWizm7dHGq2q9mwOHzJmpEQ/HzdQOdVIVwf
h16uNo90HUV56LgzpPAQpcvsp39tOSpraVkdkXQZk+4jsuqDqm1hgpXH86/m/FG+Ub8Vyonbt6wQ
xYf7/dZqx6XD20Oc2TRd6raEAclfuzggMuEdnmk/aus50ow4SOTuPyq4nueaEmeW6Vv7tdsVvi51
MugC+amXMVxYJByhf4ELUlZnkRAjIV6QoRGqB1qqwKEdtktjNn++Zc8qdLS1/SWWkCgVcBUzJIGJ
CFnkRy+bGeb8Itlfugoj6R2tsYaN4+1W7xOh+LQlquTK3xbgFx6SLKrnG0RACn6Sf0rRCXP4Over
Q79r9wdub2G6qxH25dafVL3mCn6BiBFa96zM2puP4E2yfGWnbh+ZsPaEZBQha0d0nQUdmEceD0qj
9gM5LLJSTIZjxQtDW9ScViisyVZ0JM7sQ9QkOZkhPLxwKhiu64RPvIaxd69CzqKzUNX3IvaO8br8
6/VHjQ8b4EACTD7954Yoot8UPHFuHIG6gi99pdBssUCLpzRDP6llrpcE6mNxPpyXnLHPAUIPk0jm
3gwDeDySOwO6EoEvADdXuJy0yLOlra1uIZwygUGyJu232h6/UvlE4lu5tW7FnJ6AoDoKWmBFYXzy
Oc2/+4lXJ9JTmJZ7ZCKI6UJBaFdYqdK12GibaEnoTMEHzYfoFVSda8HcSAEP9ZrJgYinih3XotHr
A/FTOGUOvLw35HA6DgtJhB+A/zvYNedQlHZ+5UnuBRRyc+0Nv0WLV6sOBK+rtzKJvHbCVQwjRDLD
2cp1uqRCdXWIO8mb4ePpkn3vVcN28Z9ayf0NksITTB8m9E6Jg6Hm0423Oub96j8FNr9BhrIKZxpF
VUy1T+RG/kIbS+TyNpbhOGlDJ3ffxWnvYsAh9AxnsMxuW3Klt7ngYrq0sPrHRon3E1AEB+w1jdII
iEd7IrAqURgtNZxaeeL5GWveLDmzeJz47PbylFsglKeaRrYZ3WbZbxNiq/VMdYddxlOihOYz9Szb
lQB0A6jsIesvifc5GFERGUcUgjKnwtyBtCZJtN4chgykGZvtnd0SeMt7wv13mTnZhBqAUgRo74l0
scNUcT6xBnZuVCPe3nKa+mXN4Ks8ZhKku9OBsDEaYTyt1Nqb0ziz7MmJ/Ysl0FqhJfZ/hSjkZu2v
bYwLSWEK60hpmre93aazk+srk/dJgaMugc5+zevkthD+e5CB+sUVmgfWi5KM2OH9aCLNX9uTAr8f
OXZu+RW3fQmbmWIDui37XJhihrHy+5++wsj8fNx3U6L/WVboXTmESbOSGI+LToww0Fd2X6TwOw/V
idMGBNmlt0CjhdQtwRgvnplle7l900L/BDTBSL343DhqqjXoCQ73f1YZE9lkfkgJYUvzHhITznB6
dnJouztPoQ5Rykvelbg61JtjQYB/luBKmvCMvt2LdXF4a6ITss9gKj5XUYsoMy50Si75JkvDK/AX
VMge6ghrNdqE2qLpdHMQRpHujXsM/h1RemLWZ0Li2B7YHWPXJUAuMeeYiVpzSSh4cusk19pk3g+4
Gah8t6ZJH8Ruw5N1JQF/fcrO0g7KWGez7PunxcSjiH/D6CHHqww6XvvgmPp+TZ8UXjxo33KMUNAg
k2radnOkDk1xc9kTCugKqBOIswWq5NI4zoZ5H+Vjm2hhItl9s+renrkqKTKYav96dYeRjsryIajx
L8AAtNXmEjlKhze3gVKK4YMjSfejoVNFIMSKtD9Db6zf0oIKoImU2dKK06xzbsugmch1hxCRaWfJ
x9L8nB/2kTd0+1ai/mNiWrtWuHdNsSv86c0Yt3yhIysmXI/JBNKH6Uj39t2pmUcBi2AAjUsCE4vc
azEqDF+LfdHIkRZnhXwFRj3XpVTTRUXJX4iPpGYX8lhbQNq9K+onmg61l8J1eO9JYKQ21gnHB733
npYJsi6ZUq+Kshg3GA67aMvCr2JvIW/3k0lgWWi4lpxfBjY2XOQ9kMAu2mPHu0Edb2fMNKBMIps3
T6MFmcfs6JCVc89UYQYOiVkLuD+uOILxXIQQitAYPQW26SiN7Ng0TkAAibsNIhnLkVHuELHq05/O
y0SFJYgVWrIRrsO8HcphixNrHHBVwmr/UvAddjo8d0twV9zy33dd5kW4pyEMjAR+IwOe8JPlTVp5
QhqCUPG08w9Cxs5wBBaL0S4n5SYlM3D3SnUD8xG+WhwR8mXl4XaNn4OanxzNPeFwRvSBMSErHq3y
uWusjNmQ/Uy20udI/19zNVkjslbpfquAHWRScjDSupbaiF8UltF/LGHY/cIV/Dw72hAc9PZr4Ej4
C7hPkZ8l3txXMZfcf8D+mgK6LXDp4BJcFNkfN0dcGIXi2OCZNva+nzLuL+F0QfCiYKWphvIciZ58
D8UKTC0ga7QwDYiBKAPeYBZvWDovHCLViN+yu7jxi7C9DuXo/3BiNX9KMjzs1tE+DHPUjbxq6j6S
FWx5H3sgBGbhoJcWrzWqiCdxLzK47EH8pYsKJkVp2+gIjnkEb39NW/niiSGvutRlF95d6XiufBxs
UmKm4728kbuDOwXfz2Y4ol0H2qoaaLBhh+gxoaDURUWX9KQ0/0fmfWRAsfPUU8Eu08K/4S9/xKAi
dDx6tU21slKydZgvpgqwcrHyjH/w4KXslkYTpL9gbf8eq01UKhvK8SdekgIwXZsdLOuhark5ahJc
iJi/EEjR4tRe6FYyCsKGurH7VB/Nl2v49zl3iv5WDftV8G0KI5Il8X3LUiSOag4wGqC8fEXreQd/
2kFaFcg4/1gyalHi4XYb5ADWyvuOK8K0AZl0g8+RkZncVCGtMXsZ3JeVZq6H43IJShZbZSF2ReBu
XUnCrVX+ePA1FpzNJr7/VeLrcm4XYD/sany7uES9LEksLPtNXUJs1LlC0Y+jq8RNLHbi7j41GXd2
GYEewzVjWJCoJFYzwLreP9kARm30IdgIKE7YwFw8QnzB5ahEaCu7Cf7LzwSiN2G4xh7OOMvibVfs
MtvU9tZTaI0zfl35o4HbD5qzyK5105YWGdbLhPE1evHxIhVSz8wInToMo4MBO7NiSjX0moQQdYrL
z5/dPuRNe8aYMUEZMUsjDvA4TLJJWdVXmzyLBHQqPVYuwmi2eJS52aaPclMejMUaVHzPlDsvJDPk
dqzfDv6rG36+9G+q+juyfTVwlRuSYAH0NzRrkeEEcYrjE889RMKcQCajKfR7u4Yibg1BBfvkS3pg
lagdG+Bz45n9tytGDNrVg+By0rn5lRxm5i5H6Umxztr1hSxwLRZysTTfu08I3PTgnXoJyss7GDpI
hFEutf5sNuQ9EOCCVXrEE9nJLBvVMbi2wRjXlmKIQq/tdL/0571/PuGbVYtp0qRnhIwCxj9le5sT
gY4qsUWaPH0JJvY7nI68saBWUWzBU1pF6IX3SL9ZxcD8CuEOsG4cjVi19ayec7w1b/YuI4wOnhhl
YsohBkBwCYcikLiNyH20+px0ZbHNA9Fah7WkBu3chde4E4EgaLf/seBUShZD9h9Gwtya9eKyGfn7
/gUd3pxejoYFEv/duvAJLxYjI6TwTtmmKJm7abkzmpt0wEAtaYsKias7ZcLUKXiCWz7plLS1Jza9
XWa0rXKnBTOkzgY03kQS0hETE3IfTFcC8anvCKzsz++O63ArwKFK+8f1TVMzQwJcbMRwFiNkgwNj
QH2byaisTkdAlkoGgv9BDMx0dklenWaVs24wimykjLHg5GbG4Pue7AkriqfelsR3nsV7U5wyKTyF
V1A3x+zLWJ07O2T5BA7G9aPB1jolmbtGRH1kCO4VQtcR33bXh7zj28cHkW55x9SoFAjHXZXDiSO7
2gG6OXU6eAjinE22C9Q9O6zx957/1w7ZcuW7yWcgEK6/aljhZDADmgomN/yrNxhNGZmR1aTyjDgM
B230NJIlPGGQvuvSs9aSCJsQETU6pT8L0vMEsIiGOBTQqfne5+THHE5HKmSbn7dKlULMfQzheMnS
M+KOAuonc2ijjZVA3owwCDsNWLL2dZho42H+/8yPFB5iDEhseR6KW59vwJIwmG/VivsJurZF53o/
4V1ZsgPTcF9f+Q81oVsTTaO6uDtjp0tt8haL8LLwQatLcdhbEa3ovv+lYwzZnkOU+Um1xVyxISTV
OTzUEB4PFoiOJax9s1oV/hpyyYM7qGwgg/SBmOTD2VciBdwk84QzAKHWY/2YMg2oP2K3NqyrH7Kz
/vhZiSG1gWLPm0/XxZr4Z+LJqtVkKSqxZEEthVP8ErGV5IwbLFY0DotOLXxYkR5sBzV0W+DDpjBe
Z4v0IB35U52z5txJmCXH3nBftFCasKwcHAV/vxCDmygxO8ircYAufD8EnytkMIY1pQWu1L09mEbF
AU4e+uOXqm7RU+Y8PxP92nm89anAoHhRpuVt/DmBPs6D4zi7HRHuGCRCve7AihquZ9P0osw8JDz2
kwdd5Gq4crlWCH4wVPWGpdpiBo6hce0CPphtDshUJUlmsF2SQfvFJA79etPPq8lKOuXrb/L/gS0A
xLudoVDc80KZk2PNRA0+2zaUYL7XokWCIK8CTBT7okphFfJ2gZ2NZapvlTyMfhrlzbZIzU5Uwa1U
qLIzJAh+kyX4Y5RUBLnds0mKnBvUztodR+v08XcRZLknSqCQ3FDMBETJmj/n0QEf1gDu8OJhuFVX
gTb7CtXVpdKk8wrOoYrU9vFQfPBNX0uxoeeM9eJrYgi5hHq8m4VvksCh3kiqUragTP7MF05yaVYo
b/Q3aUlvMbVdCIlkYUDAPRfm5QcuZptnq05gnMhv+qLhKsqalCSPzFRCh18rnECwtQmkmKpH4RDL
W2DYtU47E4Axo11U7JbWfWpjruvGSovl/aNaiLgJOd6JHlUPl9Lm/upgIfWqUUtB7fkDxudBwh3N
mdqKi6dCiXqAw2KOrKirx0589LAI4UksZXJno+hyOmiTPscUKT43/7azSrDHs6JBBCcJ6xAi0/Gm
YPlPatZSA/n8bl9TRSRgZVbrf9nm+vJn2GFQ/+eqLdllKyU8tmsej1QqHaOVH9GgWX86jH4f2vRv
gyUkBFoSLLlccT9YfMm6FGgqpBK8I/U2G/1ooYoJhx31E8ib3c05HdEjpf9B8v3nQwlR/sy4PMjT
udd3AAGw7bKhK2u7pJIy4DxT5atnlCdo++XZCmQlX8484ZBA7W8TR7i4saTTLyjMyyL+vULMuxD3
5D5Uqe7+pJrNUf1UOP//9+DdlRajgHuhqmDnTrZEwYBWgwPdmWRhzGUoF9j+qnccIbvxERXygRrr
nsGvEDM559sv5/Gh8rMH/7Aqdi3YE4j/KEsabrScmmpZlJkUsDE/zgBvB9PTjOxdDkuL1f7JyBrw
HI7BEINa208wRQLhPkbxniYQHhCD2f3HAHDJHNfEBaxStPwHvEVrxq+GE4Z3v40ZF+mRhn/ZR++e
1z+gxQFz4hAWspiNHpMtCpTE2AUX7v7krnsw7UReC72ONDKZWo6vjMbvXjK0l+TQLa3Z7U5mY3VY
PpBWIX2ODoURQITegjhcmb9xUxRRVQwdjc7wTUKMCuf15C5+Rs9jcR7Ays6TV0V5wtmbWXdo+TcN
s54GlGD1vF7pfdw+WIX3Uxl7SlyHmnrG0e7L8DT/AO0FJGaM/y8Xv/VJgGM6zjVzivy3ATZABNfb
CrGczm4JIB1JIm56NGSntkNveONJf3cXHeXoDvT/H1ermyEpP9hvyqXaNtRHzzb2mbSzUiLs9XOe
IeIB/19n/JZ6hfFKW1ktm2WDP+qszNQA15FeGBnVuKCWw23Hc0JoUm/y+sgYoixBeJKdPrGpOw85
DgHQ2e3sJHxiAk5QjEOnSXht8qruP6tJJX8SuvHon3mgZ4y4WfDqGtuGYY2CZRCJkJ6pGkzyJjnt
UCYC1/v/v4CKmwTph43WFyXNJQV+USTEMVRNGy/hkcSdcEjMzxDdl4LZ1CVLgHzzYkco4dt3NN/N
UgB+r2tCraIn13nmNMBVDPyHHNAt1H1A5Km8on4cdNo5Nni4EvvV+amY2B0IUXU6qg5vqNbc0Uy1
BXOlTAe19BzdldonjBrYkH5T6j1ydHW79IODp3Q3lhMUlYftKrhyciTS+YaYx20IpanHBbePInXY
W9cwtW8r3cb+3gDzxDdSsq9f+O80YJwwOiOfch5uoEk2WnUxBNpi0HdjWZoEjBUzFB/QrKj48Xbw
ZL8T846XAl5ttssbeE2DFQduoSwNp4Hq4WCh8AL3YYmcJQU8JmlpW4Bi3t+d33VAXbKSNaX1KH+G
ZUqXuQ672K9jOG+A08T6DAm+R9RnoP0Qg1gGZ13Igd1okM11KK3xHUOj4KjcDghaSa5RmsPi2we3
pIi50S+CgFYBjGL7RtU7amMBiF7QmwnHgRSWaxeNwJTQeRgZfoOzVW+sDhI9NhMoIGbMvlfJ34tz
msxy9aP6Hefibvi2WeoX83+KF5fxjUWKxeRY5Gjls5Zhk9lP4UIQHIsG/RFgG3M1E6iRhx8EL2Gz
QujfSka1hMeEDJULu0Wl9CzwStajQN8kpuEW/F16s1vEcriBicmbqv9maC5HwPgw/Vdh4yUTw9Rr
shCHE4Lq3670ferNi9ZgUj5qIeVdDUadGRvCStdk/G90+ZLgnxslNH9etWdepj4YI1DX/KcU53OD
ZP8h3jZznGTXkXAnFEo92XABJu/Wr3Sv6BMV92uq3iSqbqN3lX8zTXhaqzKc1NxWZsCGKdcRYjWy
tiwcMTAJpmB9PW+DuZyilbIwoSJulsg7h9BBVqfZQD0UAlqOUV5LDlvGn8HDM7LXGWt8n9HG2vBD
ryMa1MDH4TXBD4+0USEBldpvKXVn2Q8k9T7uVSaXCrsJ0KVXYUlyuVgRFD7DhKg+1EvyzUFLmSNE
Tw8zZv2XwZngPb0MoPvm+lsYCD6QelkL6hfWBa0R/WKa47CxvZdfdqdwSmO6Ls+onTKUqf/XNvK0
ZubrJ6QtAKa6TLf4TNDvml0Kf71CFBCaPEt6Q/pcgHxEQwd0uGeir7O50J73WIeQGDM1n++kM/FL
xsCV1vpRMOina1y08Y016Se8cuSsFGNaq/cHyWKsGpnsszcp5k2QyBIZYoJsf0EgnfUe7G4UdlYA
h6pD/OABL/G5qmJ5UdVl6Zy6E8fupsusC71k+O6U1GqDk+dMYBZ0UOZZbqe0hSIIAMFe34RqZoua
3BeA777oXfmTSXEgDmu3phv5+sWbd8pTDc43jk+kngctMyjqoFoqgRo6rlH/1RITtCayoG8KamzS
LcS3TOwM2aczhlKCDxIuWPp2O8jx4pDflYDwUm9twdAnoE/MIU+IUhNiLCopquJR0O1sFMoiPdgd
j+l4N4FYQNHdCwxPP/fzH7g8A78CWlXTBQDpbSTz+XQpUIlu+mcQzB7PkhmShnmQYiaK8j+2eTHx
sk2wEJv22AxLmWvf3YgG2KvNTUPzGCxngucak68qgIoYzmdlNcPoNrfXCjNG2JVq8Z4uZteFukmC
chuPrK7GYRZDoDxRmB8BMWOB6AdBB7CHGdNIKSs5qAatKOWvXAD2QFCYqWpPRCMakzTt0QQB1CnF
ifoGSl4mPsuyehcEt551eWKEdMJ+lecRDgVZF5Qzo2TECE0z7PWu1pkJIDsavRbqtc0j2nHUznKf
5Pnr3d+o14vZUzwoMN6hp+vfh+Of5gXNw6+MgdojRPeIwJvx5fGcIM5lWuABdtCrlceC481YGrm5
+Q/EAm7pPHodaehlkYLW7jZr1OHf/iJQBCa3NIsljdDI/Hc7sRrjjHVrd043GYfDbimTbEb3HI+l
nfyHFe5rFVR97muai0c2sX9DhufQ/kR8tDpXyWY2VnAr4tLoCq2p6cetTu73Kc+AqXvFgfO3SeMO
waoiTfOv7mRBPbagFTtRacnsaP9+zTKxktTsWEBV86tmFwoNa4t2kyRjUY0EPEMm9UNs7L+g6Bqa
GHZIWcRbJ07tWgXcAHAk/+3PMnAiPIm3B8tL/dC/4YocIrp9xIyYe6ylU3lHhiUeibwu6plAVDyp
uUlpdUGWKSQyKAl1IUTC+yvYi8jpOH4uQps3wd8Gk4zW/qGpnaoatuIbYiGvq5TQKk97BIZGxefy
pH/UAZlEoUemVIYdepmyG0VtL8AZ5RKNNVV01GmS15OrjlF5hh0K+djfjBAl1X3f+q6nhxK2NaM8
e0QZgrnRHS/Uzb9qsJu6PLcknjkCs/A37U/xt0yOhKBzidEl2U3DDk0weSswV0y80lBeCgAESFJh
9Q4upHl0vehaq7BuR/nfWW5ZsXK8DvPHnUnaV7lwwd994t93iy5dCnSch0Zz7qHVuherLn2qzgQA
FcMbytaJAcYHiHfr7q6snbGpwhZgbFm+RhnTFANJfFdmpDAx7k5WbkjaKL7lKKDqjRvMSVKl6poo
dtqUQRLeAVd+sLf46AkkjkIoaHzMM5VX3YMagJVeOVbjZA2U6/W6WbexYkxchXDoWmaaWtP4Rngw
iEaymQhRWfyPtw4OPcl8RrxYu/NJAGiMM9j3KnyAqJGcchduWwD6MN9Xmv1vLRBWOE/31egLCDka
eN2EUfzKAQvb20upfXyWcX5cJwkEpBuT2fMQKXbcDDRkKQWF1J2dMOr2ElDmMAbWWW3LLQi/v+Fa
LJlvk4TvlWOs13iD2UBknP+6oaosTm0kFzrroPkfArsa4g1R/y30KkmWlzPw5Gd3bD8FDzuV4yTS
dwlKN4u2d1xUuK3t6A0vs1W0cKKEdvNiaqihvsAi5rgNNH5W/XkjP7fKFwZdTGWvadWt9Nmbp/xP
QfY+nin7PsO7teG78dmlDEF3V9xMQ4F5Ge8ooV6FeXPvsZhHHz+eiig7yHn3nA5K5q7KlVeXyl89
cKb0cK5/nC31qEDW8Tzurb330WfcdJLv1l2jhb+Ig9FWeaCkCGMWiLvPe08/nlSQtVFSlGQMLOmv
o8G8ta6Nsh8rupPxgEb4EJugFI6CHxqOpDKZQYMpoTnidL9YGe2SUGAh2cikzSAhL5qFN2EGY9qz
ZLYFa6/HLxMBXHFoWaoTDect23Fx4MrcDFqDs4t1pWXchquwhJPENgXf+dX3PAMMzTVzk6z9EPuh
XfsYadAPgocknapSLhrzJhV3PcNCQtmwbYh0fvEbdCp1GdYWlg+Pbpl7gnG6qmZFfmayIwAPJJnc
XqTDSWA3jreqhumoMrDIGK64DKWlo6MPDJ/YrPs4rcakwmmJ3+y6G18gt6TMMu5G6o9HIBTjAk6Q
GCz7n2Fkk6pOizUsvGq7gxGQtWeDG8zvZLOQvHdXyn1Rv4tX0TsZ7JTqmkzxCfAOig+nzMcuMVrA
ZR3N8NAoKnt6xLbQ1FgHSpAvmyHU/UBYKG7xL+LDoF6FRdzekrjLsjUlyPgtcGBwO7Hepzyfnf7E
fMCDsMfrDxW+kWHEJvaZCCGi+yP40LZBDZ3Io3YEjuc6XsVlglBqfbbCvvVA81u92tep3MmtZb/s
euXbxv8cgfbMV2fZlxTfdYY+F8wfk1+dCvNVW181kr1AzeuO33yIEVrbZHz08/JQnIlkkTN65nmq
mnSGvECxaFYZOF6Vui1tXB5GGf88mY3Ksw0auk5P38RGDkWHkOwX0UioWDl0VApyp+8Ct9QSxpSB
R0qDF76CyP7YUWXFdDeXS6dLlZitXZH5z15ojs3PrKSvxcioVZAcldAXHz93gymRXkXl/iI2Cxcp
s1KmdAOmZZpskfvKYihYsWIGE378+617km9nzJCuOLTDxAu5solvQEKMyLIj/hTK8hAiGRaxRxjc
7HZ0XFzoKbo90ILVyP6ycOME2xmprIb+ZlGa27xbnDhbM92m6/zSqkWYHSWoEUP4CuEUZapWLnN2
cCo9IZchqFQUqKrIpt+6GxU8Xy1cZnt41t2KPzARqwBxhe7IvonbKX6JwIr8E6EliPhhHsqFTPBV
ZYNoPzlWgtj/bntZZGxroNm8Q+GV0UqbuX71pvH4PfufV/mvGPKAnC58fro2ZNFmsM+QsSbsokLm
Ov9eB6heIyuDaUUx1qzWeALKMl9L3SBosqAr3uYWkba3Mb9rLJGLZY1C/DY8n4BWeQixyGD26TOi
di3fxhl7Adp3WdBtwGZtQy6txBTMuFRrQ47Rd0nNmqWznnY0vdJICk1XCHwc0fyrPTUDhXlRxv9n
yHQm//F/HR5N69M9YoqxFNFHqSfnCuzX62IiLl6HiWnzn0BqTOlkrKDizASIdkj0CyzqhjQVSrUw
mugP3GMbV/PLH2+SqlF6dmeLEA/0ZI3/GkFPz1zxnhL9f0LUt/30vmW09zbmGeVL0LtYyxeP1QXb
+MYzRVuZljR3bectdW3iX/FPePhucxlHzwWi4AG7sIiwJcdix0BvvO4ntQ+RfHO2Qvfg3NZz57h3
xoCwGhDgo+yxlJVFbkNDT79kmYpMDIc+fzst5XpRTyIOLDAJByB8QyOH/Ek9BD7kaA1c+5EFo8LE
lQrtZDbJp/LCCSaXxREGlOY2OWPy6R+5U9darBKZltfBNFO4PXWL9GIGr1Zv7ReOT3umtkqsklqQ
UwWeiB8wo3NwH5l1yNF+RNQviwBNBQWYjnfpjO2hoWDrW+5y6aqM330Q0IwL5FLaTP66xGCRkn4s
rRkkVsfoSAPHyQNffNvWlBu4RDFJwWEj8hpbH0cztTLXK/OHTn0Xv6ZcixJI/nia1s6J5JmwBnz8
98C5pc7yCI9mog3Kq64XFbK6YQ06mMd1VHIiV9xTdbor0J1XJ4ssLo85cnFeRRicL+u4cWFhekEA
wdA8ZAxkI3miG/yivvHh58z7M1d59sKwkpUEpBqIEPaJc6SjZNY4S41+FTf0nFc9W0XlUnk/ayh2
fN7/ZoyyEbNszYhKNhgLtjmgHq+jaeQdd56RUiZW+9nj7lzRwGXgGTBrsFY2CHPvVWyi3XEaqtll
i2lIc3w8gQGRGyE4fysu2seYLJL0N8G+3Acf/xAdmir+OBuFe4IYigqwGO0tPeAEkppAFP1iayZd
xiDLMPDADdsCoutvi1cii0u59MnhZ264jDWqNLb2oplkgP6zMubTSQmeuwosMFQMXNk7pZgsu3LL
gKL2nfbS9uyJ4bhcRIA8iPfF5E58IKOUyTeiJ4YE2TtAIkdS5lnKhU57An9kgj4jor6amy/+yUr5
M2lj6dIvG+S8DI93VU6yJ2sLI65mtU2TEHOKG++uuD1ARBpNmjPnkDQodXxPmLyvNXJGkltZB99Y
tEs5UGd5Ac2C2tiUL5n0lsDxVTHomJRYNdHrafWOndiGnpsD7SWMXV5Xgl5XF65y4rNQ8qrDSyCN
yo9rla9RW88yrEZn26qi+ox7464qa9zZhctTH3vWxFXbbUW3LerVYK8u7TJ4RZmc24kwd4DqqIvi
/6Fg/gqOWaIKvZcipfJNhQfz/riN2kIfj8qdCJqjUhSkLGnpE8rrnAmMe80jJH9NvShEa8Ab6/VF
sYcgFPnvJaUt1ggQnFMKnvMHpQnHo42fzh4Kt2HoVqgDA8BdOnoS5UOYbbmFe0tTS6dQ9yUsiaLR
qiyDvyslJJeDPYgY4rBTYEbvoHA2q/o7zxVPZ9zOpTihlPXs3wg0fud701Cc86rPSCe9YtXb1LeM
HMK2W6LEpzptExZsxfiyg9KF4XSDH4nZXvVKKV++r3pgl/QfmLYqC4+qnBLnY9m/l03WeJ7fE2UK
+xN3VVNOAPK8XPu89/LJ5t1rgAOrfe6Vf9pgE43QuyDB3hjwi9ZqdkPFzG9XoS46Cw4vRhJMbhzC
1vUvk5gISudyk+A86aA5HsfOFEY2URcYujW32XbaKmO4kQoRCodCMpLrGRWnFUoYaxwluCkIh3xQ
I3ncrl9ilYphQZ2ZFeUqBu8YByjP10lJuiTUjvjUB+i+CVkLJxnS+mbLOtNsFiOS6sE7uIvZ3qIX
Vw2IcXL/56X1FJQ/EStWxDKOganyksUPZBYiWRyl+P8ZBRqS50VrUGXtzLcvqfy1RDde9NraYcn8
exDcxIvxh2D40fx4qkw+D50J+T8A64k0uTC7mcxfA7gdT6JEzKxdQqRJphK0xZbHJ2lAmKWW3jo3
Eb8P1896TP22e28DD6iMZagammoIvghpmjs2UNa8lUWXYJ+aiOCx1gUMMcggC+6XBLxXCf5dCDo+
QBTlGe8sq4O7P+YS3L8VwycJA5A2HA1ErUgAMLMbGY2muN6i/RXMLakUtWWgUK6L7nlDjHokn2Od
tLe49B5QcArvaK89/bTr7rwq09QnSidwkFLgDEW54qdXK+U9OYha2PF9I+sVp1F7AgfEK4qRJQFX
oqy643PXxK5UdcRjMMkvZZfgyD5wZTglgm4D7K8EnG58ZQ2kP0BqmlQjGsSCHXMSNrgd4TPwm6hd
RKb3ofvm7Nlx0isHUqFp0Ymx/3xdGJhejfdVFFvv9smjS75iiF/hEINxovSyy8QYkReXjCMLDOUV
8GCVqa85N0uX33qu1fExuNCa/h8TgzeSo9FzoPCLhuaP2mB/b5xCbGlg9repggTsxPTGjHz6SY2f
u3T+Oe52la7lkhQTGqrNPL8CDb7nloxrTqVcxtv4/dOkbEbX47sI6LhO1RPaahDnFq5N4mCIEFv2
TiQn0YlQslz6fXP8v9x90fLDBgYt7a9zZh7fSo7ecNU27d7+GrO8YajEbFOVVQ6/nV3q2Q12E4w0
I+y300iYZH4dmZjpArV9422v+DsyuN/VDSU3/QDqjR1/1mVz3IriCTh8XAE6O4E4vh9WPe0boGeI
ookFO/QMyDGoSYk0qmAvyPu3Voc0KAxtlT2In/np2/B+FrCUDgLWbG/Q7OnG4OS6RRKpL192PKte
Q51M7R7zLAR5Pw4A+WA4sE3y5nl+9TgeAXLXgGm5I5VJ6m5ZDk6kuEW8yuqfTOMpH873pBg74p8g
Z2fY0FjyKTKdR+tqI7h77+FE1PEcPbE5BqkTGYC+8YoUhTk0Ont3WqQqg69bI23KHjiI+A91c+Rx
on1KEGPr4oxF98x8zlf1wNngld15z31z1JpQIo/GMCF0JHDQrI3Gt3IAcHMXOQFcasBIMhuWlcty
FVOVcHKucz6RER24nT4kSAd7HP/5+XS5QMJPe74Q6vSjfpepOIDNzdrZ0gRJbiGM9s6Vq4dtxPGg
iTzoil2wlQVaA5upo/UJDX6y7CyRDlkYWxj+VRTnpxY8LBPkCEBfPxxLaZW48U+o0BMoDJnNPABX
6s5NuJfRDlFRgAHU02dHtgy0cWywgpGunprczdi4XqCkx9urva0y52ouRyN2AT0ZsvviErHYslCc
A5s5K4392ya34n9ifOFkkLgFmyKanOaVasSuk0ddtH080Cnhtzw5qjdEQWtVTK2cGC7YJT4sou4D
YjBGu12p/QVsJiq7VPMa/z5xTWsaO3hdEHX9am3lwgl6FELMH6VxKombD2AUVBuabaJ6Nv2da/71
JsocGckt77x5oT5Ewqo59Er3LxXMuG5qZcUEk4074sRAzXkTs/uH3ooXqp44dygnebx78oNrOPUA
BDbvC5zGQlhcHUd3No2/vKDBlbNOt9yUP2djDFnoonwOdydGwc2s2ybLZ98SSAJVKyXkRCUExDB3
Or8zjQXmvUJ14wkshL0nhEgNGH0r5Z5jY1bVZP4g4KnVa03PQ/HQo5MFFPZ2oZUUiQ7OscWNGpP/
kdHXi4CeFjSxr+yXjwIrWMRSDPSxpT96CwamsbIeE+olqnzeXIvN10gPIgfq3I3VmdRXFkvXwqTc
SC2GEpb4HHJgnltwSBA5Fh19DACBK0LFfeyeVoxbmqlHxix0TV+x7iu3RkrBpjnO9XdlN1LEXh+c
+G1FLwvlxCrHZqe2soaAHlXAf4doIvqvYcbw+ffmlDX1AGXxRH5Cg5t60geIQIHpr/rjC8ChD+HO
tGu2R/ifBEteaz0uazkHU1X39/b488vVRP2SrqJCFCcuZgs0IWL4mkqBTsZAxin9kcGF1Yg/fkBh
Z6LHWUYa99ggXYt2ucDG6wnaIS3o66PX0B5WrJbMMP8fMfXEyuaK3hQFD16rlWjUGNoA7/C7PzIj
Ms9F2jorJNX11RDMnArxBpMAS3eUMMEOke4srmDjprH45RvyfT8Rz4xHNKCw7m6lk6vgM/8VgwPQ
E7nPnbtK0B5IQl2BcHIgCmq6Uh9+220/YQnz0Wfc+7F7QbB14A3cnC0+GBtdNnuBneyFOKLFy+Zb
PBsl+KsD+oFW26gR3deSNoAlG/fEzJoDTNwRejaOQnGoaZK516Hs/j2rrtcoqAfZRgkrnGlOUuXA
oXjl14qE/q2kz12/nvOCZQuLYzevaZxuklSnyJj5pgcO0uvYNDrrBlSq95P1nBpgpvs0eReEKzpb
0ex29HYxo6R49xdyiZAzVLAWGC4u9sFBRm/gedmfY8yTFEf5oGBtWvGd5ERmuj+fkPDbwSLHUpCv
66xh1e5rH8zVyH+l2+hN0jKnrqaAgdErC1WEdvXzwHoH4afIM9Q/SYnbZD1tHjop+uAJ73yewAly
lUIMF/TWsEFNd++eVm1qMX5Bqs0jpeErreBD0BiI0yKfT8taQM/7fl2o0z+Vr/XyPwz53I7JJJaG
gP17qNVZfViF7QaPbg9LM6ncVdYftQgsQPhmguWuYM6wleo/WvVu1GarvjUgQqH93iqpqcRoVUAQ
veAKUEbLtr5HR0LeAJ0TsACMxSAe7EOT44lHEFAYzosnQYDJiYDvZe/RYlBMgFTCdqPaCQ6bcuk6
HPWSTOzVRXNjmh0oIM1MRSryCFmX3pVqCVhSyn6jhzLfHFgwvZJUjn+OwdwEN8wTRfETNwh5Bmys
qi2KdVza+lHJ6yldIz47DcL0zI4z5WFm7SOcw9mmGEtfcg+bIAGNJ8DlwQQyUI0ekNaa/KhcZhLX
Th7aXmO8rbQVQR5ZmpHG5U5QJ5s+uQ4RUJIw9NOni04Ekho8KicdBhgzxVifqjYCQLQWol1iy6GO
PQb2/J0dWzbj7FMHgD6a2dtaUYZqmvgUnT/zGqAHOM4v3h9ZuSJjdmM/vGN+ZTtU1wCnZ+tscCMs
p75fk4YACYXna7I2sDstL3alSiheDY0h2UOJbjKkEDt6YQE6LEsF/Bn5aE02q+/FPi/h4CBoLcPQ
a8uY8lm2hSG5ilRrxr9bI8strj70rdZCuaQCOAENbhj3dQe9icJQUTRxC6IUkRFtyqlL/4WzdGSp
/D1wSdUbZ/b6byAa9M+CdUnHphCjIWww1IzQ8tUuKkCSloY2UMNBA1E0QSLPvInBF20nKJBMBXI0
K9gI160ANA5r/H3uqxGaA99DBpIM1+3hZuaFZ6z/6CC8heYudQt3P9SdjZsQrKSWfQrKyQFlNvm6
ei7GomIaQegKCMHmV/x9oLraI8H8p8XNYW0n77cu5ubVzc1Bk/t5gb7DL1m2PjbudmT/xWMRDd22
mo+BVEUwix2mdPYQBA/EGNndXcrS2aSVufN1+owApvGBMNAWQX8reTZ0azyDL12H8sdGcLtfPc6x
N+iC3cLE7XK1yAYf4DsQxSSIZpsXnT1udluw9on8PlulJzVuF2q0aL53cgzVE9q8DugXUXq8OpGr
69pY8EEvEhEwL5DyfKXVaaCNUqi825QNdWuASyU6B5xOTHnC9joaAYv7Qs3rAjaCwHkyLgk+6h0A
6Basze2BePPgs2uKzuWRWVWpKMYIuwYhh/u8AWBqdd1+5Kmkhhs/eBJR213xfRulwkchYo7gsjmC
2U2CuHeGXEsoLe1VjcB55rJeukxNoTHF0Ogup1UVarof4TUYyfSZbT58zwAv9labsskIDL68HI3B
F9lftfso2Wsm3VqzGbsHnUUNk+2Kx0w+SwCHhk+PLHShSSVqXLZYK6rbY+HNwr57EPsJN12zQRxt
A+gErLJRPKZq6yiSVqVEo/xCqWGq9zIiHhtlfiXm8yZmQ5lyDt3HZWKVecigriPnWApFG476OVn+
8S3ofU1hj1wCaDG+E6e9fZLQkR6sZqYaFRYiymrmWYUAyBLx8QUZD99oUSAqSwTLuVLmcO59ny76
rIAPKCQ1i7nYSq/wo0f4VgHQ7wSkJ3iCF3mGML7qwifrISd4ZjcqE4urmHbUNyJ+WK38Vuk9I1Pe
3UP71xzPv2ZfqP/a3+LFZYd08zdOckPQYWe6JmbUtujxEu4XLuJtheQEZRUfP4kZwqBtZPXIBVlA
klWlk9XFIzXj0xWWmK2T1HSRyzJ9PJNig4c+j3bg0QxG5oZc0OVfCyF8puzxkrakbGD1/xav0ec5
u0sswm7aKXJk3J9/v7WlEPYAi/XugFRwZAS0D2g40fBjKEe7GVH+xjHWrdKDlPYnJSu40UOvYImy
dVMtv/UKvT0KrlpsUs1+gl4aahW+wHLwZoFL8OaK7ptphvs7e6KZ5MXn7MfLvgCb1IkILJoPbuDr
zAMsU7mZSLtYNj+pAfB4ngJZQ3TpvP0jQR+imYzOlYyjOs2CWt+FHdzFRrFOG6Cacw/QfQ17yMlf
lxZQg4w+IBeB1xzfX3MZ7uFCivQSs/OuV7KrqTEMq6gMvrkjhB6XdQl6NM047sXmE+KLCn/edk3n
XkH1JvrX/h5X6ei6vPakYSQWdkVXXzu8e+fM/HlwP3kz1+tA0ra9Z7FrO97vsQK+L21FOq7Jb/Wc
PfJfAjK1ILJ0DinUi7tHY+hAn0iuA+pdTAi4nxsScocLhU/9EOqDoCUKB6SibhVpq1W3zl4gPnH2
v0k04aaVoDFUgnlWtWfLnxPJJkjr/S75GpuTKi57oOhGn6pUB1/YZjtxOUbLm+ovYvdr/Lm3VHHi
xtj9EWEz7AHOwRRZ+kK6EZYNl16MjU4ZRyl3Zglh3bxXMxjE0LBV8KUGV26KMQ58iAxB6QpAJsz3
sCNlm+qVKRC3FI2lIuyTadhJx1Xc3rLGtUXr/1bOIJ/XvN4DJqH8I+88rGtnXA5qmNCspL7MMlmN
tL7ZBeaXi3ai1entRAZr1ccfgSa/VL288e7P/0+KoZEmC/rA5/SGj/ORk3BrWoY6/sj0XnSRkeDP
g6wZBvFPcedWrZdG9Ch4YJEauAhFXLT+qjYHKT2Zi1DIoRkwOtphrAczWXWzyUj/ivxyVUL4Gy7X
zqxtT/JAn6kMq5hKigeiaUml1tspqJ+J5SiZ7F+uzYo3ZRXmMECCug73QUN18fLR624RcsFZCFMM
GF/aofLWHASKW7AO04d3qwsQBknogY2e1HExJdHtBmY4Gl2MO9vmbB07R8ABU3JVzMLGbN2rQpfj
6cD18YnWu7KtamoYi9kHY+FBdSv2lfK7nv4XZPVQp1ovSPN+J/j2ElgewRgnuaLtl5fJmUhGrEZa
JA6bOWrYGwv7hK9q05pL+bhIKx1Pft3c2+XqcbojKYfFGIjzx9B2hGbt5x0jN+GyrUkZOJfNj5QH
mz6toddkxJUhmB3O3gLxaOsmSCQQSqcYj3+m6GE9TKH/Z0jM1AfjE63yo5l/tBXXcn4Qa7DmF/gm
lSJe/42m8h4INInZafh2UAlXZo+BS+YXPKU6ik++HWLR7wDdcCFOsBJt7BCCnRMkpi3XcyQrNfnt
Cp2iITfXCi6x15eYbIwMuE+2m1andgsUxu+tiapa29UViy6ExMI1c2tlymUo/0SLTdG6O76cRGe2
gnamKJvp3ydWiMbuePaQNE83lm6efGpq8rTwEYLSnZlUI75kT5u7sGmvANzstvSHL7BeTwteE924
G/FZuAVwJ40L/vbrf9Yiwi0k1vpO8hyO2zQxt91N2h+jzAcP7Zb+7G+Yc4Y6eSpDpuh68YC2Xnor
Xpj2Z5QGLJO+IPK4ErBBuwZyMl9S3d3k5SF4V7hbh1nz3K3Dzuad/JbegMQTC8zIICsFqmWvzkLM
IPo4shLsI+4Ef6q10ohqHsAXOHtd2pUP7HKGFda3phIwZeWVaTC2ZbXC/bgihNB8YtOPSCEHI5eq
x6CBSbneIcvpyy+OWsHAf97fVuS+2ERh+og33/xNtJonB3oADxCLrBiZ/3vM578BRXxdnJ29ubqO
NBoP/UZYCxtiI5GDel6zgEUYHcABeEVsonZlo4g3tCTiShZhZQ8k/Bu9PfIyZTTONaoBT7I0zlbq
PaoOl2scsF6vkkvjyshF6DW4Ll0gEzLy/aKoxfGEZNCE9lZpkioHyTfep6DRwdgbJ23VzCRXgR+x
Ls0YqcdKPurd00+pBILsGAGl0JJeyIDvJOZFEqngbQAPhyvCrnecsI2ZxfNkfki9McDc1FEBKvUv
yHygViONTPKQeXHlukXtc2xxUBnkFcx4D5ZAGPq0w+dgc+/Prq7K27j/NZTMk8DGS+AdSC+MqBXu
jpQvu8pQqTPwZJFb+qAGuhsVJt9uS/EqGBsKhgboQ2Sv8BGuIZ7TNKxYyz5140xKH3PVnFfqAgx5
PuUP1czctX5VSm7IhqTO0F6S3xA4SYjYjDOUpsK4LH9rQ9F05ewybJN/OIAOVm3P0I27vaTDGPnR
WySOWATrl9FjvX1OVRFk2EFYoreu4nhjVt9a0CSWjmL8CkZNHslycXioClRRTF0t+rzTt7MIfziw
G1N4MuqlQJ7YTw5OUU7WouJdgRLJUsV9dGV+vtF/Xgml1Fi71D8eKwRN2gjU51zzyWqEW0FSQOgN
bWQUqPdrHz2CQsYefeMH63f3VPpKCUMex1qHT1VDsBdZD11ekpNtVyOxID6OyYTwCFupqAIKgc30
GO7ZL7RCdwFmREpf5A0PzAdUszIljV0M5eAxtDi/WeY/vqmjWllO5Jdg9Z5jl97y0MOyHI0UE0Wo
Z26GmXLDZ+isfqnrzModkC62R+Df2BLdkt+BN8lJ1Z9zWVSjEHkQ0EbWO/7/Y9sjnKxCLnjAzAtk
xng2pqfiRdwAGA1sw/u1vxZmT36SzGnUJbJLSqxwEpZdX6bRJXj8OEqocyj/mIZEqTGfz7ixCF8g
JZoA0gH8Nab+Kvmk9NfLnp/2mzNrE3msTl32a0WNdb3KyAJZybaFnz79tQX1qrIfF8SFyx1UAuBq
v1dEss7lprnXHXqIT+glQHMhIATA1yx4a77FvH3n9WXH0qHrByjKa4jBR9Ipl2IqZyZQQIHsAWA7
aLzedrIhFxLvAZZXYU2jw5suioHu92e1PrzCK9TCVnmPqNFX2Tc1XPE7f0JTxLgc26ACyLhcGYnD
9D1TNSvG2nA1MPLqg8E1zYmaO75Zen5ibbTqPegReAdofebDPRUCqXzckZQL2ru71gPC3BSkAC4J
qTj1DlFFu0YOVBfCvlShfSRnwsj/1XRihMKRibp3OCW0fTDIh3g2Ak4iPC4/VkvYbLwIvS4hmSiH
EncOlPfCEP5vD197Xeu3497trHqrYhETFuBJO19iNrRiCXEoAvhLLIYb8Yuy5JBAm+ckW871pjdk
nu3PM8reUq8I8D48Lbx9N/RenQfEiHIyeRhTQRDLSdoU28DXblFSfuBlHL+2lzIItcyoWdcTQB8f
ZU7VO9d8aguQIzGpR1A4EJhNDYl2jxGV3IUJiszzFwaC6FuvlkUaAQhedYT+mHpQMeU2MmJQE1s3
dKC9p+5xviPUL2vGP4OWhVRJVLODk8FKtOqtJPmxcB3r05y9jMesXMwaP0bxd0BNUo0qwgb3MGo9
MxegsInGvHl0tzttZWLJ1sKcqMMZxC7yUM1Xu+DH7zJF6cXoP3pkrQMIjU1hnVo7cIrqsc2f4N92
esVulM8A6UaNFQj713QE0wRi8ipzixciLGXM8GOluGduoE8y76MdaYrRSTNc9SSrzJTGaqzKBEhL
WnjSgqdyMDuFYh7C+Jm+vDsSu+hZZHNCEgYT3gfBqaD1TfRdD5SVJQ+welkUssVHcoi7eq2pKfMc
OSrKvQl+/MdM/pRbKdVQfzMX6BuNppF9vqGdE2WgdNv96DJC6msXfgZphEx7oC6vVmMyyEt3DlPU
p90JVzEvBdipIyMWupmeKR63Q44qvNErVthIjjA40MOKm1eEzYBmZ/oBKzvtO3Bz0i0MZyi7pH7g
tHuG8E8m70AgE2OpskKztmmQrWd6UAybT6S6/rD/xiepdrwZqy25x+tBRNH0i6Bn9MnVRVKR3NJD
AQbZTAycU7OOSQgitGtGrKXtAp9BNvM3GJEtMEYGj22tQfs+L5yVw4uNHQ6aJmATZFMNADxetldQ
qbuFQJFwPGI7zWs4BlBwUX6geJkGKREL85HD1IBVIP4eBoqGVZxZ/saKPilvpU98zjDIlF2k4WOf
wElyAoHF8boPSLiqSlEEdEHZROnfxyhE/tHla52t4pUDuqkcDYVbE/H5j+4LlczrvAF4KwScNiDe
9nIB9WmZM+BX3Wg64eBRF+dnFLlLPefmNu3NTpxs88RAo9L1gY53pl6ARMtWIy2Y59v9eCnyS8IL
B1g5uZ900JFmhagoWIEWSc3SYBvPO8GBVPPM4LvVemeX4y7FpqmvhHyD2hIUj+4SGnq8fDc4fWkk
ZsL6/QUIRiIBk56Ow1gABFFIKvqSQHu50lR7vrRzXCz3CCqS+BCt+Eln4RRl5z85YAjo6Mp/tMC9
izWrlw6BxEhiBDu36/21XoY7m6fThgpP1JBmC/Zx9Y4QM7IAJuuHHhuZfIODD7cwX2N3ieDMphzz
dhRNVmJixjbi4JuN9866t0ySdwYRWsp855A9iiGPwWOKQqaoLprNKroNmNYEnSxZXccpW72ZHVC1
XBTRUIOUTchLc30Iyngt2MJslZIot0jbNEYN5piLFjd6CKCnwPrtKt6eKY8w3x6ywUqMAg6t8h82
MxiKyxX73wlzuo0A+H9t23VXkHI5cGDDV7tRfmJi7CoxQyhcmiot75p3J7W7HAizHpQWQkq90ucU
dc7XXrZ7AEAS+09juoykIB8oy9RahqhxDQnaR8CwqLFJVX7NmfxWF/c4k7a/VTAdy4qYJZ6jCiI2
+xLQXznWYPa2MhXf7qwjChBgBiDjBFMAWT9hng7e9YkcgEgNABxv1hTIMne1scLBVJjoJzCN+4Rz
fEWpgl6Y33H/N/OW/tNVIkUaTmwYPJ9lcKzIC2O5/oyCuzWqo4P+blx3c0oUCg0u9aEw7npj6Ixl
o9h/MAXTOiAZw34SaZViPKnXt5WvO0UEYkds9KfDETikBAMBIhuMGqpIW4CSknL5M/PhLodnSovM
v1rN62DPeb6wa8h/sBlULmBo+UfE8lT2M+qiDahvIddJcS+b1dPis8PQsv3Yb8Xe2ZhILSTVEGqH
Bb6S8h+EbrO69BmION3U7P8w14up2H6Fn/gzeTy6dorzMwjNWO6TLaEnAZxwONvlMN7yKCTVdTvv
OT5Eki5e3LhXMJCyMgmyigiVTbd4huLU6PlzGh1fMI3Dl7n3ertn/LpY11aN8V6oT/qdcFgBy4yk
L22z6voqAVqOOLvEjXvSmJCwP4VChdLJlpms7yHoudIA3ESJD0lEtfpFTtau5APRAWjn0dezxq0b
Jcco76YkseC63ZplrW8iOm9J381mphw/r9I3oaOeRjKJ1jI9c9aS3UNSJ7+3JBOe8DQ6meWmYjzo
XhLiTwdiIShxZFkc//7msl6F3TcA4tH2rGtO/1XgevkvLZNuFKvg8fjcffrzljVY2h+wZQBhjabl
9pY0SYC/yB+HzDxNVb9WffH0PUwf93LmM1z78RDG0oNjuPBn+UdIajG++luzqKKXUop4fQCB3UNF
GPHyILnBcG5OLRbG3sMmKHVkXlHmjWbvqm8IRyaCWpaqNgcXdclIBmEmi9qaqvCxrzubK13cbi4z
HqrDBu6WAB55QpH+fynMgsAHr8HfGsKAPVXwZo9H6zuAuKLD2kTF3RqTZHBsknhKRHKAg4Yab8ra
EJP7uzeTbscvCVDTw4m8kQjwEXMWAlEisftGxz4bzoj+K88ctEEkanMl1LHLPsX1v5FNLBxIJzFb
Ov+WIncihFWO2acNuv/hPn28lPrbxGXFH3gLU7ZU2BkPdt3rE6nxWwjAkLY62fyM5aMtuh47LEs1
BpVLULGw7pVbspee/LRHoh2aue4/C13SenP/SfrguuVnAQHX7zRzNhps1QqFKWdSDTK66gw+50xH
ZgNysTPovVAisbNuSkoBF5OtlpVdB79/uV0Wc/LfYKZc/IX481eNhi7CnFZG/0WniYdRHrNkoAfi
eypKz1THsVFF28RR3IbL+B0NCBc56Xw8HW81X7BQ/XHWATNuvW4ZHba6dnjlzJoBB1F/majoNuL9
BpvQH3GqCHioU34nzOz/2acwVfDx0hohz1rX0bdez5pk3XhciLjeFsfuth3SFbF4wbPoKcoSY9XF
dh+zEImGHIf5xOZxAg21nKhU/4Bze2Y8hjmT1HYlczA67C4cDp6V7p2ZS5f+pzNW64RbRUjqxV8r
SsqZUjEt9buRDZeyQ/7h8GKltq4W1eAlSYvAozWZ2FN1eok9VzI//TeNx57g5xtH3yfxBelMF+n1
8Bl2Nj7/pSJ+jqZL6GllbXGSBuwOig2U06bPGYCirV1IkD0qmzjs5r1PdLbgbe6NPsrndTABezKV
O83M3qNAIYHb5tftBW89Gd4MkyMqq9Ls9HYWekSevRWj/8RAmb/pTifVLCnfQceLVC6NzzaOf6mn
3zYfMmx+Ttuxrsqb7r+jBCXlO+taz+tI9m0AK3a2s2ods0P9RZRFK387PvlnQ3KjQKc7BLSIU09i
iEYt6L1YJ6SEoFWISPCSxj3eJAffXBQ/aTZKOTafMTlbUUH6phuTtvRHujGCKjbC1hHaYCpTWI0m
PQYT0V5rhtwKIastTaok2XOr9Kn8xXuZwEKq5zaFlmX5npBRAKBnHEAeX93X0nDoBi8hHc58T+bx
SmA07Re1Lr/EstXd02ABU7I3qXXFpljdINFC59VX3sErJn4XGpOq1RFcIqYYeHaCzdE0KxaZB1Oa
q2WXTW0W7ZbeQt9qfdj8+PZIEHi0c8wkJNQ2AZh78oLF08LUvafS8B6XFPK0MqwNiMmi0+alvR0b
UJpAxZlcM9+csbUJ+zB/OEySptPOxBpSfYFIfHIf2E3snC3KeyL1NBNSwroAB2+s5MMs7gu4zhsZ
qdzbfBxmM8ibCxQozrjFmqtM8yk1A+wHlK9/sUJmwRR4swLCpVqrbb9nerpa/TyauWM5ib/XPt2Z
YP0XD+P7xpyDByzsOuA8s2rlIKkmBNUuRIaMSGQISVmUtp0Z8SxV8C/Q7o7PMsk9PUBZNvcFwSNb
Q7KBYjBEuDnLYMjMwF2LrbyzxXAnUSu2pulyJBhIoUeBwNNU+ZfFC3DdFeJXCWuglxJ2h08XTodw
Q/gDkwDnM+S2yHjz+4jtJcbtrFYtOBJgW3WTqRZT9cwr5YR/jGd2xeNcHgEa2EuLp6G7q6sWlO2i
Cu5J0VqS0sOP5VMBQdPp+sPO/Xe6CmlJ67QSVxaLi74V67HR7Bwn/ZKuHufSjzo7yKI3FP/UbCAv
KRmclXSm920wWCKwImSlh0IFYdm1el8Y0xTbkew+Z7Tlv30W12SAxEVF4iEvvqA1WDM7+MQ49SGB
ta4DwqPCDF9BQvdYQNLGfWvFphQvg/7gYPwDFYa2TEQjsZfyuprsSmqtxa0C4y8mSJXVDedrUltK
lsMZChw+mJ5PYACfUg9glWYPGQRZhbSu/2kRAIEpgtE7J3T+zRgAqCbrdEubGRqPLkMxPBuHPSfA
y6Vju0hBe1plLNztJ4ldrskSZfhdN/DzQMULxodfEidoDuxiQG7lv6/m2qYKKC+256e6WeFswQ4/
mWMGKUXykt+DRdUb9rznr/pwAHEY/CMyQEMFFCJVHDU48aooEXuIKPIQ1M838RY9xo1C5MzHvJfY
4bn3ISqPAw6UBqLqRsXeUMwvKav4nPzJ3Crl7gEvwPp9e0jYZPoYo3XLhfmaDVKgryfd496t50st
ae63Brk5HwHa5dGkIAYqEhpoadU+OMEyMcdV+cX0U9dPJv5u3ZseLPO1xwaGdDm3TpvctnRirEKJ
S9CwlO7qyiYpoZ8+cWVLbFFMomqxq8HHNngaC5MkP08kNs8YdPZwo9BggHuz2RVhZd7t2H5XVtUk
/Z4nsicgwzc4f2jhs69lWbFK6GB/Hcpurvt1B8fJxnWtSVrI37GrSB6/+2PpYsno+nTzQOIHGI4I
vjk+QcO5WRojXO7naYnHP8UOHNtRI+hsXFHdvEH2eiim4LH/MmepARu29NESposf5mA/i5CJ4XuJ
8b+PVxo9eHvXGURBZ/zMq738+IXl9F8Nw8OKIagFYAKwH3N+eQ9hOC/gdYQ72sIZkjXCGRFnAk96
RhbCCY+BtQk5Fc334Y/cOC0SGiFgX/+s9m1cfKL3OsB15PVp3gEpEV2ajpSLg+V08tfBKaSyAXeK
3xYQXev0WVSJ52fDyQjVXTn9UH9M/hlGaYoXHgHCOHL5wKqx5RruISA4EmrRstseLZ4nkDDiDcVJ
jOYcs9siQZINeBl8c+JcktZwBbfdEB7eAXzuul6QRt3Fb/QUADFS/fCRqx7PMs8kfGpcT9C+S6DX
QpLQfKpJO46xcNm+8X9SZkYCrACd6np/l9Iui3xlKRuy+bqVVR/KHob5K7e5Hfy/TXAGK4kyS3Oo
q73m7IklOi6+pM3DcI0pz+xe1JwO/NtjDdeB3IVES+/AyJa4yaW0d/gPmIubxp9pPP/UIzatTNKT
eJSD72iEAX4sOlajC4fBv8NtdbKt5UO1f6eN3jBMr9K4srwLpWoHpHs55YRwXrEpEt0E7ntjfZ+J
WF3ehPHKWcp/Gi8Sv5bM6spmr9Cjmv7HnbmTwl/YIWd9Uq95BmUqeXrhszd14Ab08xBFDyY+BxgB
n0T/iTpeGIIA5EO9QvH6Jr2If8QlTAYSky+sBjgG+XB483aIBPlL2/xABO5xW9zU+dqSeWKoheSM
lzYQSEQtQvZ+vArXBjYvbfrsBvxrXW4zgduU5l8HZ/5thvmL+zb8GyXfS7/q4qDS41+vVA9cN0C/
fJQ8Kpxyltz7uPl6Nn1NE8xu2GhOWR6HgpckFzr/gABphNlulKq1Rk7oG9BnbFep1Ptm9dq7bykZ
yi2AFny49YrnwmX9ZMSoy6k3HI3u0bVvnCAz3XGf79VpikSu2DzYb4PNT4CU5PQ4bGlbw8W3ZvAl
Bq3ujQ7yAcezdoF7KEXvGmh2jzvNW3n4LFrIQeOk5IH18UqHbUhBWsYzLtbMURSB2h0JCyCWdfuA
WNsryjaBiYO20d95/4kbB78vi63iFf1r0q2jmlIYJRDibaCfrsC8kn/F/wGx8zmP/SXlsD+xcOWP
uod8Vd+AB1BUBGxhofK1FBoQ8pkYZjOedaxH/UffG+xWJ/pPOhhUmXuInlrYlHRBtAeVPkWZpnzB
kW9Vs4M/0TV2NZ3LLLkparWmtpPmkHjJw2GZHiF5F+mZGKeZWEmwEUVKdvF20T2mDvo2OvOjj5pj
QynodwnM8G9Acw5lKNmm9HNN7R3dK0bkLKp7mC/U8jW0F05hGXLIrNfF1Wg9LE/smczYbp/okd1i
jsl71Bp43w+yZBeSW7kTPvvsIoaEQFIfWN27esXLRkr6YAusRs2QSZllwGgBP7jfGYZzvkdIFege
NnoMUxXSNvlShPbiinoQuFzhoilvvDyR+rcxxNZfY4eDU0fkyPfJvg6gJRi47Mays5W+NxeSdmLk
jGvzvSlnuWpMDUpYhE65WCF1SURXZ1zbLFRiYUuV10xWefNj9fYHmOeAtbGv1dt5q6pmbk1UjhLV
eHHHVv334T5tTaEDpOc//rAvDjBd412nmDz1P7/kkn/XyRMdtNX2lXtepEslm9GcgyRiCbBqNTth
nVFiArYQccvJwFKTQ4ThDeEf1AUq+WwS61Oec4aEyU1x6t+JwnDcAGZu0Qsu3CDCH37w1CG3b8Fg
VMVGiYrUIdWTINTcA+vfLhHZZjgt4D3qmPPRrlKTatK/v+OcUlCqi/M2T7xo+M3CX7u5QZVUO9YQ
6HOf6FBSXSZBT2Vm1r9Rc3YaeM3Lbb/ZBC7yBsMjvXMOTnM9Tc7usWUPJ/CssPIEaLn+60wDQlBj
WoVLy0tGSCgK8lImfVNsgSagfKz6CWo+VSUikM0yQ7vPfKtb7cKqDK9lcj48KiK89Hkn70LJmXS9
kBNJmsxkhR/m/9pv9dHlWPnj6Py4A0c6giYaiWAczSevY2eJcoqBiRMv7DOGJxOWEQuG6NS8GPux
Zsp7KiF9vaGe/6MxWgyuSoFtZZFcqpokv/PzYZyaDEBAlF2T096J/WeGRm4AkpJx0RTpfOi93e0t
60Zo4c0QZkFD6/vmqv0m3b+5Ene9KGO4m+0SHR0YPJumgBMXQgNHFNOGejrpNRAvWIfPiBo4DABj
kX68A6LXbTHYedAt8vLgfSVLqvMfhLqGiHmnK6vjgUaNfZve4a2zrhN+to28ApA6BmmwsEHMvKs8
J3/sNiJjp/zPuYX5b41aBvtH8FMBzHGbz6xxFcKQUzMwg8maXanVQtd4mI7IShn9Ms86c6ye92ax
DtvbJLWc55X/+kJkTOO0gq1XdR/jAeMeYRDhk5NZlqOzo9hwE4bf8iOQpf76uhgphjk5E/+LUILu
mUdrNcOnrxyBCvy4bgpQClvXnq+5zhCLsuUbUZKhaoQnkFCtvTWoVu0y+MXEqpv+zfC1tDkbtv9K
CGDTl2QrtaVXpNBd83k+TAMDbuMPlGtXzpcOAwuF4juu6KqQDluPKv3+7M2fJqA6KTmok6iBQWaa
QBQ78fwRBJtLbrgrtBhfQQroRiz9AAa1A2WdVEVsGUno8vxlPvvRg04kAzznuUAimya8TpWZGu8l
O2Cx6KWmU+zNddDKVt15yj68dcSydMNdHEBDlG4/dqddZDAi4wS1iPE6ExXoRHMejtLaH094j8Xh
vlYjq4Zxf6AnMj8KnTJym2FFOFm/1a9uv4ahz7PgGJe0JKOG4vZUHAazb4BCDovE3oJePR1Ce2ft
KUqkmNGckigFPBejOFjoTw7XFO2PLGYY+v11ewLUt4yr8yRj6bQeGd1N5NlEVsFOYK/LJ7uRBtjH
e4tFvba50KmOuq2UKbNs6xpSAYRL1S/qyzLRkB81jqKXD/8b5VtIYUlfsTIfBL7mYoXp7UTvzMbq
TQbXziZgBSPqYFM8SR0lyQgXoVAq1jL0mK3qMJNj7E6SQrRMgzmHNe4slsuHmyW0Eb5aSwToOq1R
3r9dQO0SOaw9i4YFNe83L5iijfE1kP7Tis38iEPaMe4d/vmh4epDdyoAsuISiMMUuTl/8s1tfjot
g8lM34mrZd+ovEN650ClMp1+G8U2MVIVnwf2yZSaorSpzjh25SfQOWwm3CnihpdyAY7mcnmy0QM/
IBhwSut74L5qnCGfmG1AknT8Bqsu86sWD3vAtcK5h65HbRft3YUF7yhzyDbkw1jDt9cDOoBkLSCX
j1ELwQPnJTa1yu1nzCrnOilVuIQ6iJ2SbsL3cLDtJk9OOhhLtjLW99GZmKj/D0OnQdZKb60GQ8cb
yVnWsobv8nQC6rubMqW1Qwuxp8OjUDCiEkB7/Uwp/+frb+ZBHdhYzicEQIA82azZY3/ZXxSlh7nG
QEtBKL/PXWzwOniAiU9SeHwpbaZMDs2e63n5T7un/XBk76eYimJ7eD3M7xIyRul+LUTx5l846x8O
ZgSKubXORlYXs0sqFC/VQ0TBkJNsvG9wiTGzbsKJSoBtRIqEWgzzztYqAbqTa6gfgLpgO/xrQZEn
QBGEeohakNrWXR/sqhdDxDwjXqaPbVudIaifEQw9byCGxsxqkHxI+VdBB6GQ1Akhl3Xi0VEFpJgO
tz/Z0TSt+IBdxJ1oVFhnnOXPv3SHMiYgrm26Ih/oKfMqq8QyzyMHsyaR1XlqQczvh47ZmFfTOIix
L+BlqGRV26G9bx+bZP3wjV5Bbl8k6pROdf5qahF0LJfVCNnfA+oKAIVx5BfkkvIFDWMzVF10O6J3
py5rGAJlsQecaSqTNnJ6PO1S7qm5my1n/gj+26bKp7jJJJ/m70V/0j4HHl3u6lW1+Oh8TEC9ACea
LGBvzuxphg168NHtOIbC9Qh6x3u0v4yIkW6ItpZRAHopZLnElvITdeZ4LMwmKSerzhwm+ahUnP2g
BYxKJLqvPJ+x+lIsCKrgoiuUBypCnXO0VUH4/ct7byj0M7u84mcHhYtEususuzssJxWWH4kf8Qjn
qxvGTHarBzD8EtldSvlWDkM4ebcQ+TigEzN+pZspgKPO6iYvBl9zNtNeMhEWv8jwMQdZkYWDgo2j
gogJVSS9A986G73rvL5lif6XsPksuaXHEgoX+haTkyPofLZs6bW/+6kgakA2/AhN/oPFYX/ZD4YT
dCdPqGx5VqKY1erEWQmFzHgbcTUV0C1oUUqv0IbAU+EBQXAeJBK5JrJzR7e+WN/liquMtAJwoczD
atV2bLdjlhHpL4fJCs6vK7LM0xnBO/rDdsZhPPw3liCFZ1cpa1Bi47ikSANCZFCUsR8MLwkZZO42
NDdXxyBLW+Xy8BIhRK0iQMtzyHzuFIPXEIEZzqYRH4N/8gfmAXAZJf7WgabzAK++6UbdTK5Rt54M
aOHHVyScw8UDp0PFb1S2uQVAy7O6Zni8jThfXDtIKQ4VsJJXLEC/P8grUICtPUIDmOddK6sI2wOf
RkADVWnokWfe5hILX6V9lBPKhgGvgl4OWGBzWQXOuDwGur5Ca3iUEJn40ONFmorLkoWNKgcg5uB1
lgXVvJp4x3bRkHRXL5l8P2jqDSpE8Aqt1XIkQ678dV2yxTVWmhWSQTc4oK6ajnUmwCTRcoGcWkCa
bllLi66WFAIK3XvBLSJ5L3T1DCIG4R+w8vF8QVg3gdbhPalOTvyhpIXPx3zfHAlgjX+0cXZnFpH3
VAt3v2HxD3h5/SkOvBQe0LEShoWRagu7gtiQ986EuU0q/1m90lMYPYOmft4uY5NTgRBpDFZ1+vwX
nPK9JUsCKdA5egTthXLyMuvSE2iew0CAqnOUj2wrbDBGLL0nf4YUHXqsp06HrDSJxADZ4JNPAsd0
qKCvk8SbIjJcdpRWg8thhrPsmnskWOGKgZl2PUfQpIvrvjDjAt6+m7digzDRAFx+s2XP6/VeKRdl
SFnywKpZ6gRKBK+U4NBF2phImf57V3WFVUGq7f2O5r2klYM7izgH0gdNJDtQ0gR4XfkakCajzL42
a/AOelDX0g3MYkPOZF0vB5hEDMJJBT9p2eGZa0tD2jEVOMsvbHOKZH0NLMXLi4Jh8QH+9pqfA623
NZj1hYYfzBQ4vy1bZjDN2DiYXZLx3vPRKnbWQ/YwHhIxW/D6gkeyJQrr6WDV9Wy7F3xNNrFlTSX6
vEwV4K5kuiZE6ndBI62PGzGrQdenatOiX3iUMWJoXqznOeH7znYH8TUUq16QoJr1OQmM09eCAzAF
1jeKrx0oAJ7NBMBUPvBZear3F4wCsBY6j6NGrWwE8oIjjqbnSOhBxbPKFfjdNsfElVhTQfrcdtnW
xLVGI5IA9htR8TWPnj9Uj3jU3+mKyDyfWRdqOWyh6RZnlmhEoKZRp+42ySPV2MJruFlFtvKTwLFN
NCCKa62q3tWirqFIRx3i5IhPIEbXgsflb9A0pz0APO4av9TP4w9zYsWI3uDe8kUcNoAOBZxQEQNy
xSeWVsEf9u0euGioe7U8Vi8C/hpLG5AIUt0WepJTNj4vLoJ2OouEw2NasSwJT8EDGwHDIgwnMWPV
hTVeGjlxXJrESuU66aTAIRYbL1OAg4ryabEl1vZ9tVd1P4yRpyREA+TSHcWfk9Wca4NcMkY/rfX1
ZBejp4eCdO5JDZypxztLosdCyc7sCjZhG4g6QZJyAhwSdzYagw4EQ/Wk6nI3kmT8oh6y4IHliYdW
+nKWro/GO4UQzY3hOHJzS9IPJOuNHT0bgmyAri07dMNVRedcsF0PBasEz/FBxovCnm/3v7m98ct5
RwNYhkVjvPPWDGiUF7FjTCnRTlU7V++D286xkNj/yxyPTxWL1DB0JZKOoq3bStLFm9QV/z9HvtvB
HoeX6xB/DagFRWJu3KCyo65GjgyO8naYZ+PeLT2TcmFvrCDsjZ6W/aQP7V9zhSiVxWL88EOZhBAf
4D86e8MSVOZMlgYoeMh0Xetb+q872mx+9FGc0tVanw3OGD8w+hrd0Xq+oXNskwKD/8gpmxBNgY5+
7YnTmGm4xxwJVXfraMrEapfEomIt5SZCvztAajujHXVldm5tQklkuJIBjt7bjeS75pZDDlA33f9x
5NOr67xdUZrArZL9S2lGJ9ibUDy1dw2uHkh7sqTnezUJgHIW92hDbkKVTeDBx9L8+R/KKXq9Hz0o
y1JAcJ+snJ9s0GD4W+2ot6Dba7D4krfaP2N2qBQh47Yez0Nv8oLDUhb5j2jDWS677kYIx8456mZX
NNg8wbSJYumMQKHresHjGJxm3d6+uZMqMsGPQIsRSKu2TlHEWgeNENH4qW9GjyKvlv47ZYlh6Ck7
TIZG72cdNDjvLKO7RojG6cc8yVB5wjb/pnaw59zA5YBW5rvDgRPYNJrYr+Qr3gaHufjnsUAZ7Mfs
22IDB8qViMYtIqO9g1d/eV8Meo++lWP0Cn6IGzWgqEkSGVm2/R6YrNhq3ZouNAQItIdevXVJZNrP
MN3stLV2jLC8zYMHqv2i4q+se2iyztDj4f2Ki4VC+mZHngOaetY1p+j0AHKXO4xJ9RBGKYYJwD1s
F+ysvywNIctwwnLKE1HLMGFJflk3GSsqck99ECTRrgXDEpktERg+93hKfFnD1RkEKdRS1J6LaHkl
LqmBTT4rFh8ar5W+bYzt96kfaWPXQPjLoO2WRi2BcT+dWx029bJlHTQjWFi1f5z976n6hF2wD3+8
oexIXn9Eq8lLwPaitI2peBsD0kVb9YFvNphdFORbSXiJujWNvlayPOKRHyPd49kjX86Vn2lkdtGg
XMI375O5ENrOvsovQpLgF2IV4kvTR6W37tQxxD5pFCFnEVpTbZWh4FZncjLyqXTpupauAyrWaEER
Lw7dTKnTk0/U3RXanGy+oNKzo4Qb8dDIJ2buHfCiscu0pB49cGhJRUYKaEzvEpiv7wmCa+tloIYn
AD4qvpqs/cwIHYVPG4DuwZ5MIYykr8d4oFor1jmM2QwPdOtfE/ROyDGbMpuDg5KH3AkXR8uq4Dwc
EbbV+oQSk7wXKAwfiV6FBJYIItROH7Ts7TqUoeC+JlClyT7icFsZhW2ZqoP+MSwoTn9n2k11VXnR
i0Q0/aFrHOdNnhZrz0fJ0edn5JfWcEDRN/JpTi+LYlIkz9agr3xbk4XfFzRP7P4x05kOnqUiB2Ow
fWCL26RCwRNmdnU+eJVXGpS8R3jlHlVg+H70SlLfAtRNjVSVwnP2nyoZciwWwfzfwz1dWUlmJZGT
xVGLqDvqrp7AfZS+Ni0t0/2TSbpHbzMog0aJRiyKxzJAMjU3D8sQR9FIm6/+R4UI8coB91lP+DFT
Go778btUDG6G6mlBx6XFSfqjH/98XTbu5cdIV8X0VarPWg6aRKMMg3UG7Z0P/NzHR0HUEog1Eruc
yOkSCc0C02qNtCfK3+31aIICeLZfj/CqTmxG7yw9VuD+V9fLoc0wCYUrmcJkoI/xS0U/WBVivEZ7
jNXlKnYF+CVgxG1da5zGo2mCodreKD8dc5OX9/WsehUUjp2vX4uui7ca6IY+3jiXH2rtHrBias1x
VXkpEmWZcYlUi8Gx6Fj5IfNwkF0NOGJOB8VwaQ9izILiZVk1q+k1krK36Hvz8PvNe5X0YQpdskur
qUKzptdHcu90kSZevSVYxF2pzstIoJjgN4NvgCusdwwHoHlTQpH/6jEiDmJbZFwEnh6p7FGzuajS
bhee54SAb7Taw/Of/lZrVa9Tii4QvMXuI3qsXmuoommW9fcfIaFkcaBZpDRxv/ELVc8PzmgP71oy
Daz23LKQyYEZIamV01SpD8iU40abt2WfZpWtKQ+1Fpg2gdf+iCMw0bHkDenw37rwEF7+Qb4qZptC
GmrRGBkZJkv/kR1/yU4DzZxMYZ5n1SC6DV+P4vq8k+kQVQ15X+rhn8EwvRCT4nNSRBes3IAbKF/i
P5CGHGK2K08vTq486J/t/7K6EYLYmUqkQJgPIpcOvSdrElIXkaz7Nmmpu7pqv2GLTvLPqn8sJe0Z
Gz7IiUfGJhukkvLBbf3rFUyrwvHLG4bgtlMi5C0Wt5VmkHP17fMyUa6ljACJU2FipoEU2HRYRO6C
sxClyJonTACbc/BKXx6UkbAUuJp33cWucIW1qmn2TxIXmUKD0PRd25tgBK9HtQJ94g+XHjNvBYbQ
ynGdZjcKGYEIQF8vWFa4pUUQEOqksZRzTeSW2PFrwW7QQmQB3Wv0DwRNlunzAMQi+w1iw47pliV3
VCHDDzuIY/bHLWzYG80jsQ2c5UGZAo8zNdKaO+KKpB0fXzZKesEGqv75gvyYo0fxB9VHKK/tHDRy
B4yZXqBLVy44JovWLWqTu5xam9sIH+fQk+qt+S4vZEsZFsP3GLFZNT5h16r+Ab7sTJCLVuk+zFjH
gTnXaaQISbgSs/AWeS5uxOLPleWOuPYUf3uTcDaTmFm5N8/5UqyiJHlcG8JHHLZ8+MblSIaCM9YX
4SX9dDOhkMblSed8tz1v86Gs+tv00fcBpCPRuxUFL5QZuNpeg0v9AP9MQmSeDcAJwQnC/kMUzQu8
LMUcv+wijfsJ/gwcZQSy5Cj0gEjOyU9tfTNSHSWbLdgFmGbHIpNATM1Bp81BmMXIwN8gwqNRIohf
aOcblMADwqnzmHbQh1k9kqYxF8ym6bnmFuYGh8VwQse/fWZLqCa7doQA7gJxlznXG7GXyfrqdX4K
/OQpuWtAOXagN4z99J+sTeBkhx0ZR6x+mWwdt+6EeDp1v64S5fmkYD0wAI5K7Ekl8eRhJmp88xdj
v1n8eO7d7Q59Y5lOLCxBW/15ZLVCgFQzT67D9W+xeON9d/RC2N6DXGv+yd75AgwplWq6HRtSrmLW
4J7tLWb08QJPlRCCQQdN1dXG87T7hzULldVG0ifrkNqpgSy3bnncoT7edfs8XZX8ZhnSxH6woQtI
1UUth3gXovXHHgAzMH2o9NnWH0fj428RDCvNe73dsODwP3WGaDjke488FfS09NvNhcHkPl0DN7iY
VBXlueKiE8mJ/9itIdEgelOP3u8kjN7y75OPptcqR8VCSy3ONxpWXhZJx3jAGliyyB1w/f84yM0O
VJdRkATPFuAh9QPYpe7Pgzyw4xde1STZJ5MhW4YwBzGwgB0ZYy4pJpqvfk56DbhPAjUNI7DV0xJw
+6LQANPeG1POGyQ+d8odj9R9tYFbvT1KtgRFICTDubfv6kriuXS8Y3ckPTvPPXw/w3zZWiEpQWZF
YD1eR7oWI27VWBfpjY5JFX49Nam7NDik49P8tZGpkFbZLePezxSpmua5Vk26vYlPNNjoV/SAOCh0
AKCub39lz9Xa8VFH/nDLOOOwGdQSHLRcC5vWwX9wbLAiZSU8DTH9Ljoyf6ORD5JWRcvZUdt1elU0
izaZx5RIZJGHP9Oyo73wLxi845WMYB7KeiQXLZ93Qfmo1QmglLddqaYQIfNLlRjN+biAUMVw0TJC
MbP1lZjQPoWYHku5AgIcLS3dWftXs6GwvcBYsjI1fb36G4jYMz8bNa2lsCZGNU9q9xl+5WMRL1dO
Imbk16eMLnG9AkxuUOpmjGG+dBYGbeMee32fj1D0Scx0YN3n8cisfQ0DfY5az4q04YS0YsNFMwXw
BtTnoKeILXq/xkBWAo6CbQL5SLU1jrtGFlZMw1V6vAWMBHy82MTcXoU24HIfOd9bULvGGvDAvNws
ej5RpQr9UCTbTKUUd8Lgvnjw7f9o/NacDxqgqKlhaZ7zAC66iCBbNW5In5HLvwQ21zdY5NQVPcvS
yGdGJ5+tKkF8RpVbHPaz3KTIFAlii9rP7mNIWyR1JZErDcc4CpouHktQuEnLX+qvz2ipNjnMzhqf
fqAHqHg8Fj0DTBrnH7iwvnxTY4chEUnYhwqpePw8spvHw0x5hi7g5RFTUnqsj/13Eb56QF8o3HON
waDDU2QzF39oOO5jeqH9itnymxatsVFX/DovDkDVw42mv0MbYwxJbr94+gVzkTssxoM8wfNGqiUy
Hvfgvksaa+/7nmGc8pwb6v56rN6sKRyObso0Pb7PVNkUUOntR5oaMCBRuDIUyzu5unIkpm2Pjiph
eCmogEi48iKTSoshz3BDHlScc5sN3s2MixPf97SkbOAYsXcu+NhemvNI+htozWlsxdm+a6l2YI8O
eEWkIhq+vJY5Xxofm3HWVyO6JWtD1rjmG7PsUrHrrv8RboFOznwAOLUgoQvKUBR0A/oZYv6qpPb7
IE7lWZuiHbZCj5fZOU4eegxu1grmRIGr9hxQOZ6MVhQDIjt5ceo0V/vL+UrJ6ZlZgWcorN7kqJt6
41xUoiSQQZHewf6mPwlsXlx+PDrI2GhJCvar+Z3kPsH4TXYZrRLPUQ37OOQ2R8+CjVbn7W2yAYO4
5rRGAPSaiY+6/U1LFKdp/UlstVdMUZF586OMGzSDxEIqjrDaXl9jP5Npi3DVdpcj4xfto29jqGUi
2AYVMq2tD1aVvioDFwUPwsFZaJU+3h9ONZhtMZKAKPrl0hf2CSITxqZuVmWb0EE8CU52wdZR2FHS
1T/GyStPXhNZRGxQG8KlreV/HHWtHjsQ85tdXBWwiwagUWP+jcYcUjUuaxwYpC/eiZegWEahZka7
LjImvOYnao73JLpwuwYpOOw9zjwjpRhHX6MrANqR34ig/pbJus1yvgUA9dH6jBfiST76pZFZRYAN
sS7hTtho7avz9C1qRtmOsKCoujpaBUV7E9ir8GiTXmLktet+iHiQ2maHsIHEoVR2a58h3chRAARs
guM1rkwHFJSHmU737/xnZu3SmTfFMgOco2wDsHDPNW+tzfxXdwzCcUY6ZxEzngoY2igYXUKPo6RG
AUGV9+PucNBhFycVzj4MmazB7FtGZyoSSBCpQ6r5BP9O1OcUkbw7v7wCYL2rmEcLHCvZo3PhK4fj
nSGwrdUTA71vtBCel+WqXulmJWM6KPEcthdvE3JWiz4hF2LmmJUB+kQPQVYdcj3higCKccS/bRAY
iNbGZK1O+kMo/cAfd+4e798fra3KkacPdiGkmvptsMiTA3A3lGOOa/vYPFQMa1BNnPSCVHDUhoTv
awdRbahhjhj3U8tPTaHqfte8cpi6mpmOp3Mn4m/pnXv+pVjpGE7SAD3NW1GOQdx3OpHEd9tuBnL8
akqGWYCDF+mHoyFdZv1n9lXNwkYvwvwLT69iX/t/M5jjaw37xDeb9wH6yR36jdCfVYcYCJrnd32p
H+RH5Xo/IG2VM27yFnqTKoFw3E1h35V7yIi0pAdjQeAOzzXA3LLvFf3XY4e2TOyzXeSkAT7Rv4js
dy8l5RXLLthqoR1tEoXpDaDStD27qJPI1ro+prHUR9qHNVbtFZcbBcJmqFb89d9vvbNKcFmRGslq
vozP/kzdFE3y0fSe/pEy/k0YUrn4t4qB5V4P7/1AlW7Rk16jtX7CALu886tOLZ4lJWCZXxOhdO2+
V89QchbZAn9ce4IBsbhYov/xsNn+lUtqR/1A/3ubFBRrfL3XoZlbHiY+dBqaOlkPEQNjYBLaXFsa
psECqfFVAXCZjHSMY6+rGU3ntoMI80whBkHA4Hby0jo3zObRt0hncMTNBe5WHSc+8iQoHbWE7FAl
J6r0I+joodGaRqCijzYjKjzNPNsCrRDO+lG2tfXiU/2pUAHmouozfxN/OUveLfCz1cFMYbVWWvKN
+PTJ9U0yFU0M0Xhq7UX8noYSmDDWsWdF/MfJ6nRkc3VgFqEjv1XCg2n71NDEEGxgxDbLQKTuJ5VE
1tzWXbpFwd3Pa13BZDrFLMHNEjj13E2qC/absa44TBnU7thL7UkHtdNrK8XJ0GNgEVy6IuPVUPhL
v8TA00+5PFxRbNzLYgqwjsJaYQl/MddV4hCEMyERPYcVanQmtN0rTbmltu9cuGx1wG3FjDeqcUsE
x1kRoOAIstyw50JTD2SgwOTZSpED9Oq6GLq5gdlu6D4tCBGpZMGdDXFcRUkDbbsVJCuQdM9jLFef
UpP7t2cL2PsOpD1HZp0AQ6G6HHXATzjzhTV1uN3sP5h5FWVJqCIWcuircHZoyMSwHybpua6Dw8ta
vicO5F5nO9QuDi6q+PTKjrb9ilN1ihV3P1/fgxDyjXqIe3gCyHt/95W/f06TokFKIJb8+Q1fs3FL
uFWzr438X7hjo2omPM+T9WkJJxMXXLyyLtVvpCAVGtyq3LBEDVjSeTa7uBBUr7TzlT1iUc4B6xEW
bfuX3qi52fOITB8WWfkbcIW1q5c0lhaPGR/TNkygh05HEb1FVXHys97x5xG60WRVGecz3zuYk1q9
hQLfm7jd2NA4xqrtG8ig0qggm22p9nF06ePLN0fXCtgSrNdIplI1fe6bnwn55H9WbXQiGQF2A0DP
Mtwy+lr9DD8HDb+v3Szid5hPH/39n4HpcMNmB2Z7QVPiAt+f7FOGtR88BfI2Rl2NG0XfoA1CVg6f
Ne47jM6tLO8Tmdxg1M0D88U8l02Qi53JsFFxSZWzVDs8k0b6b6csYT74MDqhlA6GJUsUdUBakdOG
NFSlNzuZQNDYC9ZZiftgjo44EnH+gkNgsEBgpkNphjowcERA+LkqUd47SaOPlYtIwT4hgE4KaqR6
pDuQZrD4dSk2Vk2vqjjUTrzqTsVkSmJGvgrGLofyXvxILGinmfBa7VCn+c5U5Aod7tcGBykD/tsP
/pxCUmtRXjCAVfm9v4V7uego4k69O75brSz6iNsL7PGtgg2lPRqaynrTgEAwY2WGv/VC7eHjs5u9
uSr2+P5CJ6V/XUb5SOzuK4UOrRPSZ0XBGLm2y4EhVDJeScJI0fHuTPOe+ra1IJEo2swwUmkJUWfk
gMMRqDDUDQqlFyzM5o0YuVzITg0Vnp7e4M+VBMbd6CmjmqpPgTSTgtnDBIOYg8Zw/vsW46p+kTbH
nn0kGBtoWFXNk2x50nk4sLof6NhuCleSJSLtNv0PBvUFRyj3cQdKv7NV2WML7he9w7dDkj/CT3Jl
0H6U6kJ0kTvzMxh9Q+ahFpIqLY0e0aejVKs/4be53B42m48EZ9bRQfu5ESYCxibyBUnwYdS34YGL
UVOuf5TOotYsHQSz/FbxiBMn51RkptMjDhWN2wyPQhoUbimqt2FFDUfY8nHTHbUe4BUyTd//Y1GI
tLQQjPSdPFtZORtcYPg9eXCyWEJKkImqX1Gzywp8+mTILH/KfNoPyHueblyFzE+k1b9LwOnji053
KgczuideKCl4+9bMksnTxURFeCe7q4xFeW73rKSPiZl7bXmkfRNiaYWOgPPn+s0YP+xUgaXVleUA
WHQeHGH3txhGdSauy6WxntYKGoaeiu9jnEyp7EtnPxDRjIJwfo6xlVTDOL75Re7DmfhiOr7ehEpU
XooAqLUk+AvZEusrg5laYojXyIbxBcwVo88wiyEScMRPSOBfk6/UU5ETCthdanRclwAuVlUu24pU
6fFeyOt7PKkyKhgkR+GOfDZAf4neuE1rXBEr3tvGAp4KqeiePgoho2+vhdDfBmw1tKNOUT671Tt3
6z5lFVNd0VQD7bKbPZGOEX8Qs4mAKpgXANDJvWHRILtg1fEbPq5WZwHbGxKAX9oYOWzoBPJBCqqq
NATUT1SDJi2NU231CIdsYpsFPWJcUzQ55kf0zGvYkN5E8IBmXmwSXrQlacfEWMamrQiCXn+CFduu
uxkU8wxCRM8TLssDRAouARpr2o9VAvKTb3JKUFJjaFVHc573dbgQBB4NpcAblxexHHbmHTtutB/d
g9Sdupaf48h7A4nL/9i13GiWiYo2+Sj/BebgL8kyQMlSvMhd+RlEdNbsOj/HWX966EvWtULf5WRt
d1fTHaRRxqrA0/TEVCW7X1Je3M5c1HENMQh6FKa2F0GoTjQn+HR+vbws3ayoRNvC+fV3XkcvdU36
1F5TMQ16VW0Ne8+6gZWKzgA6N3XrW8m3KRlzi2Ovym9kAK1aZXpJBfxyDMEqVxvimrYY3fUle0hh
UAgY6Dd7LhEbnH0W389OszPW2r+O2mFBavCqMbjhfnn4ZWmhZ3wb1GGlHibnsKANGN+uL9BWSdyu
bQ+Ytb2AGEvWqNC7/5p7EzkUkX7k++aAL93wK7T4D3nllDAaveumAORH3AgcULZj+FsMk/SISaSD
QxRTRbOyal6vF930vJ1rQSLUPLHTtFUw90RJtXBr5VkXcCcnKlYh4l+I6/2ILHeTpB6eK2d8WN7v
cKs9hCsXhWTaiNWC/Km8L1s4/jXkr66ApqJW8YUyAhWnrWTRaqFUVqlTtkMS3HXdS44Ww1KLE44m
QDcoYmAaD/YWpaxXozcWnPyvlMDKcTT6wEszZNTXEAT4pHXv+aGppAnCr7yPxeYU6H0HZ+rAeCLf
0FyHx128G9REcfmiYR0xVFR5iADeyE/ssyVzpSM/iXvNsLo6TfCpYt+3reCoXTlBphulPOf3ZIcJ
m3hK4LNuYopwij9Jtlx87AqnS4pZfdaNnOoimVArk8AiUd9/oRbuzUKGqjrr9ZSPyq245k9cthIx
uVDBpspsJAv8xngpKOVDo1RN/b0BtCGgNZAlGi757qKGR4B29vihh1aN4lOURrcMFx53d0/V1DcK
gvZF64QMIoID8MIu8XjrkSv4iRc9G68JeHo0c8naoE+c5gdtkb4Y2PaYgNSpzU8qAZFZBqa1R3Qi
yXYFFhl9Tl8nddakSBLLPgZSx/3xDLlrIt9HqMAyFvyBCKWhXpscam8qWVBTZR9AEnBS5y1k63ed
cbaZYrMwUuzyHRWXb0ZvbtEKjIb7e6jJ71M5zCm7p7Uq+n2xKXsvEI6pMsmdGjx3iyJpzGsSwram
zmNQCz5nGw/tqmhdTAfp1Z3J/31C5cV6mje3G8T00JRjSxGr98LalBxkM9e0/tBtfYVvSeCAqgbj
bfgBpiTuZ0x8VSRQ9JfpCQgrQskKMwEHNNl1E3Gbd4grMQZIvmnJSdKbkrvqtRM2/UNDGTeZqRbF
6CKIEbrV1Cw0RyD/a9NspaB3qkCo1/kez3Yzz1J9VVMxZlvqxlYgWIcxKvvTM8eQjyCoVpatrJim
7AXMPkc8JSLnmZnr0CxoGpcIs/26BoSpSCOFejm3on+kOphco1+ZMk7sAEbnO36BzCZDg3BdVnEH
3GD2RjEUtAsbjlig6BaMr0EDUO6vYAuzlnTHeUJDfP+h/nIMnZScpCokax6pqnS/yorD2+2abDOR
P/h/T+xCYP1TwYX+MIYkjZo2rr2+Jyl546xJwK/Jvp+TccKAywoWlrK8L0n5ZN7BdqTFT7z2Cw8o
xt8YQQSBYaIGSrWPQ3evlolDMrz42BJvSmBOYfLMFSBFv5zmwJIA9QXoz8iwdTJSQcIruEOdNEz4
k3FMmYh5CLc5Jpsc8S7h0wxrBxc3u9GoOXNRi0IS7wwUn2z6A4Bd3FGEX5O3HqH/tTfUxta6pc+W
8PQRn/M2UNH2G40yJzVNMDo4x+TkJPsJ4xh4QWHi4sjYoujzajG2pK3JWKzjWcoU0yxezdXknpgv
hz9wPXddtWegFwxET/SXppbZbR317kEPnK7r+l+diIz/RS68Pau62FdKmN0GouU1s/ODiLtQZnyY
YWoG8NcDbOXqcxNcJH3fswookzpxzqCU/Kl7yPvzFoTaQ71RWDRWKMojwa0idSx2QoAVOE97Je/1
MwoAVTmv4O3YgSQsDXnMkZ5+G+3YAieHbZEHKT+qNLcCqGVXLzG5R1pCVFgH3FyoAO/yF6U5hbuj
bMen8W2LH/49PNXdPMMDdJDXHTycWuFPyI2WupLkO1C4ANpTPbXkyzRsMCcmCpHGRXyHsCC2wh/F
yGRJx5Z9X+yk9pqmlDeMjwRns/Lep4l7pHe8qtb5W9hlIzDD5BmId8QEVOqSTtAmXWPKXoElredu
A5AeiX5I/HzZcRuRo6g70BeBTGFQ+0mEtNAIyIqAdd1GPZfBceLvJkiC+/isdpgBKNzg/FK04cgt
XygG5M3DdQhuCkLIp0byLvhoSuqhVGeOhSoHwr82udBNvQbu4WICUbBvzNJ+yS2N81MMTXuB22cx
3RjJ4EiFMdA4Ni7f57nplQWoQ4ySk9MGIgRv3t9QK8+11P0EhEG7lauv/4T3u90lc9MfOFBW5wc4
65sGrdTTgyj1uSakaJyZ9++5Z+6qvO6hpW1+J5M7l2T7lsGAmZEOhH6hjerZfE2CL0BFSdZH0Esb
xrqpUFHb/SPX07WRpBlBIhnbwjgr3Pl28L1mphyOcKj03CK6o6IDCSPcXWva69OUtkmPPv77oRPg
IDR0B1rZ/SxW5FwHa1kp0Jukua6s5q3isGXyW1WaQQ5uBFWnvALYHaffNNSslxWo5DTZ9ayk96QE
iuYIJu527vZ3Bl9MskwAbWLOFEydmipYwFcEeDaTMEK2jkA/0uJw2O+g80D8+uMOTRh/XYLmTTQh
K7KOzS0jxbOJjFD2cbWe4X2wSYSeh9wDq9gP/i+YItpAU3VXGX2JqOwVE1H+dVYZYoNnoNNNpam8
/nX7U407nvOFApivD5sX+/Qh493JZzxxcFJq5I84OBvchSoLJtnST3UtQfUB3MGn3Mi8irfhnSj6
T0OX7H4b+5YCuqiTfxPPOrfTY/27GxwWPDIBayHtde4XBJjPXDpgXnRE0IQy/RFkUvmAwkwWB6Gs
v0aUANI4lYl/lNugql6e57/wxweHnYK4CWFjmt59P6pdYKrH9qOmJphPP5fzNGcTIxmfVIrMC+/M
iWxwUaoNQT4pBY0+z9CTUcBNQumCpnxrVd9b0UcXyDpgj6b/+AFY+tyj5OR2f0Ae61WVG0IcCFdP
dHdHyMZqgvKAFZ/HLsbaMgIHpQZ4RWnQdr0OYOW1JAYJOnE8Pt11Ul+uV64yU0OwTJkeZ2AIOf64
IGm/cvGnPIx3Cgvgm4LQNycjyZ0E7sdfFKKtAD4zffcBBpaC/PTWhnvvrnuIUF+H2czcJg/A6jK6
TW0++57j5v+JzfcTvAClYs/zq/bVIPbK1v1FMCY82G5PGNTie2ETlh1mH0U7AkCSon3pRFCMbZKc
N52hkS04x7iVSi74L6p+ucOs3wM8mKfJtdOokywcpCyqRoK6Abq1itMJdHBJGcObOo7nb1f+xrrW
Wc/vF6ua7FU7vz+RR0kNm/Su2iW/5Y3b/m49XohylQcNVcpH7Jz2JTsqwPR1zvffvaBo15Grji9o
/Ua7Uo4X9zgOUuP/2vuUAGNExumxBTnpFiccUsFwG4TT3S/Ykt2nWgnmiwJ94M8KjE7ldgg1dPZO
HUUL4e5ugYhVY/hdwr8JEIWU8Sd5N3ZHAJTWQblHBI5aDI9mQKx3+eTx0S2vImvL0zE1RMRdtTvt
ZmAqCBrWfBNrtZbIq0bN7it2sBtEJUZ8P5lta/iuuIv5i0Ioi/LpG6+pTUJQ2eaWXiNvVXW7uV0Y
5jk6OXxIiWaxK1y/q0ba3FXwIpjd9LQYPCBCJiclUgU5RXHXKIF15TBfJAhxgSk3X53+rf7QeIad
6kU9kS7ZaKUxnKMqutqUxcSYvFSF7M/wIGZrQSX8ts8K8Avnj05+0PQXOZqLV8aI5lFL4x8v0fCw
zkazE6wqrbXuPxG0GDGvBwYi9q63Y3twMFWHTdriEj/fkaN1qjVaX4gT4TSAFexgBKuGlqDWaddt
8Wmto7CnWf91VuZvjzZZMQLF+HuDYkU8HlDsr6XduGWMlzp6bLqgnmBvEvP6xfVmejYN9h3RlqMy
+9QLJDkHF+A/0g2rPOMvQzRhyLswXn0b8/DhU6V1xE6hAc9NjdjyYznuZcKhM0ln82HOtf5EWCBF
vcQLiKQPT5o4DUXrv8MFsQgy+5Nm0TE/KaGiFNlb18+W/0QGPRc1tL1dx8RXKJbqR+owvg7OorjP
weIZeFgvYPwUvxqiPGeNQ9iw+Yh4heDRBdqGQMIkQAeRUooxHVOxkZFSnefyjY1kxrHjl7ybdo06
hwznFvnt/3jYZ/YqAx4lse7XBEvALLje5ZrV90go9FVgo00kjs+quW3yS+/vW6bIFTiGwhKve668
YcZVAk9dGQlUDw0acnDex/C0FIaSxVYUO/eaI32QCkoqQg5PK/B02FMNFK3cnIIXIPHKRQi6Nznk
ZsPLAJxF1KwkLkN12OsFfu2pjIMtH2jCXlua7z6Pyo5rjqSE0gkoKs37t1OlYauvZ6XKpjMymPVw
h/Z7jywwGSFR2dfKX4cpUcbIdIWaNIAHNhD5C8OlP7fISIqHJS+aenBvOvSMqasCTUEmKWWpSkgT
efQesdhCCglU19qxy+v40+/tQ72fII4Dk/AY8eeiy1pn96Eb7j4FqmDQSY06+nbHZdTR5OxGYvNh
yUJAecMNRV5VF/8MRkQsKiQVqMPiFYh0xTX5oUwib5NRVYQ2PHgPVqdXvAqsxnkjYfOdCiqWUcxz
0yXTvRFxC9euuAFNfq0Uix3S+Z64kAepDo/GggtUDs9XZbNLmeOl00B42bZ1aKx74GHvCbhdyAgS
ZwqufQPydq323mXRUZxtHDkXq3anE86GPJg9Bukgj5/mAORRF1LT90XYApN7/gcxN1VhSAy0tx+M
ids4GQJ8lC2YjqxiNCN2h+1EnWg+Ogr0ocy9nYq4p5lbrZpGI5pEshjGO3RvDYQfiHNQAbE0Y9Go
qDCvf8bj0aIgDGp+xnrWAluP3zqFAdokz2rk8W0YwJq5qFF+RTqiMnAWOBNCswzBFy/BJBj5ZQFA
u6AHQJ5cDeLQcHlSMBET6nBDv5PKJC3axhQuSRiV41sMhg+8f224jBa7wCojwXOYw9o+LWPD0E2u
KvucxgD/90de0rTF3TWIcQJfZynTMXj1QnNHLTUofvpDIRbC4f7dIVsUhxFH6qTGnKGmAhfGwH43
TYPbDq/ELqJcUQsMckqGKrK6/FsqEuz6jvWpKoeJHRPL6iMEskBgWz2BPhbjl0oss6Az4EccmEEa
yL2vPxPSgeB6ZpqpHEgFj7WRSCdVRQDM/jnONIvHsyxg03HacPxYi7L2YYVsbyrRSl8wEUJpgF+3
caWFYzEmyZzTOz7rLAJZAFH8zdRpxvKKEbbCUqstcC0f5IYvMXj2/NgG9rln8vfjfpzt+Wjyq5Qv
Mesky3x9U7WQJEzej0HIxbjSeg7QFt3LA/IaVn/7nDDb96RoP+x11BNBVniOiUpf+kkhTwcTJtKU
vLsBKNoGCxD4aeFH8bZ7+8ki6EKRu9GFhZnm3Zg2pHHgQ+43sSSN4ayqCKzmY0d9SsgXYFbYDu2p
ZFsXaZVTWYSIRS5S4VT1VAoWxajkOFuopP4N2wdg2QoIEieDbdGGYNyK4G6m70A0o2rRQ41rpBv2
uGFPyIAI8sZrPXNj4LY53gcu3d5kSVH0LRwYcr5pY1eG3mIQ3eidnEpGZmOyNNcLFdWZfRAomGty
J9K+sLnNjiEn7uB3TbTq0MK3LOoo5SKVQZJQZ3FeYGdRv4xKZ0Jq93lnEqDs34w6zDBPy8/z0JzV
arVOv4nuT20q4OWkgnjh1fmgL6fcS7O8PWu0HQSl/XSWP+sdkQyRGpCo8EdwPseRGG4rDPpoc+SM
iD+p9W4hbkHqQFg+mj3NeTjmYALWKfzYxonDrz9tpyJpr4RP5ivoafKfY2gdP+D8DbGNQSgbhbsk
beDXHdzFG8FtcHJohxUzX9ehAbWNXZcnS4zFEMRPGJkkwU5ifDn13YDw/nEC/m0/b+Qbs1wALSsp
w0uqjTt8PSLzTrPVbaDw+nNJv1hbtoAkRh7lMUaG7Ai7nZysyiprzgiYi2Ykm82bGjYG40PMYNjC
rW8LW8TBf74av6B8qoWaOGU8QSlKTIVCRM3aHKV5hTiMNEWZrXZiXyrSWNvMbeQukPaE/S+3VtYQ
b+PqM7lyVIxhW9UUzgnGcSEoQR/FnCaxYH9+IphMGTaaGHT3s4lpeYwQ0zSnH4mInvawt30da1zc
VNrXqCOaFHVvddo9O+CpJucaRidkgDWNVrlOC4hrdkRsDfiYoLlwmlaLUtoSbavg0pgNU+N8x9HA
q7U9aapxbX9mp9+kiNkMWWTKCKDnS9NHeh4E9nsy+ffIB/jQCrjYBWSVK0aMAR8xEXBI1Cz4AJ54
o8P2RPoiRNQyUU/Pw+fNifsEKD7K9iC+wsGMSINOrZ2CBJd67PWZt2FTw9AmgSvpHGhMbxclDxNe
r2ZBhzGuhdt28l9LbrcWbY7ZqWJ+Mfbig5b7CevlUs4gxXhmExr5R/n4zslmEW5+X7Rpa1QWFC7H
hmjCsn4TaYRXs7ciGZdNR/S2qHQ39jDWTjxdCUnMkGcQYi4dD+cY31miP6qFkT7fI+klyFKtjnTb
WSwKN0Nrw2g3eDf8AmLbkWCTOGWx/jMa8Bezm2M2xXgQ2f/qg1JVbL2t4sXpCIo6YzVWzplzhJ6l
Gj2S1SElkIgrewCf7lDui9I5BjeoPdFapifeRal6W9CdydLpRm6c3OyZIy2cHWnOtqzgwrwkVcgh
uog1CB5m+AhO0c3ODrTsTQHeRLlFEJkq1hxwVEt1ZmBhKY1ERc58GRB8W5S2ex8B1dimV/Rl/zQm
Y0Q54tpBViNOblnOd9FVOWZoFv9z4N0LgWPsYrX/tPCc4D+lp5ONIr06h7nSfVeUhFkVRwE1Xxii
2WoP/Snc9CylT1WAfF1NcCeYZZqv15YHzFMFuIaqA7MskfnkGefJZxIUF7TxytZ2iT8MPJ2Ofi+N
1u0cNprodN+AkAwJSCkgUV6pPhgutvQLyOBq74u98lPP+lRg0R8MTQO+nJbErf05jc2qBcRngUsV
VdYqLfsohKqMx3ZYykUNXpIRL0fu6XVOZwimayLnvktDJqSKGI8EjOsk+DSrP43n3sQPZGImbHd4
3Ow1W1w1rm0xtgATARW0vZcHxETKI/XxKCms47FSkh46pyHZdHl5ZbJhDBSBJaMYtWt00cu5zXSC
hVeHazXcr3TqHw29Twp1yGs212Ky5yqiaQCsE6eIvEcaRNli/1tLJSK/T957QiwOwa1VwBDPaXtE
r0LOEaTYWSGfTLibwRRfE7ZoFIL8+x6uTdlGywutbsab17Ak4FAcxNJNRlbJ3hqNCFfTyktFoW0r
q1Pntgd9b6uBPFiwtAU0UpY8gWWMTcmtuifNTWF4bNDcTFYSfUCbsZh/AZFWFvC6ATyXhsXK6hrf
JUWUWZzGc52f4pjrhKaJG1rHfaubQxofTSSc/2FtoqJ/8WJ2i5VsVUqGdV9905CBl096assKB1xj
3EZQ94uCeGhGbMBPWtB/SymgvR2j8SRFkmEJrbkX7ePwCAQfKiqgNgW+mcA1DEqKxxLP314ULvjb
6bOWm+BkeZG8wUYcBZqy3/kogAKBY9QjvN4zY6u/m50hYpUSkd9w9BijZyuxkKr0a9h4VjIVASUz
eAHNvjBgDS+ODgYlqORFHsidFkw+9yGmo+3fY7v2vur/5wpi7eeLoH6OFTd5y6AdhiOpH024n6UY
WsWmqIWGsBSPTnlQnUB+EzChtwHIyFYRity5A/U4cLg79DZTTN3m3ZlrgMqwbbaKfcXcIlEbSMlf
ZPV1esu4AY3aAnWOeJ97zfwYnlDe1GHktY1fm4qIu1qe6vYf3Am9nuZRcDGhRpxDrQ6c0HAtK7qy
UlyMsFdr1YDBVW7Ng09N3zVKiEYjIcbig99n48/OHTgJVdKfuxZkYgpuv3ajlB1hFw5EyLNqiwMG
Ljr35ie/vz0TY3IzZpHxZSON5+I4H88OD9y3TjFPsLx7fAsfn1XrSSPiZ0U/6a7Hihx5g9jlGVLc
5xbjVB7i8AzNo0nVUPvR/e30P05+Hy2/eDTS2Wz0yHhmcGm54Z4YBEiQs7vwl52v2HsUOGF5NrDL
iGETf7RNz2kEQzE0QFZJXr16xjQAF65GL5tMhy0tZte0gVI50szfonDiRe3FfwE7Lsz90zCGK5jU
8GtVANUBrltVTgpajM2di15tDWxUZtwJLq+Ob8gKUMm0ZXfkWAxKCbQoBpedvurVvFQqRYjLYMVI
UkMt0QC2aZmIAHZDlqj1r/12IQL8Grtv0TFHghD4F8MB2icvyn+FAU/qiCiGkU1mjgOxZoFZhvZw
itkfi7ILDcEquhMWlYRju4Qrh8/Sffmbj+ZFZeXwh3EoBcntoNO5B1NfmPV2WQnzTR7v9hg5crx9
SRLFAQ95YPgbkciNStfk8IuvqnHO2IUJbZEJE93xVhwVZsIHSl4YMYj1j/WKOK3ZpwO2zQYEXRCn
kY5uyC40RVNJBz+hqmDalOC0zrRDw9mQ+rqjzFhEtDJLEznAwZgOLR3rD+j1DF4BHVf5V+V8gyvR
E8w925LdovlgscUj/2Vyr236RxOSJtAof25Q6qNzIYU7oCprL/678PYcm6HFxrENuhSpfuhW/leC
Qri+JtxpoLHOuB0fwCA0do6Ag2KOrBu9tJVG9bJBdewfCLr71P22ATnV9xJJ6+g9VRe1xb+qLYgF
/YFJXBzl4sWActw8BfYMKVUlQCzgwDHh5D4/nafwdzdXLQQN+zmO5og78HluB1vqE+NesH6O8mR9
VoMMxapuCEVDL3hFq71KrfZdkUMqyHKJqI4X6bKoAKqFg42WBRkTKpChwlXzMI/2SG+9sbWBgBXe
+KdNLQnSnEF/z/gfaB5ovLK2CTkZEmGvpkCK2d13jcpfcJI3FP2wfkrFYyBxo6gTIAUujy7GBuAG
PX59K787EfniXsrlZWdQ3Mca6FFYTONNxxsL5CUd4eZBF2ZS8EVJAuQU1SiK3edVr2o0y8YgOuv/
SuNdJBfatHqPNWzkJOVYeIO5KlUvHi5a/sUPIGvRreOzvRCEUC9+VffvjlCvaA0HDhDU6+i3Tu5c
8HZ0z01Q7PLB4j+/JjnBL/imfsusUbc2lOC26lxf/HyKiU5ZjdvAxGtDO4S7BITEStIljOvlO3MH
gqqMU3ssFwM8pjjOfpX3haCuH55I0jvE9dMPlC9spHM0/dLS2udrVuKui2fn99ndIvueQp3IGV1o
yfrifWyXtyIZCVooaJanfvT5+B3wWuHuJGpolmPWa1seVWgSje9byX/VvZFO3yZYI3lMAbd5fsT6
e0OwJHvNN4aeb4KlNLtQB48Q/L/HSKG5ciPKlZTmuReHbHaQCr0fG9KuujzCEfhrHFl+22lDCrhB
SMSxXRgBzffgZAChnpMsba6JVOTU2WD/nYR7oUyflpU+n/eD2FnQ/EPs0zjnNGlYPMsj2d9obDk0
uFsKzP/p3qkT49lF4seLiFLCXarYTDnNOfgHhm5qRZxLOmHsl3mL9Y4JMZ28+WTWSmeFSvrI/blB
hoeBI8qk7XY9GAgFKfEDM+tKy44yw7D2rZzTrtY6dkP+cSXWeH4oXdob+D1XQhyl3+E3OjPQHKnJ
+43+nnrtSIQCSdF9+nxx0/OsHEP1Juu3bW0QwlCoyMlDpHuk8DkR5pAhsLiSEcUZZ+QThdh2aIxw
/0ZDMXLkvAtWMzW6c6gpAPZIq0fs4/gj85l9gAjkO1bLvRxTidSVkBKjbgySDkKVc865ZdndIvOs
Y32rq9KiCGwAo8nMMbAEIaSQ/cIla3XXyqiiGjG82FZSh5z65/IRf6frQ4zEfp9O+SRyniWKHgeX
Xy0sMEyhYijH59MJX/XjjzgfXGyWJHbcB4AvfzK03lUGngQ6hkN6nZ+lbakF6hwm78U8cYZiBtgb
Y8dwLX1kI8ktwnQeeG0rCzv9Gsxzbe5LA79p+P51qYwTOZ+CczN9DJkezjc1G27DCdn4oZqVDLQv
THVRPA1U+BxkLDAsVoEbHg4a3fr1QoGxBMP/9mAXsewwVoev3Au1dFtN41qhNV5WvbBupAiqL4Nh
mu8SbUfeEh2dHSoqcV8f+M6EZ/B9L4ozNas4bqc7rJ96kHpuaJ3Kb0YAoykR7q4zUv2Dc2cmR1I8
iEQiXAS4M76yE5iS8R/MIXnowPe6u90DbO+KGriMGjvDAMy8ZnzRcioNLjvlLNjAY26bGK3c4uDL
L0Df6bCI3yXxhamF02mefCceX2YZn48nP8yK5GSydrXbc5UJ1MyF8bJQevcPvni6UeYIXZsKAf5E
E3ECZBIEMkiwQuisy2Jwc0svfWVC79Oy7N9/1WWG3FUiFmc44aspA7p4D2I6FrfLxMFa7lwLnuME
NTc4YhWDZQDHLnRGuApZf0kryddqoZVC6tpe+0HOt1rPFDqw9wXswYU7S4pgSCmZq7+6qUIApHmr
0lSRg7X3JadYdkijdlGss+Dddl/bnFywoFue0dBd3d96Ck7iIY75AdDfUYTpsow2Im01nLngSlaB
3l0ZO5I8gC+diTrjoTmk4YF+dflrF0njYmeLo9W+j4w/E/ZKA2l3GD39gCF7qWjqSrFAIFQaPUo0
PiGOw389MAYmG6ZRakXq0aDWWIuinHY3q5iYZxoUGPgNOBfEdg3ynRMgaBWLsDCaVAPG+rRQktDL
XsBVIFwrlydZq808cZ2wBMxGc17hf6bv012l+oXRI02HGEnlbnwR1HO1y+/xLCBOT9VQBxS8njVF
EAXReVriNXrkhsE4djCKtvoGaEfu4gUIt1v20Rp30m335HqS8Yn7G+dCfTEl7wNms8zP+pluUcEd
b101yCi6ewbI0e9gHQFPeIsrVJlse13ShhfSi0RJVXq8VCdBM/B/Y6eWN8ONXQk+xwB66jwwebdx
DdGn191RHDFRG3pMzGyKrI1+sMYyPiNEzNtO5RJR4ORkr2JnwEHJnNBNadP3xFhscdgi6+drWS7k
aV/jegg7TJfygXmbqDyAtjthdqBE9mszw3gANeb/ZOL6WOnMt9/OdzJ1HeYvBoRvtHlodacGQHIJ
ZYZ+JUcb6w3kgiDWXZI9Se0bdOUi4aVk7j7V+1Enwf2FfshrGH9FWG1ddS6R7ONoLaVCKlT1pDHF
ZZkTgP+JxdEvFE0U9eTDH5r5pVtRts412aK6Zu27hVIRD7SS0fsCF87BdwBbUvOW+bxiqpL0zUoJ
j7th+qrTI8V1nYFRaOsF89IkJ6+bbaTfVxWXuCKgNGbocr9MBZtK55lv6VKKIwBTiRUriwA4mJys
RNIezD2ZwcJG+iZOKtUXhM/pz+BYPHTn/TFFC/YGMsEQVpVACcVPAhHV58VX/s1Oq9jlNMca9U8v
H5yEGvf2+GVIAWHDAheBVt5l4l/M3mvyLtBZz68Y/qT0XMmlRQEz7fgOjaLi0WfOxaynTgiwrvFP
hA2rPOEP4k24Gcpl4ctRzYcYyiPXHnMiUSbfqbZ5YczfTQ2LKkgAgjom4oaIUFf6t8Sk6HPIaoyl
lwEOXrhvv6wyC0TicJ+r5BqWjbjgvfwYW7Su5ya4opA4ZnPkRNLNYXyImOdQafAgn7nb1vrOJZM0
RxXSij2cXawB+4T5WdGfYBWclDyYsXsT2H+bqOo8WPf3xfIy65KG+Qrnmpy01zBc5BCk9kPQG6Z2
h3AK8o2CKb1eZ00BCr9C4p/U3bpLpPePkgxfvjsVaox/Z2VoGc6YhJr1ATpG4VfG4ZJ6xk5Imi4l
pc0yhwyVdHQAXGLIV+QIxCi7gkpNHw2UGE2mRLoGyHn+LVl4H5N4d+4du/SH6ZDVMVW2FqixxBqR
y3cu5/EIGHgdPntFgOdvFODodowQ0kU/QzRyjE6rtErfucEXRtDEB5Ga+cK08jok+zb+KMKu2IU9
ru9GkE0koHwmVWwB8qj2vrWB2kcBUBR4WCFGKIgf1YE4e1Wlp5eos4PCY+Edf6USU4rY1D72QPhy
/3sa/omI7pPdA8eCZsmpbKYNp8XdI6HODEG9XSuxHdougFW4v/mqXi8pxnEhMQjZvs++SxCXE0Cf
nXxBxoFYZvx2Nm9dA9WE7QusuYVmdfzJkN0jwmSrVaEGvxsXTjgmho9SE/qHBTqWEy8DBw/omek6
eev+Z3XHYIlIRTGX1ANVcawa54X4iWjNMICeTB8VMNUtj02k/7Xx501/2ULdbcbni9fFrvEsNiIx
3tTLg+xyaBVSUdG0BYgiC3iqBEqI299aokpXhjHF+AENnkLn5DFclvcOpoGIYDkQXYtX1QHlAY74
2vPuXfDyoEd4+CnNi6yrOHzLxScraJJJy+D/YFbFFqHoyM6xIvE+C/c5aJvi3PbdxMFaOn7fuyrI
ztsXpS6uH7wOwBfCRvAHH4UctJjksZCZ8zs6FPL3EM5/NKo+3lUdHLuRYNjJL7i/5tM3KmLwtbbm
qZE9vrbkEaKhNy1M5E0TIAq6yxR5GMTZpTwZ09BpZ8NK5fsH+O1dgECEN44hhn7KYyT2JQXuE6GO
7FRA/gZYBL+Mutvc8NhRNxjrizTcicv7r/KoQqTMay32arWZCzeKXrZ0ud7nkd71HZ/a3m4yLKm6
CqcvCpyXjWn8UmqqjxcUGhnsREh/+HL8B+Rbzl+hCgl0/mAzdfzO9Vm7ptKg8OrJBZx90b3u78BV
MdzZn8aYe4G6WkZP/uyDzLjYogt4eowTy9J/TlReb4ztXIitK+YwH2BtuksbaNn+chfCDO4O7fju
2QAJH+brPhN6xsIhMdLHsIGqvGEz+od5HNDRc1FUCKW7yjqiI5v736hCP5SJ5BfvrQD9ZFkOE3bT
UG7WNqUWOUk43gwnOIFv8Xd9ZotUXUYuiucx02ffXoKFkd39noHqmSN6uQdvk7EGfj2qsYn3CQ3t
cnBlSQUWL6eo7IiXpTe4HJGURVqgWOF9BO12BDE0ZD4pohCA03+pqFU6JWgrPW7DWnEX8y8GyxEo
i67cxXMrm/98OKsEtp3THHO+Ez+TkCtTUcxlWcsMhMpZkrht4MFpFxVSSWl/Tt7z0jNf0uMbCcxc
wqAnjy0McA05wCAKFN58LY+x8lgA3b4n6cOIF31qnRBdqBps98KHkVtPjhty6RIGMV3YIIgeIPaO
XiiRoCEpEbPzth3rb/dF90vnSeAV5uAGXuPuxEUI/2p9MM5Q6iKrS8Ty9os2MaQDG/uUsNSpJX5E
udwjhWCHS4HPxVzFpT6hxk9rZAMeq6qRlXqy5NuG3298wQe6uHow1Kz9u9+wLDBPJn5z5XWNFVGp
MQcv2YiYtdPoc4zR2AwHc5N7osVNdSfFr/r1U1WCR3i3CDOfS34mcc+t/f96dTA43p1YMWRAb6lU
dx7mFA6kfq7Q0nE95ECLYKzr5Ptq2lan6nIB0rvXSYZMOZ2AlbVJWJgz0pZ6f0ID0bZtIAFSOCNm
8HAyryqOlHJHuT6F/p66rAox2fZh96/HjD0cVCMaUSpdZBJkgQ9yVbIP5rdzXz0IjWUx8AR+lgy5
YdOWX5/Iz4lpgvGbBK/6MBS9ILxX+BqPucTdAs7djW42oC6WwoJXgJdTp1lHb6N+w+fOD9+ykAS7
4Iu9rR8sSsu5B7KMSYk5qMw5Y1QRAVcMx9fHQwBtg94dSh533yGSnSIL04s8Po4Ag4k6J4BtCnk4
GIR6WKsdo7qNctwrc19pmC9OcPYYb8tngedLluSqdyNtzuebMcpKz885yWilfyccjds6JMx7nXYi
B6BwzCLUY2HXmUxkOFn/+tfA8kC2CKMd26yPwtCzNNz3xAj34mRUXw3Ymyf0Lb9Qi8IDBlwVsdmn
xZ42vo1w4/XZI6iTeuPP5RJk//aBz+J+lhyymB8NBYcvi+qEG0Z5bQ708djLJ0/JlXGwT3opvCky
sIHlFJapD8upcA01VXx4smn7Si2fye4fvu40acn67lkLFqkRSITtV+L8qrZ92jmgMVbfxfihm03D
KJGmtYlrconlUejA6XJJBXn0Ns3HwBiPm9FzIdK2I/49EmejnP8eYwsYzdOJf69auHZl+/vYPjDD
T0pJcDP/pbty2uoq1gv+y3FeKKVeyyxSqmZ+S5LTIz13sXXD4fVqBO+YIKZmrLaU6/uYGOKrXTWx
lUZFwsR7lZtPUmTO+5ICWdTS1qyFpEPihnkvmIqTePXmSaXH/ARIFiMVq4JylU0X1HVOx+f5Xp5e
TeHDh50kOApt53LcPG2PGKQ3NZnwYKYdF6SLRVRI3gdGi9Ey3X3ChOfrhUvU297xYoUIElRFtulH
OBE7s6GGkcYiEbKTibiBpJ5LBuhwtMM/RuSQRIAXHA4Tn+uL8kySMZqFaJY4p+4D8cUUAOEByQU+
QTSg4UnZZZM6fQj/GacJrwlB0CU/ZGFRU7Tvr3huiIeVttHdx1OA5i1Wr1KICHXn/SZGm9fXU20k
/8dfOy24NafWTJX0RArpa8zB5DbXdPHl5c4AAjvKL7CP6mj8kGYcko0jq4e+GFMW88C0aYwYixTN
ZwKN1ALwLcORnTtQaKMK9Ek67mcjxfvt/HgXui0ZVt2g1O5pjFhPMzdYqCuyPoqvTN6VVCKsUJBJ
qD98Cz1+xKfKdhFjXIaWkjf/qkWMrW03X5g1Mydu3Ek5YdVtU6SdBIiqJzYwiE7tkH4gMWJDOLW+
whfDs6hsL8SeYf37NI9f/94g8W9EhEEdjvBRTMpAntdgwVsR/oK2Z2ZiHgq9vEd4C7ce5V5Pbzt7
V62rdFLgQ94cVCYR1p4UIXDgKkgohdJ8k1997W3RtmufEPplEi4iTETy6fnJaVhAp0Z4t66wunRU
EqHto4XKF82JUzDnGaBVVbNG/e2L/yfsEEDALi387LY7xpTCT5l2CgTxB7bQrr9vvx2g094ZCoCX
J5DUVDMj2Kdvyw7TIRpaeyCLggWGeIWWX9O/+NuA8slyIwJ/sH+PNRGWkXJnx1r69q+HfL/x5AK4
Xn0OfZLMXLAA6IriEA1HhXul1WmbaGXsDs11eAj+C7LHcBdpcvog7ScyPPPbYhsB4jU2CngzYT2g
J1b9QJsBe0Kt+gpEWP26/9psqOhJIctuVbcdIJ1x/2kDzqtkfQk3HjKBe7o3QFpcDAg13W3/FUvJ
+afM0ynbdQU+Tr6S6gZgPBcReb6kEbq+6zFyrk41ilJdQRK+N6ImDdtIA2ztu8lImEFzGE6lx1vl
f3CYduQTGpSgvm0yoP15VZSts5BneybYhNAR57h9w69fF/xKvPBPqzzAn0tyH4yKbYOvs4OxzOKS
WZq0Jmjo0hfuyMyz2IZBNX4iBHkihGR09kXzmFFLNpnzGVRCkrnoeD1O8JWn6xDSQ8F3Tt6xdt+w
wvZVaphoD6lv+nIIakvztqQ3PX3Qt7xcTEVPJ+rDdNRJlM211RdBR10DTQQ3Y7Y6BDB/8YMXw7bg
hEEIRZz2toTGjzltcZRYI8p02HkQUGMTIDGSPS615DRWLS0fvsrMw+im4iwy1d+KMddpWaCoacup
cR/wXm3DMMgHwrk0f4w1YJdTd4gECPzOiexRnl1DL48wE67KOH6zuCRWgVFaa7pp5ly/KDaNB+4l
LlBeojcOIHxPcDXXVa6ZpbQN6cMSTwIUsaR3pQUnsa6X18HyFq8dBQQ6xAEdOQpFjKDpli44QYss
coWjThL/Fkdm0mDN6m8nRCPv3bRXgfw2MPWJphDORPxcd4rHbvNbXFQpcCN7AUlfM+e73x/fO3wb
JigBhbjYBsVLUZDBMVydJq4th70qnpSZxw5TJNqsONLet2qw4B8nHKMMNPYQ5pQvzCcLkdP9/XXF
GsD2dkztzJ2423yZWQqwwrFHNz+rMeDIDbpWuzuSTaHxH3uQDHapPc01RyupxcmRTF/68NT1ibek
WibfmSsDe50jyKWnpHO7FGtS54DONic/xjtD0d08gGQjOaQKuCZrQFfAinwHUwlazdHeZi0jjwAT
tLp/WHssAsWVrUkJlJgebSZaqT1nVkXSGHpWqFT6dz4xzblReCMWrQYUp49OnAVk7nvEC+gowUpG
CgDntLc5hxyaAOSyGIg965gWMyfNwnWOw5Cl+Fgoc8ycx175tn3scZlzQn3SKnmXkbniZmX5SId6
2BGP+pp3o5nvCMYU3sfrHXhD1ciHvWJVvyKiEQnRGAQq56btkwlwR+M5YfEKE6CQfW9priHn0WHe
UZNJJlRIuqN8wWEWbGenAv9Bne5OjdKdIcd5Gz5/jvqk9vt6yh8a0c9Sk7Divhux1aN62qoyi08a
Ay1C7p7k4AX0WxKtAlZS1uNqHHx4QOPTXHfeJ0/OB/9Bfb9IiSy/V49jN4DCcU7hobVnlFyzpn5h
SH/p4LIqCwmPtrnxa+VX2Cs/Z+9R3JCHe/B71fKIupWK5Nn3ANbaiAwlJMm5K+SWPi0gWX1rzgfV
bE+wXDdXEnL1PqT5fwbrG+1o5acM0mAKHry/1Dx+APid9/6fJe1ssg7UeMEhyk/0mKtjqSx/4HZO
zLgm4gy8t1xcp9UPuHnSuBZ4YbpO2wS36kLiDpw70+ZiMEWnx0+gQaJPOuUBhqAfEjBIUaFkeTvB
NqcHbYSABDWKtnHiVge3eOG6lknt9Ip6SbnyR2etaPuEKan6U4wgfRjX+yDl9XnvxH5tjfPN4JUN
NvUxjCXV7W+EBpgvaGfnnZfNCu2qsT3WkcmVZ8VdG8v125aXeHcWUz2lScuccwv3gaFoWUKQ74JP
uWtH0zR83+7w9/rXohC2hce/DcJclW89/awLu7T7lcXEOYZUlKuSObe2av9ZP+pcdSf1Ny5SgqvA
oLnC2o7nK+gfIqpHIEJu9Rt0JHChGSG/APuvi7KcNXs4OIJz/sSqD1RwqyxheSOJk1xwBeI5AzWc
bIdAJif0z8dDoR5Ac5KS5sFlu9yhF4sxrczJ98Z1lYP5CG9LqGmQCwutSQFF+7+YCTaFCyc7VzF7
2r/JgChwG4WSM6X+cfEzmLFbtcGHa5x+wRpluidLCPxGV8hgCxo00MYX0UieRZ+ED5bwjNbprahO
CT7XhAsG2y0WzmwVFfJii268o0JLdxsPXTzlNv0M2dAXJlTcunXDX7u0+deDz5O/k3InowT8zkWV
OS8MjZVnyp0J9qfk8tsWbc3c63UcwGfwAH0+lAPvwvEk++1HHtSXb/4YQLk0Us5FOsUVGsP0kYzE
YrH2prEmNkuE5l8a/ISSvF/FXPfNqD9pAgHmxt6iQsSmcJrZYHr+aIUxKKlrdBhB7D9WhEdIoFKr
lhmwy9PQodQyBek3WnkMnekxVMtrXPjSuPwZxQYCHisTztMosXQeO5wWdF+z2u7eNn0rr+Y4tf55
hBw1CdxGJ6whwTQxyhr02/IQK3rcvEL9+ffAa3EeDVVdhJPM3BwcqvxTGYQysn9+zKSHHCmetZbh
3ryWWsPhT1STjCZGGCliMkGuFTFhCVugg7d7McDZgxOe0s5A2ZJH8LVZLQJsrHEw2E57ILHgylFg
HebjvscpH6RJHmQdRby9gNOaPhiICXWmy5csAhWmZ20zLdpxgZf6zFLEGHenwY1J+Gv7oC32k0I4
ntd0Q5DTDx6KUW9wVN2L1aKjzVczRDL5Ee3eLzEM9b/X67yjTYkV/tU0j21ZTnP9TZzVXIv2DAP5
W68gnFxU+/TvOo5zgEdh/uqB33tSxhrwozPq9d6pPbAGbkx054WNH7n3eR4pqayW4lcbRrhvI7Te
y3FLwiD2/fHSVjkhXKLPy+W4MWgXizy4MKLvOGHsgxqaJDP1uATUGKymFS+GBrGeQdaylLRR+Zpb
cUKbhXbEuUNLW+npfliOhqemfH59MnxaT+uFXvCHaTQXAAsu3cXxdye5+d0hkPQ+XJZnf/MNTF+C
4aPvHtrnnqaf5xEoQKO7bu5wnTfJrCesBEEBwmsttCoR3rn4Gs7QWvTspewFL63M+yBwc+0I3/hg
Wq05cH88klBa7frAh0YJm1yylyqCdwd6U9VtMM5FxXpknxRngkY8+I3wCqsqmcKeP6RRp3DAJCfU
3VjUaiqHL1D89eowpXCBTejhW6ZSduIlmYmZR5VZ0xoTbDW3lKl9dlIGbBOEFsgLEHkF+2cG8MUp
RHzIHSytM0yArSH5HSJwNZx9ZAGbYYCh84IzA2n2gJp35Fg3VKdLoGGAVGjjsPG0IKHr6m/zRV6n
HfjD7vrWJdwD8G5HqutiwwdTiFqXb++AuduZTfb3px49Y8TFK6qOlZpF0wwaCXEeRmpSa450FKQl
4b9lQAzZMQPXFh31i65I+9n7zVFzAiziPsbqWrt/ljGU4j5hrS33kfBefzNfQcYKTHzSqfBlTR48
HQfpi6usty2ssvGmdCFkyGwMxMkmpuOhW3er5UtvN/JtARk8FO8d1Fkx0RDUkG+JIcXXVAT3u1JU
AnWCEC7m8fBMqJtaXAUYdRZmu35vODJ0urIC2Kn06lxFmjt9uV73l6iQg7UR2Ylgpj36+/HMbogm
76YtwRbDUnYu2plxpcspm12mfl1So81QKY5LGTbQJMvqqwmPVfbHvqt7xcSNOLFDgh3wbS6ERWhd
GRTtIDOvYw3tMavWhOHRaRyeRFh8QqIeyocQmiXfLcbACM0P53Zz2dl9XaEiEO1lfAWkQDbmsQ+V
aXJU+6p87XLrd8KrkshIRdHMdw1ZAB3+8vp+lIkYkWdeGfn9a/2pvT0oM2WON1SjhzapQdYNiKFk
FiHTX1idukLFuSBMXPfKM5LJ7B3Q/QCrxVqW/gihRDDDRvA5To3xdy7OPbIB+aFtCJZ3J9V5pcZZ
tN8PY41fhJILtI1Z5iqvxJbfwOFtUmxCBPnkXsOPsQ0Liv9JJxh8LXTcsSnOzv6YHmRV9ZKXFV4e
gXHPggNzDBd0S68Fz9SOdIblfpmFJDKPK4QOX+fyPyUcmD8daU1i5B2nOmbyJm308MQrWnuvzrwz
KF0AbLBtRFI1HL/EwACoIREzdNXsbPwmECibnzv16OCA3cx2vDmg017GogFvM6v5ym9nsRxS0BTZ
AWsWmDY7VrAIY8gpyO5waPA5TIdwb8EFL5GUbBFQHmNqd72rRP/0gtmkZqYrhwbuGu2gO20qh5ww
zitUTWdtx4AxPMGyZJwOeGHeh8Z0/qcTaTvlQqckpqlI7sExsgo8RQ61htU12ASfgSqyge5KMd/l
XYnIwvT6TVCQCpWLA4qVW1h4GsdwJIHE6y3Hnrv55IT1VFcw1xKAoeK3boAgKCjcCQ0UAnzpyG8E
kxl1HX0BOLtsHBVzpUsFG4E21qVXPQAatXqhUd5B78gcKE+2iwMaRgFp0Rn2Fo9rlhBhI38ImiUK
iQAl1kLOcTf+RRkC8w29nGnZ8EDqwK4lLFERU3B/ZnBm4C+bH68Sia48hgD6PHtrzi3Ge0TQ/osb
eGCBVhDe44YQ02cTC68Mf7XT08bzz2XUgszC+w7Kso5O2TUxWEybaQptn/HMEZzogd2TLIBWVz8b
cKxqKErjPB+cOfBay6bl268DQj2XNVJ/7uvhDFAdH36PJ20K9ZdhFu1Fe4VoX68kDGhFIvwaWc/O
NEHut6e8HuPK91pOX0U96z7vOQ8EvuimocFzZqwXm18fyxigKGXiKo+dGaAo0svz3CKZMygDR8ds
go0ViBt9Xw/OY7kvUq0w2fuCerSSnq+PYF0co3JYdsdCaUrhkYiERIyGeb68819YvPLGNmnIGzSY
wHK+BKbUJa3iMoFpAgu7fgT32hxHScaizgeRuYPThjOZH1L+a1tGEa8FrMyQAgOaYeT9MOEfz6tQ
8JVsF9RHiaaTeFcCeex+CwADyeOHlTbKkG6sOoDH9ax7oi5LJH1knfTi/eF9AoYkNyXGqxQe8etX
cNejkKtcqxeRxpb2ivXfe+2jCGhnCzjN9EN7XOLM3oyUoHGywu/oWUpSd+S5gK0KUSJYp6PR5zCT
xVtl0cRIg+zke/bDU3M1cNo2OtT9YwMxb5H3WKxklkkelqTYWfVlKshiPvAQMDNIGW5QZbcZVXhN
tSl8omSqX7BlxooywI/93ekdhmS/BqpjI5uyHwhj5FmcVrKUnmO2ySeXmnWjjpBlhqv1mgvRWK4A
HeXcpmNJExpe2Q6+8QMfqyPIKzYdaUHNf6Sh9jl9dhwHDYpMP9FQ/ohTYZwlJjT6Ax8TvJATMyH7
+lPFXlYBTIVBvHbqRqIvD57vQY/WRQRSHLCfkpt+wM/wGyZpTnMlE2kYvfx/KxT3UDg0aORKgkqb
2qjLFp2S4wmZMb9Dyzj+t3R4gmtE3o1FddTb9tshCYf11eXnRRi/7rO0yG+6WTtI7tFxH9AHh+1w
3mQDbUBIJhTzPGbUz5hAj+nBJESUjecBijGVTP/N/9j8+1Z4WNM7wtQ00NoVUtdkOcCLStZ9ugXB
43WPPmY2lm5EtBlubGLUtptU46FFvWAy138RWpYDYnfUSdiAJab+ITa5vWVqusxeIDdVDT2FDk70
JZ1SfeEiV4RrT3sG00mWCukJwlAKhzphI9xOKs90++DZjl9y8pxUNcxzylEq/Ekui6WZPa7WkoyG
ua2RTH4A37Le6wT4C8/Wku/TxjhrZNDKuBNJf/WPjXmv0nfb0B93QK81Z9ecuD2n2R74y7ClOxvN
aOOg/bXktm1syujQ/BvVjGvE18qKt/txUEIGpBOLA+rr5xHIdZ0Topiw9cz6CySBrbXtMzLkMb/t
SbEBKNmctZre1Z+ZPXtsB9wcJ6+nMdwfywMYODltW/WQWv6/b12vgfyrHrDboXNWnB27Ry16qpUx
1ZX5kZowH9N9UzBvt9GpuAwmTZBNjBd8nMrg/sH7jzAuEOMNX4DyQ9+2yIOp88OQCzo2ieVroISu
6yNt3yDKcDUbfT1pSZSH86cFaQQqB8MYlELbqqlMJ3eMsyqaneOHMoENeKf5AZaFe9Mu9herKTr5
SDIjDsolMZ0y2Sl2Z3H6r44PpQ92kzxp0vK1ODo3PVyx0/HSa7wqT99aNKh6mH4gce9CBU/CFpTN
4v+C3jlu59tT8E6qdJmQoU/XD42jU6AQXONexREpPDu4A86qrOn6J8OudIf4p0mxQrLBTrDAYN8z
3J+wGWdw3CpxFEb2QtVSidAZcZ38lzdidL9v7ceSvQfhaAT1JibKEccqHt2mRVT1RxqyFtCoLyc5
2EAw9MnL3NM1UQdtEbY0otJ9GU1FzKm7pD486iuxfv0xtaI548ggnBvvqoq7nLb/QgjDbsNEWPDW
NZ5K9dwbmp0YfJbqX/3MECpVyKjBz+JLTSt9lay56oCiPPuwq9Nsnwo6gi/mw19YfQz1ZW0vWW+i
ZgNFvp0IitbTHwrw3WAQtkc36l9KV0aZhH58WtvD6Z2GZxf90a/kynJ5Nmyb8FU12ZGh/1YNJfe0
gUF2KDPxdAtSJSgHJkDVtaXQioMo95DOuN4/xLI3gur4b1DZsTD2rC4GdKl3aphG7/yElKIkQGa9
P9msH9p2rAHgowRPKXu7fPfkf9f9aAqyy52+vO4+oCPmf/NnWdQ9jp1c1RyuIgA9YsVmTJ1DRUWc
isAP6y5rfBFrM0jzW1buRjDscpAU5+tLi7Rs+/xasGOsa12SYbb4Oc2IgMmt4SbeYtbMI6INUeKv
snYHGTcu1MDLuuhCn/xZvSTrWh3Tgu2mTNpKvBfTf5bINBR7GfVeicfeTHEE798PajSs2T+o6GhD
D0jIX4/cznN2jd/CLd9JzQki/IiZ1wLoOEsItusCR4cTznmPuXMS71jH6mOphAse24t6Axb+6RWC
B+Ywzb9SiQWSzLy3mMqUXx9jXQTr3KQ9TaI4ZUh/f8+0n5I6cPtSihYDLszsSPsUqWhtI6h7iW3q
n9PXeYBhER/Q0yztn9rSHNvU3nKDJniYJ6WGMOergL0su+FbUooFj2hOW2nWB4nfmkLe22Qj/rS7
g0Wdsf9bb9mHAbfpJ4JyZd1HVaCMS+gCPx7uTHydws3tnpa7TSFFrGRNspoVViK0tVioj0495R90
gTGuU1z+3JV2/2szBE84GvLVIpr9f5FRCBiMKDIsqfe6Zow485i7mZ/oRFci+JMgq0kQ79azZbs5
Z/pu1lEvqHgXOG9M6WnDPeKcXV78V6vG0FogtBFqGxwGHYqfP8NFkHkXzEAvTQ5upfvYNMgpBS7B
ppQ76FnPnvxUpV7AV69DGw5gVmuK9hm/3KT6D+nKPZQyjw+oWav/t2I61kHRxrWpwWHpk4NJXPQ1
oQDEQK9W0sm47EQqcfNCAm9cxNXFAL5pK9eQmHTOQCFZnvt3cWu5NX63fWbiAMy5tORo733ASdNA
0Lewq+pW3TmQVOI6Ou3qSLwhspdkUbxMNtrAR6Jpah42jCIDjtvYZratOJgT5e/n+x1+kn466ql0
WzjmmO9yQ+dm8e4tZk6LplXp+QLrc5oZ1o4lsE4GP3cTxbGG/j493lPdrKrWKy01i3tu0ft9VgFT
tW1uak0CWx/v5ULhQJYlkaKj5v5J5xxY9PDRfu2DAMRXI4fXnJNah9giK6Dci0Khoa7lpXn5sIu4
ISFkv7fRzyohyAMcw15yuTbs9uY5krtKZLCR8msmjMWCiZ96t6VJMXpvj/Ma1JpDynOQEllCH0uK
W8KADoP+WmoUdDFA7u/wekR/wMlzf1WET8u2rF5xLv67FMouc9OSHekMn9pw1PWBbMn+7h45eclD
/yDMgwQhRwSitWSmMmmCWAHvL7sLbxC0m5bb91eY8saiCq25E8ePzfsZpYg1JiVhy9cfOnsoNxIz
JFu88tl/XidICvnoIwpmFiG+sVa30fK9DDVzba6zRBIJu9rROzl2ZcvxI2NygIiozMIf6LuqQChk
hDGoxrG/XAEcLfXJH7pfYobjLXCXlGeOMyMNLY/EwspLPqPDCfjLr+9dZDSbE32NGqWoaSsw4nd6
HRu5jOettUgHUBvTGvzytcUuiwlS4LJu6dnJGj4J/32I1XeE7Nk8XdzgcC17vVZyjm135Zco4YSE
VSGf7MNBGWyQfJcLSoDA3C9yTbk166KMqVWIzI/EcG4DL9J+zP85d9FZ7V46X73QGMrhG1lZWzzV
RK6+SEzvyj4uvLIb2Mpak0wNt2e77uXU1EaMhMgurz3JR8L+IY96F1u8omFr/eyRcvh8AVZ/OGlX
yoROou9zZZRrOvW1hbxC80YjDrrgkQOledpVR7UhSu4RaJWcNCDRo/bG/DPT+ThJ1tfTo5iaYPNa
OwhErWibFrrgmu1XYa3lO7E7W8ciaVrhIMobFUMDxhOc5Xsoy9TeS+MeLcUrUbbxL0jPdBeC4gzz
D6Nc0KSfv+PCV0h5Ue8RsbbfAqcuq5bHaZ0dUSL+hWnGjHL0dgCUovsPpIh+TQpJ3bHDKLBd9EyG
Ze2l7ljCtGvdANDz6UaeHsRQEpwExrOkjG5/ycurtanu8toQQjJnzLG4FVOyZTa+Zo8pfRDq3A8X
VIErzY7Qijl+NhaBj/mdcXttqLTkqn3kTTYo6g7vdMrd231LJpj/1oqsyhnVz6V/1+qDVlta1FNV
Im2pKImSuL32XcYhh7/IzngzP6NrUiX5YT7ww79L2ShRNYh9mFF6udoUvuQp5tzgCZpQHzRezOMu
9cP5ugA3hldGdEMTwDQolUrwswFnoiTn5Q2ujwLCitNMzb6Gmm+i8OGeaE1otpZv4ox93ljzTRSi
oH1G8tL6gwvRjTKwHe7Am/T4/ALwaLFHHK9OwiM9oc67pb5C4TodCqvpTERGr1klR9B6/Y2Ra9Uq
qnGeu7n/vkqZGJosSvjdyZ67kdUu1veiUPNodG60D3bH3jjQw7kIWcEMbFbgEKWyZzdGJtn7W0e+
tYvcYmXDWIkpf5CMFuGsjyIEHWU0zh78ACNzOSOAuSmouhI39l9KpazdceoNA16UFXa2LlHqF5qN
q9SJrdJmdURFaNKEvHar4gycVCF+fs1wGKe1c1l54VIgsuc6V03RLvKOEsckYTHt/pjUXFVM33PL
kTwESLLLuM3Ti1Q/L8v6Jk8v3cK8IDA9POut2lKly3cJ1PbDW7S5yyP92VW5tRoRtwwOrkCvi1pQ
r3njcQ6r+ePvZ20nnAAc31NjaR+iPClL7I7vrW+JHBg0f7nsofdU096HLyZuYl+yBk3GxG5c+luI
264zjnFiHmUGzw6xqCrukQ+FGzDoXixmONRFsdYoffUXVwIga/nCxEZDEPmtjbpoOU58YtPeVKGU
lvunmYjERuxfaKuURA7XkPzhmZDyG/gsFBYUxJagWXGmau5rX7+IEzlMHD4Nv87QBlgUGUvX5oYx
tw+CJDbmSO3g/E0HmS9jrl4x6vALayv0IhUZMlEfgUKL+gltHn47C+NOnLg+k4pFgNxDSWEBR7JG
nKlW08/SuFIbXFJGwevCxL4iUsf0shmAzpaqeRcn+bUnQxvjRCvYdzBK5cOTfsiLBUDEpy0t2whF
wfrC5lQkcFes7QxvZWv0UKCLC9IIYDaWQBJ4MeeyhGpDHP4yARsSAZAAET9CQ8CmmTe+RlJWsIn1
vTDguwCtQKuov/o42ZXjoQnr4Cn41zFLb5r2/xu5e1hUAHT0sABV+QUPgA0W/kpF+aG5Yjie+49f
BTprg7mEt5Pdn5ITw17mSeniM85UqADMPFJiysO+LrSTZw67/gC0pu0jO0TSj/8snQFquKQfVJ8F
eUji3HUPMne6msWB/BcDI1b7whPSaw0gahDhnioAhS3DsZJACjK7eKPOev7mKiBpKC1hu/BooHdY
dYLjb8EO2QzEucVAKeML/iPv5yT6dc60z8KAglV3KnQgJmOKGLtLPuIllfoKsDWzf2ya17uJTd5s
s4b0WHvaJYuaXK/I/Hm4ilMUBX1+5VOtGLf8R9tMkAZJwzK07zMbjVo+QJ808aTx8+rXhLkHstTC
3FsY2+WEYsilmTnjUxxtm1NS2k1c3qUId9Q5jvxTBpHsEpPE5BfGZ0WBqqU4j1C1dO+cXyj5SpmW
HA/88BaGf8iiF+kaMFXmPjrSo112Quqm4e/FNIY4NlMJ4f8tlaZR3kA1J8XRb/hAneQ4CNeq6r+3
ojYTmSWVH/guAwoH7JqZAccrqTygPm6gzr3qjKqiPm1kIKqQX8VDDPZKHKA29ovNaypxOlgnQ0Vf
cqyLrbeCOt3qmtSr9PAsyjEcJ1qrxgKQ0sBiIR3eKc326uTQYJvpI+7WXGd0vNaJiH88ox6kTJ+D
Bup1HAk02ZQm0Kf0TmbiJJDHnjh0LyY/REd+uTYP8bbacn+zqmW7dqxO2YQ27hYBnVpgxSy3h8OD
kXa9aIQcY8NC+tMpcVhWSy9T5MP1dHyjbahucs4OcGR+WYahhquXcnHpRgl0PHREoTOSAQ/fLmwg
5JU+y5Ae8h9+Xy8of96nonvAYY5AZeJvmlEZL/HpycLd6Yt8Ngw+2GjWLgXShNXJzLUFG6JLS5e+
sTmIzr1KtYsQziC8y8LHQPAopMqRWPbz+Csdk2P97U7yFPWxVuZ+tgTQArtwwaHV/ckx5TEnOiup
iC3Ns1CIpxfuJ9Rzc4/SLhOO/sn+iPUvK1LUZyA2XAOc7dkWTocYWUk+XMU46RDGGD26Aen6dj+L
UwRqPDDKwKeNe9zkRFpUQ9I53KmqM6f4rZNmwgMrUrFMa2Sww29OfRTHBOmGfT6kxgoeQXWOTzfb
rZqJDA9QLwlDASQn7UZOdv4hbp7Ju1lXgU7tVv/C0sOe9mXwqqijQfX2Y1JuettWftlTxS0IKb8Q
EGMIosPosOU1k5tVJrYKe8tlOPX82puOWSr39AlWysUj6YbmGYzSlejoGY4Tc8ZNAj+aqhQdjxa6
XVQJ67luZUCUWeTNw+r+QPvWfa7QT/sBg6xnSgjwwA/FDUOt+DhVFOgg5V4dbS35bS7E7PKHLAhk
PEXgxcoHwZi9nazsB6/y8G8Qzh4KGz3oI/Yp1eG57kIiHtpvufEWh6ewAMKV1yMEsR7k76FZCjjw
lDUMdSxMeSxkc32ExphUA9RFuxJt5+FO0lpQVcFEVpKKXfFCApznjiKb5quLHKzxuAX9WoEdLcgi
WhwIxgIkAzAMFZ9nmGyUcdgz3fm4gaW+HPr1QlC1QzQ2e6kyjte9IINiHFVswwyXTqhlgLH0VMJb
K1Z2XuPqZS2TJLwxqERW3gpC2+ydDpQp1/v47JRcpLI7wK6oYep6wc4dqhfvsVhSpSaKJhNlYO2x
jYZzcB+kwdv9NGmj+ZZ7vs9vR4anslBggzyTYg4jBJL1h24aepC9YqOCJFIfCQAwldFqXE0BSfTJ
j2/PRu7J7RAQDH0uaw7TD95b/MvGabu9eKbfToUunBFGytGhncR7lDQZ06tsMpQ1GUZ0PlaLNotx
mBMWL0VAb8M5BeHv3a0QiH8Edf3bdG4Jn9Sl7rcksmF6ExzikbCuDhR/PbQBvr/GEQm9Lh60CyMU
2vHTbrc1Jlb7mDyiM3gY1PAePAH81kh7pnzLYEHgqeU2FglHFfMUz7Yti8qXg+PVtv4bIo6ZNABx
XQT3J9ZrexBFW2uMsmZdPS/FFU3UCkRetILAmOtOv2uXGKLZ768/bLdIHAn6CtHF8SuqpkzWpDbM
J6gMzfegAEfY58APcbvlCPgIJN+snJ00xf35BQJHaWCz7iJOItq41JDDfReikaFtJtoBjRFMiA6O
7ZPKGmhsUAvWP73caQFcu8G5XIyYjgYuQwqfUhVTNBIX38eLgIzp5OxdJVfB0ozXFcs0VYjRGxIX
dwpU5KoPurF+3wp5dOh1y8h7HuCKS6emkemQPsVPtSGoM0cKDJubxgr0uxtEYosNFeZkBGC2sIX4
oGK6OWZyDhhEcSZhTEkboy2g7PIDZ2wyyx0pbyBWvMrwwAz0PtzP5dFEIL9Gb3BzDp+h2ywH655l
MVxjicaDRZj9Dt/sxNwak3JwndZC1UiHaM0PRRulc6pczGQSFxILh93jc8/591WcwISMH1b489Fj
QJ9yBDtYV0gBItkMBZ8UNvPDdSa9IU5ttUEqmPGS71O83X2YyCrOygYnKPw4AbPrXgaQpDgP3eXx
9gvnp0Nu0VzfnypM1sfHuYBSFHRD1vTx6OpoEl3AdzpD84ya9Bm9oykzbJ+E7binH/A1IRxW/G0V
Tuq1M9bv2lkGt0Cth8xnJ5h0CWAwjY5Du3BfzOOpTOGTmrs98zPxRzXGEAOXVgpPq1BKRX4ZqRHv
Zao+cbeTg7ny4PZFr+hHJCwTgXWPAeNaoVvD2SyGU9MhmtSrTRs42c/J6kSkShUDuwmumXhcM2+Y
/fwqKr/JDgCZOfBIW3ddnyIO26iwO0j9VRVI8UyKUiGojRrrdplJpwYgbssdGYnxEzpf5NJzqhhj
8Kon0t7hbnf9YoXHUdO0uPbbkGlcu27lgWbdCpuMb7cUqqsyeIKAJoivjki63O+FZmns/bw9gf7J
M4FIZy7eybQxB26G/q8XsF40FHacUnu3g2QEogWuhS2kUYtQXPn9hq7Xd6pI9zM/wTfIeBW3A51F
cqbnLgOPioFOYQLmR8nsZAVe+8/NTlERIsuHWjooobdvbKnPmzChJ1ZIdTmAbOzibjMjgVjOUSiw
KjTX5VEtX3YipE0BhoSq83ArTK0HuuoBucRDUZFNjhK4jNDzCZAC1Q9LoazUtZ+4M/x+QiD2Mgpu
WoFJAiXg2pXGeZmplbIAWPpxYnOD46FeWEdTbVMVrwk6gnXlDaoVUECU8GBXr27jsdogEsEOG+QU
7+yRgAAfk92xdbBy6V5NVCG32zQBvSHreTdhCrg7rCVhVG8oRUmMexP/9JhdTQMwX3vH5MgbPJTh
9Tor2ToBehkCfkq/ZzlcmJg4Jww0JbU559y60hfC94ir9EIeh16C2VKWT8ANgoqDcHpLpF4ATt5k
Q+6tB+k8tAjcLucKjRxyKzyyVGJKRoNbeuBVtZxAXNzW51ee69MH5h5nUI9bI1JMUDGK8Xa6jnJZ
JB8XMIVi9lElRXIKQe+WWkItw/9DkByF+sRcB0NMNEpL4xjmJXvbRgGoQ/ZM4Zean6ydSw9+ziQt
Ba7Tr42lMh+r2Hsz9LwDWyL8TKE24+uWrnNFafa+TOfMmU25zXF5CLN1BCP3FEwvc4SIXqwYIUIO
U5GfsZTHpSsW4wxCeyQI5ykaGt+bZl8Rf7cVlX94yHHaEZKNQl/m8NwFCRbfkshX9a/MoceBvszL
Mzabvn21tSVic836wols070FCwPnYerg5gjthswZj3pwIO3z4xuWGhJiPFj2rI283d8Kq2kj6ZN/
m2EAVVUhoIH3QKmTe+tCaHV9bL9EMSX/VHJNy5q8NW9f9N2DDkoD297M2PoUtkbK4kZsG7XRsscH
i1m/YpIeMSeP91rwqShf65t/1gR57C3sbYlRfGa5hsSIsdSgdMeULEKQFs4h8KnSqpstJ/Je3bvX
MiNliXf3apoJ3YgfYId4bUWTNCpCA/GaHdNVlng4/kScWJ0FwMGiMK2oSKXpv8xmHqEwQ47Qmmw3
r6mQFaWQwxrsMry2Kpk+YzqVgQy9LdaWDSw2gcE8VC+sDzdfeqcsGddMv9QtlnpPtU5pCyZ1iivZ
/FTog5brB2zMi4clqhBsfQ8FljcWy5Kkdq5YP93WqFuiFYThtYnJE1K4n9PbpvXrvHtgdvgg7Q1a
Txsud+mnfFSYStPcX6fAmh7PO9lZUAOzraFrUsifeXt9s2WDW5NoMWjk8af/zJvMxpt8jHIJIIek
S0yn+qNJp6sF45ERceLGW37v7BuhnaGO860XVFkGY9EXlFSwBaXu1KnLUU4Fk9q3R4Wuf/Wb1bch
GWBK9jE5F2F333Be6sskA9uA8jltWdfYE2rqse8o5QpErJ6fCIf1DvzVOuAjVK6edBTHFGieFRuo
SBxaImgVpvY+cU0VqEtck0aN4mmaK9V1uKnfgIallBNU/j5g5zYsf0PwP//1HrIiCf1UAxTCxCKS
u3zgAiOZuugpuapBAd5OiraaZkVmcRN0XwMeZqxETu91QuRQOTQkra7wGhA2eTq0+Y2qIzrDMM+Y
NUi7565tZ4e1akJzy8R0jI4toLQnhgwVT0c/FHK+qhZMcXf8kTYUj5wRcox47AgCdLqglH6Dl/Fh
MZo7AN05gFU46c4bhccIQMSche1P4ok+0+HS8SeyAl4R0rSQkatnciHWkgeNj8EkEGypllyvGFjZ
sy6pihEmSVurLtAX+xxsKoI3ceVTXCHyFcQVyYvqefaYlN9a8xXM++Rw+W2roKH/Du6kc7Kp2uB6
Dgfx7nVwlaofJ6D6Toarl6DUYnwDSp31jBXWyNin+5b/OihPiPxq2CxHCmiAoyGOa31qkyj78ZVa
IVRJw869xx47ZeNoDL2cYWF1NsZIENLpqJcV+fdSqzxRhE18ty1/9thwd071sAfcHpYaYFkrQ/du
6AKPZZK5nMlCSjG5ds1QktL/h2Vbf0y/c2w3cZIu/vDgAKKoELNpvmo67lVGjODJYx7iDZoNnqoA
HKU5NpOMI5PrmGtOlyZUsM/IYRohTCVesF2pz82H+6NfiSDAwa+Pps6Cz3vY07bl4Adcc7N1LR3s
KwWe6M9teX6rQUp4GiChRnpTQysjEYqC25moaPKUnZy71JNt+O7nbcgJqb/0JEnitbQyoJv2VZHU
jxxFCnBE1M8Pat1C6YolyF/Qx1kNuvyVzItyPoE/+isCTiNA4acABO3B/cha+xfYS24PhGWCQbN1
Kf7piIw8JfV8TPSwDuQaumG/XHTo0B01KetzvHQYY6o0du7h7m7EoNKwNUav4G1cZuSeZ2MLnOP8
MUU2zEPxoFWRWoZ4oCID6e+fhriCV75EHe8PEgGGIJAFtXF3wNMptpae9XPWeVchk+I1G3j+utVk
Pai5W1B68eaf+S1QpmPVh2DdvMEw9h4RMX58zpkRqymu1N+iu+FmduJ/YIubfWQZnuq3zodtSQG1
99j0E/TZo8PajkkEo3s8XQUr2tPAONdAT7/SqyT0MFc+9dm9BlTWrNofR7gfqjJFJTI1eaYM6X8w
61YpUiAwXeKBK/+GksJIPwNWaewVFLyrFlPxTkWujGkuPOU+eS9xaqZmckuW9cAvbde7j5Gve4Oi
l9rML17ghSpr7EFfgRK3oGS+3hwvwaizn+3FmJSF22nf0fZOfV1zUC+tfFvJdGAjVwkE2r/OnLke
LZ7cQGpQMsW/dAkkl47fpEpanrhs8xP75+xLBCNx4+keL8HiXPddVPTGOr7/YIbviPoxnQblpx0U
s2/nyu/BEp7++ObNgisaSrtjaDetpEBijh+TTtBCYdxpDqtRzh0CphtIGQOHrHAkc+Ry3VTk37Ou
8k7w/Xo5M7dTjYUpMcrBPVHyETR1oDWavKL7TG01/r+42/VEnkbOaMIzDqYTMJCsIToYn8dyPuGX
IyePvHPtaPoa1GeUK27QT3Sr1s+ml59dQT2d1Su5cmx9/O8i/P+t1hZ4oeyGqj/HTOkWumMrbg/z
aZf8AG/iXEKMxegBAqxw5AehbrAXj4jtjxznWrhFQMLWjhJbDm5LDAnoX3H/6mm5vEKfvueHvrTk
xpIIjgjkfPaa5fC7Vc6aNaAG7aQHee3HRxwIpMh0kdt3lS2D98zivmW9swCTLXS/1URM9OyobwV6
jWbBTyj3ewX1IlCvPwaflFMBZRNng5VXr77Q8AoWDC5ACh3Jve2Atzl9YfJUgviXA506GI7sehsV
SvaUk35YnCZ+l7fomG+2FH72y377QQ/e787UZChtiQeLTGwBH9ktTRWcRrouZMg+QmA//4wRYYe2
67A4QobDlyarf59Zvvj3/EgeLPvKRg6DLBnCUG3t7HULHvuU79AFgPFw3syivm06rbxgME1HwM68
syzhVQ1EqiY4Ucds7mqvpXNdVbAraqAuSNiRv3nGzJDp11Ixr35iCb1hg4IOWGF2gGRknmoNYwN5
snNbwuO6VqzomC3UjuH9kyB04ivLu1/aJP49mEvMNjUH5KDm4c2wv+AaKlPtX6qIVOsEUlWUeyyW
zViiTLWtmh430btRUcAL8MD6mfQqkxKwgmWwg6vNpem9thu3VVA8bxqhQiX/xKznDAOJgzeSSEsn
cQmOqIFPoBpnwhJEOYt4p+m7xrgVl+kwmwCoA9aYYXptuGSyeFvJ7oroDqqcWraSqWcmnKdAGtUI
vZ54Fcu1Xoo8/sbgtpFkakOiILqZub0eIgNToF6vBJViXHh75Eu3iNIA9oKR8HssOv47hJ7C1SV7
2mXaI6nMLba6DZ6UlF7OJScrHSzLPKRjt6rAp1tF/OOhmpLYBXJWMAKfR7A7QfJL2rSqJl19z9Or
Jih69G3F8hSWehppGgzbCeEMUCs2uNOevdT1vbLkWRmjVoJzd5ArT9cwVwl6XcsbsaeoJq9fxOKW
xqNiYeF8oIBiz84TkJEI6tCWZa0C4aIdEDSZwvigQ3905FuXxL/NnmFn0PCPu9f/r0zqgxMm3AUO
1czMnizfVMCtFOUSY7dXfK+Lgj640oReTC1rRdIPRJ7xgcs8biBU1P+0cnsuj7C9l/E8lotrVzVR
kdJjgOORfLCq8jf8PyLuGTvK2eBRluuk0g5ahTlFjTWIZONj7CMCKpVeBHmCJOWwKthVFgGpZTkZ
ABTGpwpBI94v3YBfygTqrgVzZOO+fyQHgSD73TgFEJkZM19ZjsyQh09AObjLK7AltJx9LaD9SOtt
6or8sEE2BPTDU2A1Cg5R1MzzG8/kJZ+RirygHpYFBz9F9sJFkxIefvpkxLVQovJ7kY30xrkCnGwi
U8FtjGVDVpQPMVl2ClCGTBNgtRuF7YNvjFLgXrG6qfEEYZWP9eHe1a7Al0xMufPKljnjpQNqveNh
DtAk5IFC0pUik2l3ckIzwZgGYhNUeJCwWdH0/MoXUBWffQk51F7nL4mnFNloQfz+pICSv9y9NAkc
PgOZ8usEScYtA97rPdns6CAgUMcnZOp5Rl2W8d95G9RathTtMa7FygDflyA7bKXWrstraggAfrT1
JFLOoibtPadJ8KDWOqD9rLHf+qPwHA+5KYghu0Ec75d6y6v9iiegDCOMcQK9Iq0oFzABZrHQ6m2S
E6XzDkM3pGOb8AiHRQJeyWD1hGp6QvMvyS96umutoNY2RPYRzBW1sH5CxUFMM2DApjjcQJBQcZvb
rzJ5NeUtHv2MZhUZI6Myo1Yi4OWlecCWnKN1Miju5zdNbwmBwgBBTS/QN1CtwA+6dD+Q43eYBAOb
YlpRJnuSbRu9AgRfAuxu9Ru055RNCdg9ypjMein6uFaShzpQ/lbyptUZljg4zXKrCUvxa5+HzKLi
zLKc5VfMyqJthSSaPIJa/q79kFytPN1ZYQNh1EO7ltQjcz3FUa9eejBRjIU04v055rJJc+8VkmNZ
KOGQe74lpocgCRrO+mYBgaLV7OywaUlyP4qpARx6GR3RS6FaUiRc0+ecC7Ih627RyHeNa05twXtY
QRNGYGVjmEeMuMhBl8DgirPtvNAYX+mFFORq860IdU+NTzer0mMpwEaZbOYjXnt9ykUMdOrSAZ8z
3hKt6XvVJoXKJjWQBm2clnIKaGcBnCSxTxUYNdF0R4szGSm7VCXpJNGtVbsy15XU7iCpcDtG9C9L
7If4BRmNNBkCyPZEf45pHNTzHAvUr93q20fRf175UXU05JTJBsnm6UQkJYtP9H5OFNlWi6RekpcH
UUGlh8aOcm2VkzpF5Cl74NOApA53X4rtN+EFC1Dp94JJF2czk9kTWc/2ktL7mZcVTlEnwWKFGAPn
+HCEGGfANpySxs96Ix3FAVaJ9eimkwdVehVnDUdMXlBtSfMeNLOYVqbPRepOFbnIfM/ggJ6J6x94
HFoChUWlb65ttlC7Ix6iUkt7d+aciL3o3f7MzSrEEcJP1g2wDMre0j0B9ujw3RUYbFEwZCGVBSkF
cgH4VMB1SPQIuv+AZFJG+KXEkWa60T4Td1HM8ZUV5B+WvAiNteN0FHvDuUD47DKiEriyMEwT5XTY
KjMoHBf58M6kIc3GjM0dqPMMZxxQEL40etb77y1PZnoqTHC0pGUe5U7mIRhdQokHfz0Xroyysau1
TRvPTYHJBtlvp+L1uSteRsj7FHIqYTKtKXhZBWMLr4PMxahdQpyy9ronLvagrEm/N9u1Y32H2UEY
0m17s2qpkLoiq2D65tCLqsrlQxHIA8pQXGE+d4Rw0NqaiLfuE593ZfRTmzf+lXd8ZUBQjJcgyijd
9ZUNxibW8E66w7q8mWBbmb3Xuw/k0yYXP2jzIsBHZ23uGe70xQxK7kSCA43v4pd+IL58k1orgbaw
2oObBQYCwEvE/5JQGl6Z++0/iBo0TTSXQdtw9wqaqbUwWtYuMKRIEjlGqjZ4Fj8x8rh6ogbuhngo
8H8G/hZVXNt7wi6sFhNqDgSnnE47kxmOJUK0EmrtMxut7snvd15wtb4qlIQ4gE/GAK7qgNNP8Jfy
lFoqkVgjd+3I5O28O7iYjSIrYZUzYySWoKknA3TiNXH8IJm2OLwikdaBXBb0hQEJo15x2Lk7mt5g
z8j8SJlSiDmHqomNP+m42nqkvr1SGqvPHc9bKG4tJF7S4A83DolU6QMWw18IhYUJy+2HYoDkYlI8
NV1R8XfUfngRPBsHEcUaGOUQ1BrQzS0KWIK2usB+Ly8hp1tbxwYsd9IDqh4kPeTbOvPlmwjofYnB
keqp/9AMVPujQoXTf5EiJnZT4UP6Ov0m4m3GAmpXka+Dnso3nS/MpuEmupxyF5jsAD2M1Y2d1Ll7
tj90GZiw9rZlXiN2199/CkCVHBqupAjd2KOPb2Y462TXeRL42ytla4guDEDJvKwiVxvDVkVzSzHE
yctxo8DN6hvcDrVUEFGni6sMdgACAu8KeWgsGJ99jYByhTg8VZGQSAjgmsjjddAhtuQI0Us5F2KO
+kaOuqh4MS/8/mNxPVvnZDbRBlzLLCL/ttev7SpAziZKSZpicE2KiLoS2twk4RSge3dDZXkel/o3
dwMZzAHZ13IwwJLYIfiTGTBpmH93EwAZ7pg2PRk23dypQMiqMYiCgx+VYT5NZyUKX6Jinrffr5CK
Z63ktzOiSpefODMrw7sSB8VixoZePc7JXLu4oCBAFdpQzt2NxsyleP+A5cQvp8AgJwUTosRjfqm1
IiKe1nDmpPIZYxTu0+j/e9KHN4qSpdMoLgivtcT6lNxaubwmCawVdSsWFlfMlU8KeS92a6ZDXZXt
1GxNnDsNVtAK39+ORNhZ4OTzwE7dxY4rFz68KS2TR+/ORgIi57FxtuwTMY5dc/nqUq/HekMT2cuP
1zi4wDwsVQ1iZ+Tddjlm0bsY0frV/E7HeL/B0AgpbzPnh3ih7mUEi+ValgfkzxR/DiphmToNIxS8
Qb0k5piEOS81K8kjFgXxDA6E+eRlvD2i6HDy55mAvuYuMn8Xf+U8blvIEV+USegFxgbrunDPv8im
G5AwIMTsJFRcvzXb3OxEYCH2stPSKj7O/1BudhhN2nQ0VzeQmffQf/NFrkpaF6rE6Bxu4fhCjiUJ
CRQ1SA7kF8oRrbZcd9rZoGwOoOdEaC/QuI0nCD0QcgNlQgcaGJ6QUtL02q0nFsC17eWVMSC5etmh
zaFcYkw9LqR2mVYNDejIY9bnxgxBE9JwGH3Xy9SyWwfeLSxKK9j4mXL14CNbmP2vp49Sd77Cv0lJ
709mNK7pindk2t0sQFd/uvrWb4OvXX+4HD0HhdZdOCHof4D2w4QIYrgft8nW8hIhPZYvGzbjzdKU
CVh6tHPzu3VJyfXIJfcq1wOmGptcRp+qKbK3aSUVq2pExlifVwLb4x3SEEdsQVm4dUqaG0M4bGZp
VswlCL3imHvtotDwgzwrWUwvtouBbwNsJNSw684T/8UqoQVdrwcrsXwhuG8oNdjQVVQAfqezuefZ
52coX/kdPrg0ec9EROIB/h2OGNjYemzH3oHtuBYQ5K3/UCyz3NSK0Xayecy7iaYLAjOOHl0ri9y/
zdlxdWGUA44Nf9K7+xZlAsQRtMrerk/E0Qosu0Gat6v0lNaUaX04acUGYMJhSFFRWozNwynVlsna
Hw/6vBt43txrAOFxGfBED4VByiKLl1ZaUn9o1NQi2MtEE9PwSrw7JpTVL9gX8X/+1DWpc07OigCc
Hg0qqVpcXBwb1IPZLGJrKKyCwLqxBX9BggvOYLhkf2/6u+OE1Vbg0YAN+tbK5TeScK16h66fg8/V
d6DBraV7jELNSWQufvJ/dlNDnuVRBMxFO+z5SdJCwVrSgWrCKAr8OZZsQG14ZwZs7NxSvGaYXLWH
9USf5omV6VJLkkXXUBDKLOSvPEmhx21hcQ1u9vTn+i7kpPcpv95hEywqld3ozTIqHegbgwf432D2
DhZNO08I378Rla1lMrDGXFJMZ8Db5E4ym4H034QzkqWSPn9um8fw/LmyOhr/FvV6VD4LvRO4nzwt
PtrpdUujpGda2hF2yyhEHRmp/NyNQiFWjyv/3xobqicYKwiroomB422qo37uBzVM3R2fUhywnro4
S5MBt51mAkJZ3uR/mCGjMNZ0qjnrbsh2yOhDEgQtbc2deaJlZGSezWaiSAE5aEotQO0/vK0iu3MP
J1PViV7gUAGcjnQtMFcixpQyKQDntEhcYtA4yIV/TXyp/septgWd5vRNYa9FunFDKY+GBLcWy4AY
v3DVXmXpCe+mZm5nNjsatzRbKf4nwaIWxEaSyDsjP8Di3j5KoEUXNzQqgNM3Nl4Loas+MOQPQjjV
lQPpb4HP9O/ZFdZLbVimKBWIgsIzLwFIWLlUiWxmBk9DxpqQ+mJykj4RQwx6zgnkXJ6MEzuPMgYz
UZFYaZsuJKME76kOxQXokj68e/AWjNb3FFUFf0x5boD7MVCHCSuWMt2Zlb04PI2YH11oUBg7cTVF
TK6ji8iG92EW0pUBqqOPZeTITqkurLuGDPnWgAKVEhKXycFmQbYE750JeKo5NVFie1jgBW5+7neN
2H7BZKP+71P9HaWOeCAaT/9Czy9vG5k+3prML15cL407h/SEz//xMyzyRnQ/eTBsFTSi28EAknB4
EdTI05t3lhxa+CsCq7e/RLZ7fu4VWsFoJWIkVEO/NLuWGA/DWq278liL/Wxe1WFDVXb8jEDLfgps
Vb6vAjrhtVIHG9eqb1vQZeUjfuMK2k2sGHGQqI2bFNLHhXP4UciYNBy4dVQDhXn+cA0o2C7KDb48
rki+U9T8abqQLexNN+nNf/1td8Nnc4xRNvm+WJ8VlrW+KyG6v7TniD/uC8BNujeu2MxMJkOuX4yB
BHbJ64IVCDeYblIeynnkrZ3Um61/wwp52W/QtH8ybrswBA1eCfgs0uuLfN6xtJbw6A6GmARwKBB0
lbkLFdwhAf9iZVbXoPZV6Qfrr5vVsvQP/MupLQ7zpRRhLP5bv/NXwcxamDbWGuNqNxCX7V/iLMuD
AdDI3kiJtMa2i+xOH5TfY5xpdiVvXbjYrb7uZuqlHwwSNbrhJtwMCftC975x3X8H1DrLYi6acKGQ
QkYilLLSkypmZpmiDDoyCII5LsFIQhbENhxHyI8qCS17byAhaHz4VmZ8qRkC98GglmNVwvPOou1f
oCfitnSuangNYAgWUlyAJARk4e62vkbYmEzTSh9cJveNHfhL3/3oSxJMMMK5pfoAiYck7xnM2V8R
pF6LJQBBQyZpr2so90mxuINn/AYhuLdbnFEqc5BdNSaFjavJs5r70Uqe2zxJMsZZREvF04fVrsBb
GuEZ5BKEjxEchAzDXHSu2SqSwsvuoEe5GbT+tnIu3JgG9psd3xre5xt9suJNFfC7L5R5PNku9sLe
fs/fqKkXTRZaJKkFdcXf2QL978biVzWbXUr2xBIuToiEvP5tmKkJUABU0di3VTU1WVLz870wIWri
Jtkqiud2aCvkN+EqzjMdNmdxR2Qb4pKsmWg2BUuoG1xxrgyeoOT4YxBCG8H+8R17YeR3coWXiQ+v
QEePZ5yj3o3s0ff+TtWUqmcRFZDgEwo+Swlnz/jgXNldHKzObqNhFSYWqo1Gqf1zihfpxKYc+8W2
UntruMm1Qs67/4XgIuZGbDed8KGTUKHBgui1+gUV3o5cICqQ3h3+gP5SuNo5vt5DIWNDO5beQxxk
Vkt3OZv4Xo3N9S1fHF5Qv79BnrCR7XMyM72yaL3oZHL04SeNiVfziY082TSrmUjnigVVY2cDIJrZ
HudkXTrlKFc1eAdgCxPEeKeAubjyVa7IlKDtnpna0DkEngSW4jm3w4ucFpqqJ6IX47YCIKfwvaz8
v5wSvDjqfvlMr4818vO2hLIYx7hBu0ak0uFQcY1fl1JvDPQgM7YA9PGiJlDPInQFa70bGe50EfRR
krMbHDK5KhTf/RwxXKw9pFQg43ZR1b2SSVITEYgXh1fYhHK6/TqjQxTs95byKykJlNMv/iDq1zyk
pMdP2XzjMfRfGWLy00OjTRYm3yBAZqJTGCb6s5npztvL6kBsUDo6NE454cd20M3KyZdcuOWEkQbF
jZu/tSvNpSpXF9YCzAKAma5jUg9XhZzlhTn8j1wlIt9EXtSxfU0NNi/3M1bxEI+fZVy3RbeGeMuW
qieJse2QZQLxPdIHvDkV1j15csm3u1Dguv7qIiyBt0dOMONlvqYNLuMtulSh452uC8xxNJOgScSM
RDCepVjc9RDktocylr38VxdR85FW4obXUa8bVzi4jsR0VNkYyiN9TDnkk+aZCR26n4G9NsqLlofc
mzRmFNYxPcE2Oa1CqiT9A4snTZYLtMygwxWEopzHqX5nx4XaPbFwcYtr8P+h8vwQm7sMcXofVfLQ
8DhOS3ly8c+RYjzAiifN/A/fsD7hfVHlY0td4PnSr4PYuy8GOOBUrDO6g4TwBZdTseP4RydJdcqA
Ic8ZNKDyyST6UGFGzL7H/4FZsvISjiSL35pDZlarLO4dnNVxmuaY57MUBPheTKzu5lsu7Sn6YTVS
l9fv8waOEgqSpSA75B7gb0fHG+sezB9nRK5dC1sWVXj1nM1XvxSi3YZkAZO1BUVIDU1wBY42yzAU
QnPvRs8BwklOktfmdHPtFRMQYq/Q0E9NCJtf8SLSobmSMkZzHTrsyL0Gtcf8+/awj4ki4j1Jmn7T
BdyhFsHKiryJ6HYPpV+u33AvBmx00pYdq2xB67zo7cKy2Fjh+0RP64meW8wEnKmVktednjVJ5aSe
nGyggZzkwF8XyJIpVEQ2yfcMUyWFDuU1vKR9b6PQP3d3+ysM3/s//4gRUJ4BHS1DvCwefPuPBk6f
bct1Pb1h+KbZFpdX96R2rTKj8SCfyxx107TM9w3yetB8e1kZg4FPwSNoO3vFjGWMUYZMdGrE12bC
Lh/EkALgqKmc74+vch6dIzFr/RdBqiK7l1O+e6IaYACVq9Qyv3MODS1Az8/QtLNSefooMSuaNg7Y
7Z8ncHnM6uyYmC3YS6ZlK8p6yVby3zgBMlP+3Aoal7ahUSem8IoL+Wobh9mshOAPaFsJCDqhefQb
fgGo+F/Y41HnhKY0nYsvXjlq0BLtxoc+E80VQgSX/tpVar8ecOR7sWBc2UqBikrtm//qYl4CYq4G
1JZM0cP3BkT8I8fXfEppwdkQGksOscbmaqJNAHZj/nt7JLrRdzT0KTDAlYMDnFRkSae9wtKiBbv5
TaqRzbsPfw3xGkq7LS+YUBZT43Cnn9iQDSdLxaZKLixQaMun446JeMQuUp6KzJIVb+GN7tshbSuB
qXJ5VmeQzNPNSPz5tFFmG2rQIw3El5N5pvhvtKkrbIuAcGiFNkdw9BiyEP21eGxHlpZyLmIp4R1u
EQlVXeV7tiLZNrIDR4qXBUy5EQq6Qhj4FmPOaSNOqq4karHYVDuqGJsOSHHxWv6M0Cua+Qh8+16Y
0tx6zkm2I/e2cXqZwwoHCy/f0+j2T+wi1FMA7GJxjmvIElIHigBCVrTnCQ3X7TMQZIhCV9ID3aG5
quR2wJT474A/d7o/Da3Q+cSzLwaiMwAZPHlrGo0fRMU4zAQQqD8ShDqJSDY2etxnpK+XYW1AlDtJ
xuMgviBcj4BZ+uQaPtJm828ngReNJ0r3fiFNzdg8Lr+srbXLdwJy/A5AiOABdDjLiRZMM4iFMiSA
r5DyfC9Et4IELsRbWWMnh/ZB9VywJDMolZV+azErMwhF1eUGt1BZL18v81pc6+CcS8wUq9qoc+jb
xW+ju1pPBQmI5Bzh62DObZQDpW1d5S5vCmkQ0i545FPbIW3JXJqbdyIFGnYM8y1zgSEqNXCAwF5n
AK38kZf6JizcSG6vj1PmKCdxXEWD+3m38K6cDnyw5jzOpvvIpKbeYELaVTJT1A5XEdriWd+qfM1r
zEKDvgDNJpp16sVvTs1D3g9HjmCLbVSAIDozS9K2+Mivszi/9a5m6s8KcMtWRQeAy2PpFEKDBUXa
zM1b8ulI2IJ7OsMBR8sqYtxAI+USNdGcLs1skiYbgk0YQGK6q52ALg1lqBq1e9AgAkhjv0U8T6Yt
P0lmlUo1rUSXfLePQFTDsyfFCiUJhqqZ1A17ioaLBrSBOH1dZDjYHsxEduN/VWTVatVkCrQGUWM+
1ypa1CrVAUTUgyoej2iqJVphDvfLRoTnEXLrr89zPCzCPYEMA5/wsk9D2PLU5QyYItnm8Qh4I7L3
Q2OZT4HVCS2/PIjDEAYM5QCTcfZLpsbsQQvjEXuNEGkxUB1q6GjUdiQecalzmucibsPTaP01052x
qdmMiwhYRCkAy8ytLkImvea4nbD5Ph9OUsHSS9AIO/HVRTct7WSjKnKtQLC1spG5ozzKbJkUI3cj
OfICXJvYHl39VAC8O+xsaXLqL55/zrBdwESrYotDKChdw/zj1fCJH5yqViA9DKf8xzKzbE2wVUx/
xCREzNiQ5kbcKx/z0GyfmYvKhnqtyPHZAfEr/mWaJFp4bTXorOMTBPYVZJ8cIkaNY11gH7LCflt9
Ia7r7AhiJ9i1aHSHidhccWPgFPuDnM2Y24DTF3JXgkUWIAKAjhLHFGp2WYf7TDKfk+moSswlhWtR
51FBLSiJDL1G6dAa27qu4V13rwAPrKvK7Eyv1zdlWp6Nh9UyNN/WqC+1Z8l29n0PZl8ZEegiPSh0
OY9Vc+dj45jn0sWdObumc/gRSMSpmGfvwRRFl6dHyoUCRQwSd6rTyV/qtV8P2m+T2EJ+9SZxwX4K
6ck3lBUuqD82ZK0cqviuoJNpozRh8g3BgcPbDipa9Ud5/2hhgiJApzxrTq4Oe/s2MoCCPfRlcHJb
aemJclfF2NFxKBP371DVy20W7jUcIzaq7cPLwhQJbtBuUzyp6LWj8tQRGgfLw8G4wKVTJYjIKBIm
11fuAZtUn2MwNcOYqKGm+SaN7SGvpvQ4Wmwq67RhV6ghzEyrb2uzNfXqocOtc27bra99lhjemGLy
yC1SW0eVTQ2dqdVr7bo48PaZY6bo+ns1tZt1Gd9bD6JtS2QHNzUvuNl4QMM3Gngy6dDRXORLJQAn
vFxInuqTPapOeFEVlHi2UEldbaNpQqgip4i3pbiuVsqQWYDTtvQDcPQHhoxmNSD8a7fNXsMtL5vq
sQ3Opc+Y4bfPlRnZQDLFv1Pv0rabJjIz21iDq+m0peYt5L+fM19fCXv3UnJhsRs7Yv9t30alPunw
G2y8bqvMcQ2vyLQVzOl++uARcVWFU93+xaU62h09/S1R8ofilqDlMgqvBXJiNe9hUOeDchNKeu4B
u0s1DrFOI7EHJRDEItz77NUKNoUpKnA3rS27cZTSjQbhcb2ZfqFx3ZFm0MuF8oW7TFmWx1w+xHDF
oOPLj0l7fX+J4zonvyhZmE3i4ZuSdVUnNxTxVTO95x54HjK+glISC0hGOl0w4oQQuB0M9uB8OqoN
6wnU7dhBIiqWjXPxHIbsNzYWTHYNKD/j2bCi9IwfvHjAR05mCunr0q8rLmGCgzXe9BsXM/yovA+i
LGqqhV0WJjA30nk5usxkwhPwj9jSsxWUcFbjYpDgH51+knupjey1H0vHh4eJf9qvvnIvoqxezy9g
x67vWTFaogYl55IOVP9loDQEIevPodR1TrV7Uq4f6hkhkj3axI3F8T7EdUgnZTJrOs4M9BbYFmKy
7e56Yp0RMyXqQ3Mh1Y+8QZe2tzQe4JL+KWvMaKx8oMH9sowSJSaf+Wz7u8wVUEafblEsbbXbKZG/
YCFzgytmkzm1fJRIrHBfiURL+240YjDGXbxtC0+Jwc+3LXbbAPCiebEF2EpCrhL6AGVgbDT4LpPH
+AR+PXn8RL4jTi1E83AT2rBetK/vD2RJmmsY6W/pWTPBs2jXlrE1GOV5UlWAh4WCFn4pznIfsGc2
KBtxzsVttPz0aL9qJ9clyMLxovZrh1k5RF5dNQEw1wNYP5INJUHamEMdtLp+FcUlMssS/IGEfFbb
pAXGY8kWF2bUa2cMiGPlB+RIl0eZwDIgL00cXDrvVd9XHcsQ3IcA5pFxcngxCQmgFELTxy5xx7ly
pZsSsbZbcA9fi01DQdEev9I3uCYGZ6veYwDgEg6C6S6PmzXVgEvKaZt8BgQDikAdPSeLMgmMnBFY
/KSsAtfrjPoUVfpUowcYb2dZu2WJF/bCU1rKvO2eGpo/uy8F20rXOKrBk/UxOl63hPxCPzoX3PBb
k1kIlxLvWSW3jlbeVSFeSy6MyDXzsnR2PEu3of60ifnAAOb5nN7qPkJpNsafmvF8DskIqhj/HcX4
D6lAYmTxIsB2s9wyxYjwosjUouEACeIzOuZ5IhbXZDOyTNmBxUIkHC885xMGVYQ1VnmeE4s0klAx
8UszALeOMBBDdl3D6Ptk+T5rpjCPOKN2gOCaaw33F4AYeW2xhfe98wXTlHY8DySp+0ji6DoYFvdW
9X+8gLRMY/EqLXtyhOPCd9kDobubAWvNZHhx45NiyAFaC0Mb2/huPSgVUDTxISgbDIqxa+Bwi0DU
CmGVmo0Ra2rheckitHG5wqS2QUKHUr1+0lMUZ35LSoPj50IJq2gCqLQYPZOi113iuel957OfJzPH
srI/0+MrujOkTslika9z8R628jOVJlHECYXX/KNPQXG0rQjljkpZ7b2ZxYODyDJD3ofdJ3SphUk+
t3jnDIqvJfNwEARuhOk21WkNQe5FUlVWyNGqZDaJvyWrzjOWpxl+7U8Dz2sUOIl9TzBvRTBKhp0Q
nqA4NARKt1pwwqq5w+Oab0vWdrftwIb0TQ3MvOqpu8js7x3DDbOH8BzmgeaCDHIjSH0SugzlNwDx
vXWdmtzLH2YLMRcHeKRc+UTxAihmDKnWyx2sYVkHkaZR3fkpCe9RDIk6NY/lPcr+Qmfno5t+sLXW
fWeUDdSEWfZkLjq/R2gurhgls6Shr1biWZKGWoCoYbX8BssqKJXKE7VsNup1m9S2bmoVAFcnX3Jc
XrXros5mEzKXqFbnTWTsj7v6v2W8EnqEXdrI4EQlFV4a8KfrSe2Xavr/IUeWeuEG9qFvWDWFkd+l
gP6743aTUQ5FS5wDrzbkABDtrsWYKmZ3WJkD106sr+s1kUD8wCTd1rnTLiC8NpX6bi68DCdE7BKB
Yi7yX45cX9+L4qr7Xj3Qoc3VzVFpg6/h5y3wIQiGPYHNNdDHxUg3VUUgsMKnAitpHGZV3+rnZydW
Q3y3yJ1MeXFszL+jrqKe+lLW9edRtk3cuJzDE9lZa+wYuftygAyzCGYUlrM4adOyDBj9skyKY13T
b/vZtoBieyzDDMMwhsTm0lQakg5roHIy22Az+t+cPhTHWlI7H8Yn4OuoaRhhl4yrnMzyTrkyOOAq
cVt9weVXbb1SKscwlMK2G94oSXSF/WFD+MriP1aTXZToPCSBoTXaDK6dsJynMclhQVdk+Z3+8fG0
f09pLS5no9TfLQmTLWvRUyQJL19FhvU3CfGP5/yRYKhofhx7QW0ey+NRSpj2NtI6jEHY72P3sTMV
3e2Y93WnZZOHecbhrnT/XrI8Nm3RjyxjSjcI10Kv+8AqynCfRkRSGQq17Bs1VOWDwIKdcNgG0JDR
Bl8zSb6lkvxj2qyTo46MQpk1huRNiX4gPHBTts3LnvcvRLjjeeD7KhoObawPFLSrNM4wgeCgY8iA
cMNxUjo7HbJtY08144/VCIQTdPIlEkKFItJC+gT5OK6c9fDzAFBmfgtHegrXA2F4z1YcWA3bAFdH
VLltnthiIGvXX8zAyOfkiQzjqgW7pA3VecbXo8WW6AuWqMMe0sxwpEI09/QupqaFPs5Hg81/+Bjk
EEfj9nIepIkQ21doq+2BkoycYVNRG8I6PNwlQULZDyED25KyXXH9VoHihSIY+Anj19TuWJld/j2M
wdpiCaFh1lMX6/EFQs4mA1T2JCiFnw8ObUkIrayczxLvZKKyuE9lVrhy7Twi5g9BsMkpa+Wooc5e
BYeYjMI1/6FXxx66Wkzf1V03GwYngUjDL4Z4f19ITiSh8/lgXWDEVSrh5Yp3XD6sLBFWFj/eRmfw
q6W745dSsDhObo3kRr8xFjioOXh0uBDD4+g7cFAEfMtqubtGMZ/T3lsHDLW/YghonefnpeFg3Evx
ztQqijCErxsmdS227YWumxz4L5iGzx84TjwszNnxUDY5lt5ji1Kevfd/7+jUJ0cVULwt6f9F3mtd
Y+ei9LVq/Q4K49Wv30YN9D3voNYkUlxB3+9QsdP1bKSlLLQEbgi7vr3Kn46pVvcEyxf/6jDEa3Ow
cdYiC3Nk3jqiI3DzOrF/XqrpUPZ29UgE2rYfusIACq2w78IGfPfagPKXzfA26U9ZohEzUVK2HC+c
PpgyCAFTCudonefRj8ztzvd8NR6g8N1IEwGvrp7W0EUVJ37NDlCFBTL6WSkC4Y1BOO2vXcC6SOaO
+8qQ4jTpUCTsdxiU852nbeYFhBKsLiXEXDm96nSKGIifQQ/NU9xLrxySXa6tyKINFenAtec1JU+g
6H4eWHx7sySzOZCcfz5CP8ynOdVCSBcAJD8q1ahN/s6k4NR4F0vvAHWw/8FsiSnqwgE/uWjBLduM
YyPLs1p5MxyH0EdNuX26cBeNinituWdmt/8Wp5w0EsbptqLkHSaJzWphntiZUEdF082FSl9WBGa6
RaECu1vu8gfhlaojwJirQJKcWnyHoypezxTecQbdqlbtSZS0h/j1IfLK4vMydj8XxL0M945HKn2n
srHaF5NfV2IkosmvKI++ipIcouJUMv89YnkJG9bw4d2diQMW6flkRlMUoDWQPv7duAcCTYukqj8/
MTFquy1mOj3rHKHj7ux+V9snWkeDkBM1oJZ5y/7C6bLMk8o+zNtvSc53G86TkjIduwUjZdsq+uha
jU40dheFegfDVd9U6+lHtqTz2IykDtNrRyfQQnuCNaedPA+bl+Yu6Dk89tNsq++a9jL4o2v/URWe
nTj8vvFqVlaWXw4JCCVd/O2XvlAGWKcAVlhaXk2YgspZJsg9SAKNLOViYbF4KUUPWIy++LBezc8v
XlK/n4StPI/aC2rCawNxKyeYaZuAsG/7EMLLzNuHCrifQacqWo1/cbALLjIb1ItL2uAU04p+I6Mm
C9M/H2flNNZ6T4/IDDFrbByehbkPRBmYNN5rDmuZitevT02JqSwC5OfoeKOzvyzU5vyEMSF9os5S
j2IByACi3Rkulw2W25ASDPe7Brj/Yq7LM7giimaW8mglniANumSPUV7rRmHFdDEfObdYOO7So9Og
lXOiMwTNoNsOJpFLwugQ5jEJL1hWuy/AXt5qVgJpoQW/4NhKpSrJIwwIW12KbUcEpwPcEmHSSn1y
tWTw/h6+pB7BQtn1H6rkyhQfU2Sgayb2OdUunDrutjf/kifyx3eWuuGftm4jlA8ISHpHo9mspC81
JPOHUUPVE59q1XBzKSdWjSxjXJXEzv8gHgTc68olbXfSiCkDEBihpottOqFUxTMas0jPbt3pSULC
SB9QXJplFR2BnV5ow1ln957ZdZ64BAZ9G9pVljHDwEtgx02BfZzvdb90WO7kwYllNKJP+h6ps3rt
QjdbGlvDLq+4rJkIFYLUm+PXnnVWk8xiFXS0UV7Xx3orqG9T9GsdT7RPPkNN7nG5ieZrutwUopfd
Kea9mDOml/Wge4iqtyAqV9p27JxjGq1rLN8xMFircYf2np0jk7WeFNsvLkTwXMEccL1VmTZnVU6c
0w/3ILIWd9qBBnjCT599zUCGnyFAj8sfzhoKyy1hOzjRz6PqliUxyUDz4GtcwN4qtCzO7Kqt57IG
ncQD/enVoRwL4goJbbxvaxtUzqTTq+nitQDHGdjevvtZ4d1RhAJJZYjZMWUQwcxkA4oW0/3fao8/
i1wFwogs1SKvRgyeyICelzSE5jjQeM/55Kso/kB5gv6c2/cyo5YV08NXwDlu/EyFw7ShSq+kzjsT
7ESH+3p/DYdEJGXQPjYV3Rz8dymZaOWWVlADLGx25VOvD6ygjvnF51JtKbn+0NtCVStTwyREVuWU
25Jm0gAFFFUcvy5nYvVY9+D11GQP66Blk/69Ai2e9cSSywkeV6OaZ454BRlun/8dhRTRwzy7Z1J5
aFXjkmX5dnWd8TkqruOaLWswjZioiadNTX/30D0Su9tWUpLVc+5iyXm17owfPv6+PW/7Tbv1lWhd
hY4ImMJoKYxDV2nJ4Q8jEZP3XKpsXkqhBpaB6jvgwEbJCbBWnClmGazaa/+JFQe3CxBJJe/6HNJU
IKjrY3Old0d+GoGXiWuTufrpLY8XUKYNj1W/0A84q3t0XGSZbFb4aufaug26k3leXb49CJpmbQuJ
PIexQr/MjsWVSjsH25GkAhQuE2AUtfD+dj9YXImVFCRhJHXCMCHudf3zBy33znrIWNdJi6aSStIH
cPSGsuYUi1YMHxlPXHmssAGQWSJIxjoCrnopEqkfwHsOkd5ymvX/2ZJxScnjlT+RfSGWWAIla08T
EbtltN92BNJwhhQdPS4H9fq9qMCt5w1o9pkc169f5dPc0OpOTicuoQLOoOAxixedixzkrViGtWM1
x4wXAy5YCQqhqJootQ6aa3BVgAf7UxHMgvwQ9uVf6GI6/5KNZzIMVAi0hs5HGCQglAGyPmsowDSE
cZ26305nyMl57BMAWj/pRXAWceF3Xcnf1A9ByIQrYDaHkaMbAwDd8xaH2JavOaBW/iZGDE72zvmd
90pMoJG0ctkO/BcsMnv6XHhln7IJHqi8rqZJWqsZwwuZfRvBOs5xI87UaumT4DA4FJ5lbluNEyiN
sCvbkAsSJITKNEOw6dfmq83P2U9sShnBhxRClisQaoUCzoj2x7x5YvYH/QNyimx4AM4g8gsqj2nD
79hGqmISLL5geLmeHJire66LXu27wbN36RGpvAEqDC2jeTlw0832as0k3elKoRGExIqQEn/sUjDE
kfjhb2onPEpC+Laknyae5rk83gmHrIkydL6hR5A7H7DWPLClvtGUKT4UnFR24hUt6Xvf31e7v6Iu
f7b5asKcQ1tMwY5vFr3l17faPaqw+S7P+jQi7sp5c8hgZK2IDsvaRIfQAZDV4UbHTRvnuvND7A5K
YAyLDi7NkPUlHG7HSTi6zjlHZ+bukMCDrPVX7PCT6IB1iKTj/8YxxfQvsGSZmQTzcwmRzjn7m44D
er8LMVzcLNhnmSJ4xDeD6GNeOOKvAEUYIhclPm+J/GT2hwX2xCVWV3wLhWmAV+05RwNtFmydIklG
MsPTl2wZNro+sGRwBh1qr7QwG6r2/mGj85jB2MWqZhqmPT+faa4RKe2aJs075iIHFk2CTnREjxhB
ZTa9UybUtNUiE79I4SC27inscJ2pwCfCkmPk1FC52+cHky4YAkdNoA4bTMxPAcUKa46sZ4mqEMrG
l/084k4DGbPsCmdaHiEZZ79L98e2oJa0MVosP8nUtlUO84H1GhSaOl8iEXHqQ9DkBlBe0BAWMs+t
RBLP1U5iCR40q1zdXwdSeiSCpK/JD7Yakr/EruW8OstrrdEBygfepg/7MeOUaJeJKSM3wyA7CSQb
A2lsmy1qGpRxZ8InDIDlxd9S7+Zge/NMDreKO0ECQ0Q/h7qm8UI4Hos4XmWrZfG7VYsiEwR6GDoo
sYiWfmwWacqvjp4Vtg/ILr9JLOv1ps/sqMvEdXI82FnPkyk6dMWNBKmRK3DpmESw1tvvcaqQZFeG
C8RB+m1V5HqSpXqkKaPhkhZjgkaudRjCKPsmdEkO6PiA7JNdAEQ7W9Yym69YvP1RQKyVU7HL03C5
1fZbukQFR86Aw++865FCJnZNiuRSGu8qKOaDQpPK3qHx4/swWVSaNNsoPH7sXDsSTN6TlM88DlIp
34j0rWsaFC9nigYfBiPOe5niQPNRNdHd7WrkWdVSug4ovlul0HM8odqUvSCqSuyZ6ZaT8nAxn8Gl
UMSFqIMm4y5GC/0HhO+WEmrsn30eeskK9OR06oRwz36sHhAYV8xO+JPNe/E5qjarOy/l53N47wDV
aPSiWRc/+oUmUpBEr2Kx0BmTTHA5PsCfkoxPqtUbJ1IGbbeKG8A9U+nvKmcn4cSlrjzMss/Qt7cf
WyRrfGVvBsE8OqTF4qLsk5iIjIKan56Y7giUHf0g193CpxenSeN9FiZJG94AHgIT9VdXjy2KA8ku
s5gGwDfbW2B5eDq1zoQ/uNFsKIkDGarJZrg92dW5BSNZw9glGQtSUKy0pbxhnBoe1eDXSI312TyV
6qfN8Wctt+g/2RSQ2RmJxAeKQ75VZOK9XbalYqs/w56bWN54TVI4R8XpehlK3Jh2KkI8GYQBuklQ
KMzwXozLpDZGngee+OMyjnxiGqaa+BGaIAWby5iiLAYm+h3re7HTsnNqhE5Fg0+OHZgED+usysmZ
Vpop4Glo9eV+kcjyQYrpOmAo1Tanch9pb4ib7S/8Hz5Ot9w+jRKtD2eCC8Nxs2mN9quqkQmTZWRa
hPDMSU5XQloRFDxRAaxZgzk+TEWu9YDhkiNbEGSyBrrmoQkHhqQO4EaARjWCgTCOrbVxKm3srjPn
f66pYWTHjphoq5hCBBoG6rA979rDB1GZG2nbQ6mouXN06Pxh/188JYzhgXV7Qg6Qa6uqCSaQA/XW
9Xgpb8RQINvr8ly2G1UnNR6o0JrxBHSpa116fNIoa+1GIeqB7yZXDqXblttkZxrW/y+a/whmUJQl
EFmVRzjQ9ytN1sJkm2ksyIg8N950mr0faTURKDRjZJ1lEMoFNSZYaQMNhOXPPYCKicH7t1GiloIP
4YOvoFXxq+BbmbmLgdSQ5RfjlpGnHt83zOoSff7exF4fMx5LeCKLVlBess286qZgkblj1KD8ybH+
90NWWoZMWBwmQ0wN8Tbky2mJLgvMaxWGHIAorXlrEe5eFe+Oz2RM1XHZ7szMFTBH/Je+wujdA5AO
Hla/2MW1XZSbscCNYYHfshyVOQSLco2Ev99cSZ4pr1OItky44G8xTNcIYa2rfw0xxJAkDOTg8mth
y3sgc42jQ/IuI5CC9KTyvdL3hSQWPDo3hVJ+yve5mf3dN1Vnqj/nZ55omP30GjyLC6Znpt7iwbGa
UW1ZuIWaRDWV8GxH+h2oxx8zenmCCOndtkY+2scAum/0pW4Z+bHvsY0vKXquqr4WxjGmd3xXMVMl
XCekGcanCwt9wSdlDY1pUUVZZcJyyfpneUr3BGu2pfiKdSeaPYGL588vAtA9DGLlcRhuTCLtr6SV
JzVyf8yazdoOtNSi9jX+aJ8N7NdiAUqVmcPHKiO7FbGJuCR4jEbh4dw7aPwUuEd/j0D60Y96bpvA
xNPtKqATGVubIfZuGaSzpd8CCJBFoFkIPQGKkVS3XbP1VFm0s/PBv3hEnYHmdChysmf+UFrsIM1M
dcroI76QSILQHQ3d7gOXaDnSaAsMGTAhBVkltAQd96uFENDTQ200qBj65d047fDWhBVe0QsHPjwV
aY9GHTuSgTuURMyWsV4O4q9F4qzMGUBF/VbBCN4eZg6sD99A/z+VBGwvUqE8OV2gSRZ2CgppbZw9
1VOLEfiLPHzYKKsEweUDUgIFkf73GgtPPMM4CMARz8pMN2Wvn20Gvz0OObYj+9Rsv0h/oqaFirEy
Vbu2pqj7tOvU52gKCqIcTxAkQT7yBqAesOG0kn/kDtObBP0ohrDuhrr0VXO6L/FrOB/KdmQ2DHOK
9n1qMMgwj8pWjKaNVLvxEYxBW38ZX6emBa11JItEyT1LHlXkM1NI5Oji9EYxuyuu125VZscEI3hW
Im663WjNhAIAqSjV7nnDh/QWk3v6QPZMHbzUiRc1ZFsqNfReInXqy5lZbkxIeRVtBwP81NtHvvtR
9y28jCzBLbvJCIOzA+xsExk7DXY8B+HuiVi2vyQzd3N4bNnUck9SVFB3sPq+QcrpoQGh4fZU4Q6Q
pa12i7Ba5lkRJ0syM6wZ22dKtFu/4tHgy7NA7fBgO/VKhGlOpqndwnaEVMwYTAVvC/4zfCePp7to
A78DIsuUagw5O0PCqrFLY7kpdcTvVU+xFpfBp6xJgXpiu28dFkibat0rKOPe5nzPB/jB1t3tmmPU
w9uLTGj37e8fMENrNv8YrSK1GwzFe2NyEVl1XmsyydbcpMXReBS52aMqlBYYJPrLZ08jCZ6DtuPz
RzSh4plni10OmF9AzIVgqJWhnk3ZLbAx+ocJC/15QLRbn/WEt00mZ57RdHmk74iYb1n37MS9sLmk
Vn6Zu2iTJPlJ1/llRJqMSm/Vy/gmyPMMv8olD0eNG3ORAtdw+ExV7GQEGW14Vn2SDFTVvSCdq0pI
tSXVx2NEV9EHdyEtkYV318GI/oQaNGAoUiwQvpYVnMM/jiT+T8a8B30HYmjnYihB3ub2WqwsbUP9
9ZZHtZ2kwa++etpt79dR6/lL5dc05dkMm2ev4JejpQF9dBcHV15BBeaNY8d/wenLZ5iUn4Gv8NaF
FFqLc64DSK2wcHmonjK2f3IekXN8b5B0UlAawkPLRsie82g3I9aQ42ywgbJbKjfV/0nYt54mVIco
e/B1IENgSHBbdzItc/aim0foJNlcxEjulGh7m8tsvG2uRjQmFXwGCxQo47RKbV6p8qO7HjsrwNr9
h5LRK5TOABYgF5EUqyG/Qe4mjx2MrQ4S8pUkgGcce0RhhV/ItopGPDmnulOlSu/Br/Fiu/ig8jZ3
vG/nHL7HaFg4LBTDn5cduhdwXZ8IPF1RFx91IgbYsW6/aAYzqr6+Rx9nzrJ1oo5cAdtPxqunqkhQ
tFBDKA4hmBqP6fFhT5CXFF3fgF2dIL4qFEhsySdIR64wabkCS/S3q4BLNEHtPvonU45NgIBkVY0Z
UqpXT0h+20tzkhJeFa/qF/IccgDt3PxDxbM22E0mU4VhlTXcOVtnfXht0MOHNjfKCGJg9R65tENN
Bb74TJpLcJ6xh6FB41LwD5hYzXQSOuoEy4tiuGeoDp5GcnWp/D+cnM7aVgW7bQfDEECM3NqM9u46
d/73IkouDMSNYgijCf26lIWUOfJX6O+HmlmvHDJwrZkVQTmZXePksF1AH+fU/Cp5u1xAUjMVVKG0
9dC8xbaAmbUrPFjGHj7AqlPfdIZ3fx1WUvDbABbJ4Zq/yNxKT3Oc7LYaBxX642dzUadUK1u38VFH
IyAqKgW5NqSsvlb91DXTha5SsLnbLsVvYmdMmG5IwZUMlS5B0KtSymwylPALL/8BvY3y09k4jCjp
PrGILB2kTKmfwgE4y6Nwa/2NfotdTrkgrCsDGNCNP5AYt1gGT7B9wbE4YHNNJ/IUjI2BY6FVa1h8
KV8Gcp+Cb00HPkmJ8PaXB+jNpu0TTVCO0bwf7Z93NlgIAkY1TAtyCK0lWrTr5y2KydfxP3qG5AmB
ktK0vNn60m/UZbNWFgC1g6zAI/VmPkw3pizIZHvgT3zaWW8TA+pcJ5xD1gAA9ecy2zuJwaczJBGg
patlj0XnerMpYLPI/l5Npv8jgDaRgApcV3hQLSXg91DyK8dJVfL04t2IWCb7l4cA+3y+W+TOihAh
cVNCYSemoMKL8MGxJVxiTR8Cn6aoNevvnZKbEpEfh55a7zv4gMGNMDEZzr+XYHCL4BEC48GwIh4q
PkQIdxSCYAZzvyGmRNUNjJxNTg6//SODs6roDr8n7qq7NMRvSrpkaucOva7XuZ3zV2aEDwcxQSdq
ifCNwAxIASpnBLJmeGJzEZCrG2Mj8OZZ2kcnBgyG5YtkkSCRe4st9HPz/TEfD7pb4V82eZqaAKsm
b6JjtMe/b+10ajmSTMJKgVs5OvfC43P2XVRWfS1aLCDIelL0a/8+XE3Dp8VEb9wDUTgKaG2HZoFD
9LXDdr+DVHw9jcrXVJicddzPo/AYZPTzETyseK54LRGLtrWjdUyqI0cFTYBh1McRVCKAre7yALNS
z0hd4RaeXlWtPjVhN/G4XahFIyXM7Z7T0d6UewRAtgeR48kz6mbI0/qtUet9FhBtuYOkbvWqLTAE
SphMUgOkt9a/2cMp+dSEXir9VqWQpSqkzk4XZJkdALUEy38S2P/9V/H6xZQa1QmN+D91WBU++EXt
J19XTX1qWQ9erb6AS6+vCKTYKsQdT9XjnRKqgUcNMMNu65kzbdrsWp0AR5JxkZ9jb4iBoE1X1Qgn
2jR3ZnybaGdUkRQuILkJctSTSrZBhVVMVXhYud9TrTCdBjamJqhpcSiAok+2VqnCwTjeR7Mx5NHy
xYjoxKWEW7i2oTg9mjdnoFlbgK1A9gwUjkL8iP9tbmNFk4b6w5/ViDEDcHVTfdEsP/uofY66L+3f
j6zSMlpl4UpUKhsjrHRi8B3MnNr+ZFvcHn6z5OYNFXMr6psM0UPNY3opfes39YVA+gy6/Z3mG/Qa
Fw5s6z1xKO+VyZvZiRtwLo6JTEr8L7o9T2tadZn746LJysxjCJG3nV9g4meFvABWJjNJVeuoTd/K
UXNxxSfZ4HRK2cgv+fWE2P4SrKJld790aeKmnV1zMSWILl0n4vNgYz1whHGyebH9xNTL1m8cymkf
dLwFuLB5rqadthiCw6Ej1hiS8rfIiCDdY2W18taT4bO2lSwozWcY+rmee3C1IJtFknWFfLmYF9+z
mDKCBFT6UJYS63OBUQE7Pe0BD2guRuoLN3LoqKhvWaTBNYwQQbHp/R3eNRwt3zew8Am4oOVEenL1
NoMX8fAX/JfIhKX5g+S0l7BHMABcnDFpSrjx0yWpDC+oc2yIKtuQkGB7T3RtcSGj/QSbYZ2o2vCe
EJtYzbsau0H23o5ScwiMvLN9o6DxTpXLS+hQlPfrBHRrZYmpfft3YxzPF93977II4txMese4077M
3LHCdpL3M7CL5fTkg7K5sfgwoxtiuUQrS8VVGoswiF5HCMMDWlE8CDpkWsCUaCiuUxZZtdxmaCt7
+uAyDkE16gPbm4OfGjczIjVUB4bXJzV48mIVD6foMtKHfW0u6b/Df7UKkxeeyWYMlvNZ9doAcUH3
+MpF9fOh8tYysjO6ycuvl8cLeg0UM9jNJbJu0zvgi0TEVorLAOKyR/U9PqfXQo7syRuEembF+Nlo
rqf0TJLOG0avHJRHgqUDUdZL4bbLIcPo7zUIv+x4gVu2L6f1+CoTl0t5OkCG4vHzpx+uD85g5G0i
D4E2lBx7vSUveuRX9T8nGrNZrdgOjSmKjdA7Szr+s8XgTixVVpWa+OMfBO4smxbVMGwq1Zqg6T+z
II5cLpnWWQYl3yWefM2ydbwkqNaMNxH4JAGI//4H8364cLh5Pc9JJILnRobXbO6XPJ5VYQgpDXru
dLav76pKn7z0KuqZ3Ystq6BbLbOHckV/z+lEzIpjQ0H82x4HR2BPi0kTMytI+uMvsBZ/0ipb0oZg
HHOpo7SGGdPEP0SW4fRHWWWNd9p5/3tQJZ/rwYMKlcpqNIcjsCZ0OndwsW6nagOx4YsLAXy2a/4W
SBBcjs3e5jcO+IJ/G5/6MjuvrJQsmDEDjGo/W2p5HWLdwG+kU0CEFwghGRsw4UbgJlNTJpLG0QHa
Y7/346HkrLIXedzS57+rt9ljLTdLAkQHLldFwarF9hpCbufwRZGCN64Gvb4/FgmsCBCdBF5Be/mm
WOzTP9AcfgGJpS8giiQaDeCJaxFg3BYSE3fxlF5DJL3TBRpXAbN2CpoIMhHeTdQc6TD+VM8PbrOY
uim6k0mdm8hXNimi+KLe48r7i/ixF/3ySMZu9XhGBh3ku+m+4bAWIi9p7vZn106o8hFPmLtW7O8i
Jd6+lOFODtWj9D5dULZsXo86Vuo4FXzfX0dJ3C0zxfDabfxEUHagXoj/nDi/6nrrY8YIS7alttH1
Cl/mfwO4fQhJE0a5BCDrsPgZHjYKJW3SgEI3RdaWNCTWPSUrMshnlAQhm7SFhjl2UQbYJJXjQGmA
8eEdyJ6w68MmCDUeMN04FODknxntxZrWah55dZB6kLNZltNgnQas0s36pVxTQu3FnkO9OosfDMH6
21/i8ZA+CrjzXYm3H6DiuFB6mNzEhO0sgg+lpXYOzgHCHfE2tf5xUVS6N+SKOMnjP/jSizkKHwpl
XofI2fbCZ+0nIIRzBenWHcB9gdmlAsZMdNyeuJUAH8LmyzNDu4y90R19rv8RVTsNTUc2lHEF1LzG
X9wSHrfJ0NnC/QZI+mmo9f/LOx76fwxv0523lB1vds896h4dN/dz/foOSUWEQ9KevbHK+8V9DlKv
AcwARCh7gJ+4uRTu0eOcdsC9Bnt82zxoccNYNhJJOtrt6oPt+tHnd4CAzOWdVRr1s0xlDyHyd5IY
xUwrZLRExEdmtKBSRV8jBS94Z/CFHGQjnY1016SkR4cuEVcjKD9iokb5hktm7N3wYJANJODTBP0h
Du7p1+O9ojrbuylLglZscYTe5bFmLLQB51Waqw4CyTOLBanhBpg2MiXUmNMNoSiSLtG62JGzUsdR
v2x6NsUShsncBxx6C+RHkNZdHWSe4J3ztWrdYoHAHtZywjmEqqpkZApprt6r3RO0KMWFpirDOsIR
A4WC/apZ/7NQYoGWc/odLn9jcNSdNyKM/E9+IDLHwI5yw3jjhRMUgtd+9LEyIGS5fYgLTawiY46R
FuKU4PD0yLQUoaEVASe9kFL91QpNnGSz/UL4hiPNyFhmPyJNh8mEvZFDxAaTME6iSuFAjfCygbL/
3HfVtoJnKU+Hvl09LhuqNgosLx65GJoYreK3OA9IP6m6Kob3WP4sJRSLYdxZqWSBeVgQs81KEh93
QQWuE/CyC0xPaZnF6MTO8VpUG3+XZX2QIrfG+5hwsyvO523jdYGYn6E1KBXIExWu9L6A5QnovqQ9
hJ6C/dr9sh0QX1s767/d2KESzpNVi7DnEKJx1P+13kl2wvWBYmBgk4r/1y05Kbsg/AU560hg0Slb
yAkmIQ6SBJOKAr5fIL/t3vszBYv3LCLxH/TGk8kiTnd4WwdPBzrA5GG1LYnFGhZ5o8pTmYuUsomu
mcZ1ZDJDS2PZJhkqbuY0hvy2M1RF90Ud0KyDjwmwnYOdOcxlcQGF84a5ymxj05yMWQ7Qy3Z5LoX4
/zw5HohsRLcCFd5eJhC+WjERK9aBKlY3zPpR0m6JtQclBhOxb+3L5JAIHCWyKdbyFj7Nwi2+gnHt
6wKeDRFd1BSRxbTs1rN4CZt513rTiuZWEQoUwFLRZU4LL54QDZejGpEeNGQKQbfR65T5GykVlJuO
/33snurRX3s+ZfwtAFR06EVgZkABg897EAS2cn419Z9ioDKN7irVInY9UjWHJ5c8C1ty8b4FdbN3
WjqPR+HFKtuH3rsrTbXeW4C6Y8Lx0lP0fieKzrzzP7Arhm64Nesaf/Xfry9Zy40ISkpRNRztfbUa
a9xn9e5flhHXj5kPdfnbcYBnG/xqKwUQwS9PMBW4JxwC8/gkOXsBgYfuZboJPYaEknY8Iggh8KFc
oC28/u/EMijG9tdU4ZwCWJ1PkR+6VMdk0S7E2RX/x+nAbSAbRfzFxtN1u6mmBR1V2F0ddXJ5KuHw
ZL4+6seZlbZk6R/l/msuGenRysUXrvBBOL0z8qp0oTg7UkvrqHw6OOpBMMBBIU7zKc8Cx1IRThrW
iZF+oTu1iCRQIIJBLy73U2jEMSVJrn7/xKmkCUGRkNyaAhYpyacdjnW+QR1tFraerU+CBgBwTn2R
wjfRKrpHHBgxWBJqDpgttOX4Cv9QaMAF6YmmwwxYXbDJDZCO3kmF4lHNobZIPOM86pagROrP72eH
yazVH2IjzUBhLrfBJAzeLIUkOmyXwOE/Uz41fLrMTZ5mJqWGO1SOMta56wE4FuH924ybgj0b97Pf
cVegkgKFHynyf7KU4dTfYIqAKb10v2w8ANMSbDWQgqOLkXELEbiHv90l0CZHvmC+A2L5YBvYw9hl
pmNLV0CcvkopIHKYjfHiV3nsV5WOtHJ9wwp0vgTwCxD0IglTuNe8wbx8TtL0lfihzbfnY/bJ7rCS
tXFfte48RApJEoI/99hqfU2Z2f9lsBBZILPnkG7fMBrJ+vNmJH7bC8fkT9z2yc3uVhDy1R4G/VAL
osGCSTShSgS3tvVMy3OpJGiFklv95k6/V87OPVUM1dfWTJmijrefaEkLDgCuTDbG4EnBA7c/HZJN
9sp9tAcKR6CABlntz05SxQI2erLjrVlUOrdwnPRaGNubs6QS4qjjkeafOTcfNwgqqPAqu6fxbRse
aTB+8galiGheWrrlCIuVTexGE0o9hDbqUEA+Lbb8E75/k6QBJM6l3b7ot44MGrgvawNDUKI1vsPm
P8obPmgcYGl5as7YBJLFB/NsnviGUthbcFnTd7RG1o1JqdsLN1ytmYWC8sykE9Gcni5xxWIytBM0
znkFUNgYmGPzQLBxTyeydSrG5k/plhrkyzxb9QjM1mBpDQI4r/19fpn8DqBtEbUoIQsZMZBkpUgc
NCq7r4HxXF0sf9rA5x4vM3Zk0xtmXh6g2iU1fA/2VqV6Bes+QsMQKmz6uLrNKVqo/Rw25AEbryuR
jO0EPUgrVIs+nH3BlREVlkXnU+jUH+0rUjit5BDFHEMr8w8M8AeRsxr4Dj8dkHYi9tKuHKl0uTYV
prQVVwfmcmYREMnzCR2P4d2GZz82w/87gvRFp9qpvBgHkWY8SyknurWXctU/ZkPb1Oz4+TUxm05X
BH/mM91HNZtDchxlAKyvBhzbQw3e1fiCltbHMsOcGnmNeiiNuOU/uoV5MKCqSJoS3WpR9E+hVOPu
CS5jwakWgAsgPyv6oM+apmuoeORy7vMJ0igBWpMybRV1aga9TP7OtvGibbteNQnX4oQzqj7g8Kck
90glvz3tF9VDhoGC9mQC0twXoRWWvLNme+iA0B2t7JjiP1EZ3WuSSnev8vnzkCReZkT3rtKOdf5s
n8/ulUYwJAh7MOMNfUh+tJoAu7Jpe/EVhXak/vqqs9zgeIDsK2xiscNvUvvZ46KJvC1OSRu20p6A
Up636sr73dS8t8oRh/55SSteeg9Tm3XEF7vV8aRMOPlrXU4oYwGBvnwmLQr0bZkJCepWvLl+okCm
xnEMY/oCpSciRRi2i8FVG3ydt9/njzB4O020zSdW7f1qgCv5mrg/2uvk1nAql/DHGt72BZMHGfbr
OiIxvorNMXOnPYD8jRf+ifs348l3fYpB2ab1ejD38f/WCh7LISKEzyF+hgrojUzPJ03YhBa29q86
fya9pft9JhW63R5ZsqwXVw6uaIjIWww3EjW1rI422tya0bB/S55NWVrltxrBUBQcn46nT5ACwo14
MakUG5Ay0NHNSUwtvjcCXuU6qjvqVHdtBbHhXsaj1GWO4/I5gAdSSMJ2q/3eteLSqsaYzwQVJMD+
3zK5eyb7cuAYyOJjFuOJcx65znFh/wdnbndFRkQtX5EYLSHaDtEzbiBI+WQrf1WpxYzdlQ4hedeY
jLZlTpyLqFufX9EuXUpDoB/HJV5EXxc21e1rFzBVrosR7Y0uDNLi2OAxsmLCcU90Fsihrs4L4h5X
hH5Cj/qkl9wyT0Y2XyCDxr+pH5oogynUnAhaUYVhfm/VWpiN8Kiu+cMcjDKOxFBkZPREfz+QUq1u
o4mzpTmZrH/D8M7Rn2Vq634cQkiiBxPGd3c5atw7gl4m+VsPKpLP5xZHzGgqkzZlWVEXbRwMPeFl
6qsk8ASKj4ZsWogKONJaoAJ6TTNxXK8P7koWEZDhT0piPXCjtAP3jReVQgDW4bNg0QGGte/vU4Cr
k60s94qTRXWZa+Jeo7XVCWVcnrj1wd9RA4Q3I7QvnfE5ciOyhRsLuTXaTOBX6y4Ll7YjtjhMxLgR
rrUhjlhkg1l00V/AIHu+I6+vsPx8uLAhojfoCSw+Snanf2f2u0a6Lp+rjaJm10IlcVqDTCtUJdcp
Kqm0yr+dxASc1wko23vmxBYzVQEYA2F+uGFDT0KFkorJ0gn20sBLi4WFi/sAycvCoTpBiiQB2iMR
U08Awm3vi38VtmAKlz8gSkEHiOotqFv2AZ1niLqIh9oaECPAV13yMbK1Dh1TmjX7rS/iy0nmd/2z
pgo60ycA2tu3J4a8MedBVEV0hA1FaO5p2p8OrPmRz4/gIGiIsFOwbrhpraV0+KhTnXS6O1IEJCbz
tzfvSNJztnff+uD9ox9CzfZ7mP8i5APo8ZqcvvXS/bhcWWMQyBg0tGm6dD68YjEzQ1M7epSqBz9G
OGtWHJn4siC0u3W7i4s17ydOczy0HS9rMdI5+wBOQk+gQObMlJOjbDCDWRJ81xHGRoJn6QzcFtKp
4KogXMvIEaUnSD5DiWsw9pdxZG0xpUP0evV6QFqeR+ybU9IxAYJA3fdcOT7ArPzfuJZWqnyJsCSs
1/QzmM5AoKfiJfloA3EJtR5azrExtIdan/kwXqsY2RLES+ld/TWm7eXLoSV5/rhFP6GkjMrpZeB6
LyCFGQuTAMjp/mV+yIWJa1MqHRL6XSMWkcy9CphO0YmMTSsAAXP+PBcBMm7Nd5Z/8uV/AKIuoKAR
efRgkXk3uSK57IgH9PyH0hQim/fUj7D9TV+xuBo2OuEoZBqDu3wWYCVBq+QreEU08BQyKDhI4Kh/
sI33fVu4qXkcAt3yhevfqcLQmW7yBuj1LUV+7rs9U6wqcdPy5ey1MTJzGqfr8/Fu6MAfeBRVG5gP
MYCjYkm+d6ay6JnahH10UvQpcJRLQpd6vqXkcAt6pFdNCExTR/eiJL0Es3/lKPCjGFumZmAN1ETa
hec/gFSTaARpc9PxxJp/l3LUmdm3ir2mvFDckDY984APXnBHrY439btjP7TXI13Eyh34C24tPIjh
Rz2K6DX0vv/wjmPTyshAefhrOs7qRNC8lWnBe2WCU+OzQQflsO5z9SsyrciCNiIVsb3cFHY1J/b1
Z6PKTWwZxtD87hnOQ0Aj9wDgaifvmq0wxb0Msd0BW4bh87tcnJiWW/V2AiZmarLQKNV4X6AP8me4
SPm5sxSt/VFgXSbFoo2tLUch0ktEi92xhXTmXyxpt+CTf8CTO6m99HiIZ49xNt+9LyfXrH1p9dlE
/R8FpU7qe733c4Sh5Jf3kuQ2E0gx8F108YdjShL+VxhMkiSJZIDxgk3asKIqRC1Xisu0PJzHB+S/
RSf93gRfMS8XQN6lc6v9dr/Snn7xv67u/G8uYQOz6cwFueR/6aha8vwhZfhbfJYqc9I6jIuFOlYC
VNKhRkkfriJQBobyEtBmMZuNggPxjDM+rItac5Bsj9HANu2wCYT3eWTc36tNWNzPAuK/FYcgycgL
Gp6yovHo3AcMIbajEuQNQMID2E1kJXPEzQWnzn8yCWFM/jwL5z6EqnSCYb6YbnaSN/1JKNXmaIOs
2AxJAV9kQ7kUCxkPadBiTBnV8CwkBwKpQGkCm+8kJPKQH67jhqy1IeK/Gi12B2px++gypess/Noy
9hsmYsfq//P6Vylg+cAKM2gXvGgtIyj6Kl7RFQURe8o4K+M5WqE1JW0usUU6umhH0Xj82FHs/fC5
c32Rcza61HE4N25l1ep+dnm2+awcjtmKIC4uVIoxC5vNjqGz8c1Gxy6IDx0E48QBrZFTqCPf2Bpj
Ll+vwjJD2D0+uoJoqYwQmPw0Hc7soz8WNOYTE37qJg0HKxkUE5TYwz/EmKd6hzBAwm2yMltLK2QE
E/3VkwlR/U9DsvGwooFpS5qYQP4IdIZ47qcJT70VF+9H1F2/ZDsLSHwivOjG9rW3gmzATfxiA/YI
ESwbQSq8lJlRNxU9/mRIl3JtFhZLMZ8G065g1hbAtxVmyLm+CD0DWENP5yMR3PWW5YgCu9ViD+fK
GaZenzdaCmYWik0yD+2Dz8ST6LD9buZ7h/+AivQV2OAEcacH+5rirntBU0v42MB/4DB7eYHD+aSj
IwgK65V0d6vfb4c4IOpsJOC3H/KGf8BaP9KDBQzeA4+ZW/zuqNptLgKY/d4ghynKq/+5WDN9Q4M5
YyJRbJAb9ednce3vH31Z/0cuYf2b2Mu5prIFDkhaH/5rxUhI8bU5O78TKnQsPxsEtOTBAPMFce77
GIDZiA4uUtVxglrW/j93vIEFXAqXzTw//s7Tj9AmqRKleD9xzOrDIQfzB/htrXrsTsfWHPSUmE29
zcuJkb4BOWw++r4IS7ngaKBRLr0i2qEt2PTQGmzhhvGAZKvT/Os446fZ/hO7rWrwlbVLDerI74uf
e5akC/58Nmjl9jzw9kNup8LNkXKw3750dbqc8zxw6RKw1FVDKQgT2InzV4WhP0ziFm4rBWdIguGK
d3fLt3P6xtZVJ60BlrmDOsBLVfP+q7+EIB+OtZiOexkxGUalOHhkvT9uW1LhXWcK2QSYagYhkNHR
/sUu2LExP1AD7LRNdYd1f5mKHXMsqP3qQQAhIX8tdRUtPNjvwfefuVBQBhl7A+G82YPek4xSeNOx
XL/sz6uSnV+gXDVztOXnyHVTS2NKLE1u0U7aUptyYn5flQmmRwfHAdmdNYg1BFs8GYg3D35h7Ju5
VIp8lnRUMmZNZqqT6nxlEImb1jARnYKODt7teWs0ia5o0Nny2HbD9sRn+W3Eyiaz5nWYbO4j5166
QifUGJz1VGkQ/3FUwZM9rN75Qqh4MYNfDRW55fmTeRt8pP1Ukr10S+KIOpz5hbWZ7Xwk9o1pc9Nf
BfHSA+knC9HaHNKTdCQBO4Vt3AsVwdiLi4N/T3RTbGgRHTZ/5Vlg/RqLp0WwPcnm6SIYLTy9sopl
W0tpp0sm0xwBnYrJySc95bLpSIJyXyDPzjzUoWnzHeULVXplfOcmc0WMpwBZJPoPs2Cvilvul7Ir
om9uwmvEn898EexHeowG5iTaWL868fbCOGYc5Sh0sjZYDR08WYTQ6K4tbc1Ecv8vIPQqDD+hEHi5
vOJV15FHKvzpU9tX4WP1JcxhqujIAEJT6VPjrz7OvDHi+GsBYjj3jrJSNF1ELVH/IjFhxkwz6k/6
8Ai0QPVoIm/Bqxby1gjsR6Idea3oMsfLLwG4tNjYufNtoiq3L0hLCPRj5t8vp4vJDoatIDLquLZh
hGDs6t4baWVebkzFHlfgvtmbL3479pHMYZRiFkMlxV/iDrTy/IB4s7HPA0XKMuFZ/XAOmJhmFnSA
taxR10aKeo+VUPX5aMbGzq0+BfBH7/mpP/4bj9Jw6aSv+QA29HumlxGtQuINUGeF7MqrUqFZsWoM
hs3ZUEXjs2li4qJfrCMexUnVEjW0Eux6PFQ4jDQfwM+EXcP9qIrPlmWfuji+hBmDs69QP2c24qdR
MU9Qrjpid9UYwOiFDgaJlpwfaYxnS65I678TtsMZPlvJrgjI0nuq3R1iohZ5e40bXFMz/w2ERzs7
L9XU+Jo7lduWKjYsDQSdIRUGRFOoEMIwh0HvSEQ9NFBi0E2CPLFHims0JsiVyVrK6URw3CcRcRM5
XMo3OXXjoTKL9fCJ880e7odZoxWBSV+6RWTAaOyY8ZcD3M0/8CCpZ120TCxTH3Cebol0dq+mEu17
oxyEueX/buR/WgcWwKJINe2RuATia6ltGKUu+CQoj7dFJyhr1fftwb9i9UCknU//2gqwe2k9HpTF
KxN1OkNCuBpEy0mFv0ALeiOKgOMqfkuMrOnnU+g9MXdT37Q7sYALbwB5JOw7x3QY6DYTKeADv4a3
ZV//2V8Zkt2MxgapInwlcwIIRERamZzdhY0QJQcGVKMyVurBAT31KaJkqSWRgjZKOObg3D8AmEcx
u4TNvHR/5oEkjTV1EVnPAbg4BXTFaIZBtF03yBil2CFXTPlKlOx4pvRCj1pCdHtC7+BCyEjM326a
mSsj6rBZMUNg++XzSci09MM4Yay1S85Pw3rityQO38o25L5qmugM83jfajVX0G3mkcWKKhVcxACG
ttsB3zHVZ44Y3tCIWyLVVBgp/BGmW1ZVWICDThR7eTZGro3+vvsTjy1G6/QJsGfxhlvjJXt5F1bN
Zeiz6lXjRNPuuY6EJaPLwmaeAugViq0JLBFm47EARTNZLNT/2mCDN/9t82ChhVknsVBkvNm6zEY/
aqeuZ2otFuWSTsxBXt8qVtItKGQ6LSfriRbFh5otW8dEfPkI+hOVjxfhSmN9o6SBSZXX4nOrEuOf
sWCo/4iQNR/SP3YbFH5xo+S8zxw+1vCY4xItO01UhZOM/QoT/a1ynrU/IGI+1MM6APuWyYVmwIRB
s1dz7E5fwsICS5WigI/+rTKJE23/J9/pggfxnipMxAum+CyszP6a903qqUvuXtTRBLdZacd4cfrc
SVw3djw65RlD+Nk+JTBNLUzDHJitptF7wb2NmmHkSqyvVwiD/HnvhSth/mvcWFGm7fBsqtCOu7fI
RrT+GfP9YSyI8t1SfRo0cTr8+EOAAJrasYAeRF+9vIaCpQIcb+Ji6xPIHUf4Jte4BS6QqtzV64Jo
gTkC87bxL6FANCMy2SNDkQ7uTNU5b7p0PUaw3MRXXUgu08Dx5/vHqOkoKOw1aob0c7t+fK6KCl+s
OXStfqd3uT49j01jAQg3VlLXHWmHD5Fx37y4mlkthmO4dGSf32Vp2iKAfygZIdN11Wd+mIlZAwng
erpP3B8uPl0x706GCnMpjuhvB2/OgRJyzVPPwV5orvFY5bPPXDNep8yZT4FhrjO5U9BfKoPN1wt3
H5ymLLI//rsCloUnTRT86hGMHG0br1mSptiD2K/MhGcrAeqSS6IsnEShwFdXOR4Q4YbQRsJapcgN
i35QWECuuTyUvkk/fp7DEjdT+YLqteiZSHPM/wgV29i60qZ+sfGwjl1jWvqdFoctXhr/wo0IRehW
mVD/karBQPH2Apenf3aPVe2Ln/mMRADtvdt/Mnl6Hzlq43t031zI/XH2FgXzNqFOwAC2Q+ha4J1p
HGojcN+TqPWG/dersxyk4QWhB5JFAV5kpHzZzDbKSGzOMnqJ6d1CIAYM1EbkK/YhMQ8OAYlc6JtV
s9KO4suxsch+qUpp4JP4jk+xt3umTf9BZwLHKMVNuXwgc+BBTyJhO4LegP+xeSVQ5CFFcjnSlqMJ
9zHSgj7vlssSuwVpHMyplBp3AiY5KXAsHf+H3B5WbxD7zv3V6wCY4ZXS6scNOEaf3HIip9Xj4Jz7
S8M7y1QhpTpBnuDeCBLWLcf/xvVT5fvWyUfVPsarPJWz/N8rE2K5fL0xPpaNkdjf2++FKSN4leSh
6hQkarmB9YQ4T1uZsmLdTzYWjR9Mt/Z5j0VY0u8i6ep5aYWNsdP3Ut7Qfz3lrHlJkcWbGz5Thw32
UpD/p1beHFGXHUI7Pk3SvH8K3eS8DNEUoiQfmM1p0kNKnUrpSrqyw6lzFry1i5b7vrPFHzB1oWQY
FN/rRguD0qwYC2Ryh4VchHg6U1cXYxqxlfizItSA7GDA7s97+CMo1fG3XY3YQ4SaZpThanvCII4I
WvRK4V6w2LmPZvEMyWpd89FxIYenNTvqyp4T8meUZsYjxV10ZPuPpVGv1XVWw9rTueJYrpvnf4uo
1BPKQtf39Wog+xRZuTGqVLRyNK4/8YtB4ZsDOb7n35Wbphc2HsLNL7Dgbzb0dcdirLkYX19D3Oo8
/XANl52KggCFIMpvP8whwcGv+WDmV5faTxCk15dUKOWrsayoUKtqdwX+WJRIQf+k3LDfdEITnoSz
P/pCBtn2cxWS5wVNfr/YQ4A5IiLvu088KlgyTPL38VzbDtl6lwFo3LgxO7P/utSEUmSoldmTEMPp
jtUY5l6GEZkSQl6irnPRQfehsOJ2uVRuab/1ymtW70GK5RYLo7dk+4qEYmkMeorxrhIPdIM8RoSs
1HiL3NZvE/1PDD9kyklmoXrNW+kCk1gsxg1+UjIhc5Fym4ipDS6Vdah24OLkcLyj1AUyHIQVFiby
ldxNknLWpju0qLL0EzHrLADNu07vaIPxm/CaooMS8ysl8nVsnLNf55IzhT5XClbLDrsp8UJfU1i0
vh1vH6rT30245l4I3ygqaTv4P3pHOQGYsvTMpxS7RSIJBbKkfJNsZ4PhQUTtHZPb1zAc3rcIIKAg
AO4kEs2zQPO+x5SfzB/JCpxPEqnj5HiS32riBnouW+eaU0OwT+aj1SVg1qwWKN6k4myUaO4nh1T5
ieno+xCez0u9m0ZCWIeyPk1iKAvvHW8ylm+GH+7/gQHavtcJ//AsqABMnEeB252F7JWVFtGGZqJ4
wSdBgixthHenU10Mh1JLhcxpihe8ZIURlZM2X59a3j7gvW6PuYBnUm278Xy/L4QFHXmMhSdonObu
SesMs7Wvw1+oG0w07LicfbgPCjgppD1WXw1AOn+y4TnAZXa7fxFl6+VOgDW6CQq6vqxTLC3sm9ok
7ROhs7Llx2mIcBdKNPHpM8zB9eq6zPY0feoHb+Der1WZMJ30ryO2Apc/SN5HiX179rCLJj8eES3i
7mJR++WkRAOHxySOxYlTnbRjSRSRaduvh5IdKqc4/50RcnSihrRP3MpYvDYrN5chR/c9rOFVDCqK
OeaHQvQUO2mbSFsWWmx2WBnEqW0Z7q0iov5Unn2uJNmee/eJdqwb8uuizgjNXRQyvQOrSR3BlDrB
DzWZ31Xv78RjpIfSHi2xtkgiyagLv9P9dWg8ikXI2NIyYY1eBwpQrWYubM9zXFpY3+1tZ4N6JyNT
ufP8uppMql6CgjfMKxsc9K+I3QtihtWYAddcWcMGW9eGkqS8S4luvskiRYrl2Zxs8UnktkO5a6AA
Hm3lTYVBFY/ZJacYDqPO/3Bwu/EcEJbTv8+oqxOHZeFzvQly5bgCkjUTHRdQvC9mHxpbViTbOqrq
rFvxrLbjkLYH+Q2RvQZJ5Y/4ReFlDW8GIOnOJe7yXzTWK4KObUp1wZWrUtAu87WVdljl/aYXiAdD
D5zFMo92LZ4AyAionIvpAZo+w1JlDnMaGy0GzshYWopTuiovvoX1zOaDdhiMn2i1qkpExeQqAjbY
wvknqHqty7rInRhXxecqDDpquqiERFJuZtjcTVCZ9rL13sCnFDd6lBhcNXRP1la7ClZvBmJS8+wV
7KICteWJg5Qv+xWFp43BtV+y2vN/jwaSzPiPvpU/ljxeZu2KpubMcqZaVT3tFJUsOKdV8CVOXJz2
pBI6ld7sREyOuHsgq/ruSQ3HCjyzYJibcFNH9qBAZ+1LYcSS1zcq0HUuYTylR9l9Z6ShPFGgaV7c
0s9y7IgcLq+AdA10nuPPdM6GsqmS6FyVUKdHFuvf/Qu6Sa/2nW/v1IJ/lwTmVusWQL+Gh+fjnEpo
LBl8i7IXShhFTUgiNIZyrSuopm3z464zJ6EH0OO6khjVi8U6Ghaa42ej4Fs12WrdgxEeFZ3qo2IS
x8hrX9TKTLa+a6oOrTto/H5mqK38ZL9cHUVSWDyQMZcdsX2oakyTClEu3alsSUOhIBH0awwhijE1
t9VTPIDT+evT5FMV5aLt6guoJfroRlgT6tHSlPsMV174I01YNttrWn6mhhjgNhmQ9NXci6E7ygt6
wlypvZKgVDjLQPqaq/eG+y/JVGXSxJVwYkwKU/vUUaeglyHpSRZ4LmTfRQWe5eIt0fWBMAqgDDiK
0OpMAoUwPoxHXOL6PBuafpMtdGV4xWyIx+5ikaisK9Z4s9vePx4k8Dv8bB4SuxRWWmCEBMZfFZ2x
hk3tGPDWhF/zh0IZN9DCm4WVJRbUkn8Kav9nw7BwAhmSM/KQjQVgLndGnVqcYOcTIo/0eJ62V7Ec
ceYUmgkUioOdjKcU7S0Kscp1V/BCqPGBJMfqJ4keatl8yJLKFgesbk7gGhKGZ20mBlVa0Kjkqe/T
lnrfBcvva9n5b7dI34fJiaoMWOU4HFwj9y0i2zVKMMTrwLn9dxT6T0OVctPpmfg4q2OiwHH2snZl
5UVZBfqEGBzFQyX2JEOnuE4i27gNvUcsvJYrcFXlNJaya7a8hWvEO2+DVa8BMUmIVMLwiGuuLom/
JCO8u29vhsd71UwuxtbgqKejT1tKqFwfpQb8ujQvFUD+ZcuUFw+sVTL0+EATfbqz7JlxaafV0h7I
9zjwZc3MxS5axj9R2LjVdmi/BaztYLUhES70cb5lwqpCZGzdbDzp9K5aWTQZUwl7O7H+zVS4NFm4
UOXJGMr2It/lhb8s3UaEfJvx0yUf/uvB2iBBgNf6DJyQtVckLF6Nk6StxeJuuu7dSauSUPFj0ryT
tcD2xn7SJPcDgdOZuDa7OuJFUl9Pf4LPXn8tj4WnHNqBJNqAdUr9tK0/Opvzpiv0WCH5QfI8+VUN
rs7qahD5c01iH4S/WqYYau2KUNW5Y0IZ85iaPlv+oVVpYjrAqaNr+fNG2TZ7rCMt3HgFbGC8unwG
QK0vXAQCjmjbk4VsdDhxSeFh9KemNzw2qNdV4gOhduVBCWmafBgfOvDxi/JF6Zg7BObrzCbtfQBj
vlKOHsYsHYDeK44mDPlZ52J6jQX8ESTx5k/wXPVv3c22kH2eSOaw1fffyI8rVurKnW7Py1YZ/iyt
7VoNT21OUcqS6mQ/AGFIKnPP1GVIaDpMgLPylG/vxo3nKIR9j//Rnm88/Fc/UWYFHxDgRaJUKdSL
NBDi0A1fVgY6oQVBSdUNgx1IzP2dVsKpNGLubKTAOEG98vMw225U/XkxaArO2Q5n9RbHH4gsfjvW
xXWVB92FNRwAi0XsjKP0A+16ix9BzmOq/HkAUp3P/lyFAB8z0IzDIiC6uvPy0+m/T6A7D0hLzD2m
ZoPWUYQd+XXFwQeL5TU0yqwbXhgakDflzOSmcP3B3P0fda4k2Y4KEfzALjqh4RGo0bp2fPJONXd1
BXcY7OIMqLCUMjOoPJwIR5Fc//ZJO+MQxZ5deVymqDpSIfBE9PfovkT6NpBKYHMRd4fj5VYRigst
Gu/R7z4lYsNBx9l2BdSy/nmvKz+DJZLud2VON+QDHOnre1ZRm0W434Z5jQU+Z2ZMc7z+QCn6X4PF
ZOdNmFFCxGnmBqFH5aEQdSXh4/nT1pb3H2tX6EX3nbqfs23iV8LUzN3j9b9fpYp5x9cYc8KjKH8h
DvMsM7BNq/TpTEGVc3fLr8fpIuLoXREZTZCbm1LK7OkiK0JpNAbQVQjBpuCSwXJwVnRIGvLwGH5F
eORGXSDyRS4DSvWO2r+SBExBsvcZcMgYWA/mK1X/m3Zhb6gFkEDYcgWC4m//tIKt7QILLgwLbPJ7
G0QMA7RL1CHL0z/ASciHONW7Fu6MhN9qk83pFaKLJ8aRF9D7wx95/tGs8dOHQZfpziahTuufQDAe
cijyRU/SSvm3E/Iz2i4OuMC4E83LaiXBXGg4mB5zxuNRCgBR9vjJHbMgYNJ0YAAKiMmh1o8gOw1X
R0kz/MZPeYMOyQXeI2WDme7tqUWpaQVhrBHwAkJ/yOKBXCt6V9PH9Sc55amf7VQb0BfDPCDSaACI
pdL2jz5gKeCCStk/Xlj9cLi3oKhiWNYMeOYn2tQnrl2aqcoULBcrtZ0nuv4KctK6dYGUyT5jKzto
mhOJkIa8/Js7YCs48GS5mtTwAcJOh1WyHEZargESS0jtLCZ1Yj55HsmF7vSNYlB/MCq+k9pYqIb6
zPKAq5fd2EMjCzUpxlSaofKots/8VetP9JMUu2gq79/2zSL3ptMwRRg54lbpAzAtq2TyWmTJaF/G
IRlkXrguZ4OE1h/fP2r/Pq53EruS9IODlHyaljxC7RvV4wWPQsaQ3br9fGgMynq4Ys6OWyaPx3aJ
0uz4JDnkJELiXIPmkNTLZ+VnBPBZCVvHSTl7LS2qbR9jWEv4Q9yekjzSbyWJWcEQ81HCW+XZdeuA
L2YIguQLpaAIzE2HLhTdzO5Pgd//fom6PFnN78RKCpj0SJouVH8Evkez+xKrKMHfPS1FjvEzIvPr
chCTNGNanL5ruF5WBN5gHkNLKdLW9DXU3CmJ0SIzsSKlW1LQ1J8xc10e4w50Y9Yoz9hHBetx7EeK
3rPniyfOljiZQRLrsKbtwxRzHhcKtwAp+cfb4YZlNhHE+EpNaEAimgbotwJ0kgVRZEZc22qN8Pds
Sl7caBEu8jUmd+9S39qQu+HE3Y94TuXU+GOMmjDpo2WFpcU3NF5MZDSwcVWVsvpD6S0zWtVsUbcR
a3tDB37eBJOfb3v3eAlk4yFNprm+cWvU6TVfrErup/MkIzpEzRiEy4Z5WGSuKURUDv1Aask/44ei
BtN5McZgdmDlzvQdWecfWJNEVAGSGWlXB0K1yMnJjKXuGypoBO4j9N1Q9QuNL5Puwwq14PvEJR+1
Nja/LYVvpzpf4EK+p86ZOp8zj2RpDI/WnI21yZxK5hUkSzOtw+SMTFudVA6nrYz0SxZiacPoMgGm
E5p75c9+BZMSm2Aubc3XtzOuIaSvpH0aNqBPxm+in67waLwGiFvTA4JJVCK1ev9Sqx49cekCdOJX
rfXUHQpXedf2TLQ2b8I3Vk2PPWJ9RGdzMKHsm8c0+FRIFOnlsoKUaMzv8j/TnsaqkhG4ScyJmpWn
kNhsW0cT0oP+x38VcSAJFaU4nhc2/KEvZf4qYKzUGPNzE9YHT9HbN4MjgX7aIlwDX538M78r/gGQ
lxbc7JWMmXghYL1WHPLtAD/vv50VetKIKKGi1rWV7b5xx4tUrXOgoeNcUVaQpkq2hryA4z5QHDW0
AmqTE9EfcSKG3bhoPDg8NlkDzWye3lZD8Hx9aDNIumKpfjRXWjzahE6FcUbTioyA0hAanwW5mLSn
e/PBUYPM3zsQZsYVkFprSIXSf4RVqoeAcESEaBcBG6/GeghEIJ7rb8e2DIG7uyDNJI3gr/Zwzdfp
4HzRqfSSkSxor6PMUyhlst3OAKxNt6Aqe5NINBTKxMqe4r8twS+Ctf+sOPAQeJQhztzyRppejtYd
sjOZKrd9QOewmuht53wYPQfV6Pa1y+Z69SHGVppSMkHLVYWiOCPaSBR+JT1KGsiUbwgU3fQ8qxzw
7362TMtT9g7PNjauTHeu5J/tt0ry9ci+iV/0Ji9QMHEhrJ3wP5buGF3cJFTfrsFhm0IqCgC9wf5V
SgvaG5Co+UgSqxPT5G6nN+Sxamuq0V86MbGLdjB+pgHz21x5hSe1tepfuFlLZinDTnFgOVG631fc
IxMcjrL7QWa/fJwpSw9RmQEIod3zHKcftOXYOfrWlf4xYmwzrcPzBKUy68yH7YVtOhN+E0GKq92k
3m2Y6jSblYgqus8M8IGQZeYv7NNrZCD2Ol9lmfzL022ziRzNGvE6rEfZL+vTeJR5lbCb6hh88Bzj
XCFzaDjjA2TAeJnq2iugdefWnSJYeAi3KYMcCENRxcz2AzBhlLy8AIu7+ngIUE20RBjpnswPT5UL
AhmwJ5SwA/CLnertIDB0eS8L7SjBlMcRZBBquQ0v0EAsqbDM8OInPd56w2P0QM7QKJEGvoNhMqHq
yBfWDQEPB6cSieD3DFQ8zBumip89xdxGVeiiFTzS5XGe/fYxNnCnsckF27QwZSd6Be9JTakUhAwt
egNgZXld94JKR5XT1/uv8F+ceD96cgNN1wc6Blv6DljaYKTo2LU1DVLwHqo48swi0/yg3/zIMM5s
ixCvqDQKxmyFqpdaouoK750Tjl9ZCAcPxENgrahEzCTIrzXqjozD7TKvcl2NGsBLPHTLvrbYAjML
nH08LbyuCNzKEvANmm4MdL7YdwycrvmvD95OnrwL6gr5wAryj6AyQF0pant0e2g8JA31pW4yZbed
nedxtYYWsx5BLxaJMeFTB8b9HLyLLg0FQGpC39kf2PcC4A+TQeGjsPD0a70wzP3TbFucaoiD4DiO
kDJUYPoIJVi2rIeZo3oRRDWiVICfd6z7xKn42nNwem2O8n+a/oSV3q+mtX0PWiRhbW4Gt5EdMlJ6
m2jFmLz4W9bQfIOgjjS+l10QFN12NOnvSh2KycBfPsxXwBo0UTjb80og7hPdYNVM6ggAcQkLj3ek
IsWqfy2b8zT89j/RTv8Ksi13J50SxH/vHxeij9AbVOtcdG4pCSLFyje4zA0w0cXUPtJBpvMyJhxH
0PiyfomoAWH5PZ3Pow7v/QOGEzzc1OCWiZBx0nHiVO5+xi1oal5yHkc3b8G1YgaIl/1K5vGT2+JX
tjNNT2/hxO6ja70EI96+grcX3uHuDJgnY+X/5TjL7uypGAlSse7nlNEcs2mhiN/Pbwog7oAnGxE4
T2vR49DZkLiGaxCt3IUXr6wiN0a9aH4asGI4/fBHXZpr8S96MVGPmIN0sXZwwTDVJABJKo6Elk77
YJF8YsxsIbPh6kd/tScKI3Pumbr4E4o8HeUCfSJuUapYi4FG9/XTmXt9nyM/xXJ7DEnLr8AuHy95
T8j9oXcsOXVgm3Y6lEk4A765mWUm89ab/TRw/sq49v2XBRxRGRmW3jSJIpaDrs2NfP1WTGAR45ET
JKXkI3yfnQcVYRGi7SXtjgoG46CgUmgJ/PuPDtd1FTD0g5FzV80LdamVzKXY503ZshQuT1ybmvj7
Vz3sWeg+UBCzo5Lnod8522KBNLk0IbSicr5vflOowk/UkTUCOGrMkIyN+xmr4/ozFLklyRBHSYWt
4e/5ZJ+m5gNPRBvFgQi8T0CWmDCi3koQJbzf2y/Lt5RJWv8cVs+bIkAJS3sZVD7c3j+iW40BeW2x
ec6ftAbd6sueOOgAB6b/OdAl6yCAJWgzeSz4oQ5stk/q1AG4Zyojc5HzaVmcEO/1XWNLovjJ5HT6
ja1z+KrVtKmp2uo+wih8xx234M7VWxQgjMduKGpt7gZmNhwDFglNDQYODuYoI78kzNEBm8T4fcXJ
xDh3rblDCC/ZQTkKx3x1sBYlH5QNd+M3wjCZBcTf9JtkDRk4aGV7r8IJLREjr6HZ5lkK4grwofHL
fUAewccrNhgBUIjRPrkv9Gu/fC0Zi/toFXg+ffBVKLcYgAepwyyZ+I/GsLxnDdFCm+CTOfcwx/yY
wK50b3EY7gZj1nB7llWgFjw+2qI6GcEs5VkysrjrXFo2x0uObITHHr/ooHa2+kP/jB1xFG0YkAXi
X179kIAmFUnPj+8SoJFLZrEikPguTkp37IL+qoCp+MOQNk0WrTW4HRiRTewbKhTOmvhGub7DiAiU
dVXJcBp/TaC2AfcQeP6i1fcjX9cAJDBVSrHKjJXjhW03tRLlkIFEXLGHjGK+NlhYRRKVEoiImbnI
PBEFn540DpSB1QxGPHrxWc/FUU9QSbtPxRrwuNMzQJwJLYHri9al9x/d3jskZoxuqNjCahSQXprA
RJtZ1kTkAZGTqXD1u6RldB1OricwnsTAcri96CDa361S/PVhsm31MGXUHLa5uW77tZ9tPK1DMLrg
WNl5Z9h82D783EucG29keDUuQYLs0La3SUFiIbeDSXlj3Q2rxDOjcT0kS73CrnsQjxwb0ddhsPu8
35F1BZ92H9xv/GOyFpJJTRNgdQHQy40C0sEWei/sU6GjQoew70Tv/LIm9o4bFulCnHJdRf9exk9J
y4NxmZaRNA52r/f0kSIDwcRneo1SEltJVslzJYmejg/u8j333XE1cgsvGF8YTj1FNmro0Zr2X6Om
YdsmBPPMojymNPa3kvEuKnPJt629AT0QN4SC+WdfFZYpKHxsFeYwZcTqI+1s2IVyPiakqBRNmyjD
MzvtiATWRWtJ4DniIbdmvWGfy9vviO60SiqDVyw2Rq6tEGRakkaeqUZ/1iWv/DjdmXvaXYBv12gZ
7OTWsD6KwB5BdX11wYbb85+Hpyf+Kvl61Bd11jGp6xFGadAJ1WIqE2e2PnMg+e449TpJvQ3oQYJC
cowlC5sfDARUvkJVHh6DLq1tpF9e1aAub9gyF8VZQnxzagDTBXYn9Cx6f7qz3ZQKSo1tSEJlQ/64
bze37UsG4GHLuchjUVoOFLBoHOG/jFSr3/YlbQf349uGuxioLoyTnryDtRczyWX7S0h2ILzCDKXv
TDjWi8eE7f8DupInHH7xbNHOhBjAqkbNjYyRAH3jKLF9yf05YJFrST7W3REjACd6PCoo+ohMiKSf
q9eQXItR2eGtvYkM0hFLkyyKzcDe0G8+hL/FY/z3poPqmlCqbiaQUOWkXnEaG5nX0wuyCSPkZ52e
MaUU8b+HZwqG4ELvJsrxe6SWAwWrTGLXreq0jFBAlYCKQR/ZM9UpOEqb3wmt6O1byaLa+kCfwDUb
5ha705dS1cr/PhenYE4JxFAhlk+JI32/7JvT8BnKP/KeqqGjU9Ph92D6do+oQAXAXna0SzFn96Yw
xco4Mp8X+ZfCmZGr5v/Lm45IA+mUQYH8c+Hr5j/MScpb3JczGBHtL7FcdjnWUcKNM0m4gHEVFOxT
cgF7zqoBtAKRJ1R1VdO2SOdlJkGUxEo0UGsQBNOWs4iJl6dzkaXkA5TDfE/Kgf1/rAxGiQXAt8Eb
vcNTZOiUHbuAHfPTiLxtJDx4X8OsmITSD3AGY4Fko7PML9dwqifn9zfwfb43HDRMiD4MGGFeJdeN
a7wTcHk6k7wmPAiFFJS/CuPfP02P10B3GnQ3aKxv/Koigct2UpYDNQguZpbEHQml+Vqcj9A9sCgz
CH9+qD8a/F35npJznMH7fTWWouEdXb5JD2dI9gLv/UrZwmZV+WIVwzT/zN9Nvrxz8GCu7zxMfNWT
GjRD3c2O4JMavetlcZb7bhVU3QIPr3SCxu7mEfsEjBrS+3ITV54l20HjYckAHTxF9sveQdqKQqkh
OpkzRurh74oWJK+L0/zUdHcfExjxgvzzJCUj6qIQTbmWqV4uGyg+OsEQuZ8uU91rApoUOMSUrPjM
hZ/EZsbx9GIWXcq5/qEhRmKc2rwRAtgSUhD3b5pLgJfbXcVPkWiOUiOWM6TBWSZEJPDwtKasPW09
9HbgKPG7A9jJzi+wuB4afSRVe1S2f4vS9XpZECmsEH5yMFBMyBZhXJQ2Xb5Qvgc9I7uTijL8hXFX
uELnqtYAyiw/kOE151bp6IUCicHMp0lhxeUERxFGFD6M9nydmpOexStAnAPjdQ+0MzmP7xIExgzI
9XPDDf6UsXU3oI1HiHTZKwD6Aom+m8VDzR9PoOuAmz/a2pfrA+ipa/ORz+SUTH4uMrGYk4XdyvXg
ydcKsSwpHTieZqe0fr1rt0qx1kCAesKX8XLPBHhN5SG4E7DT3glovo1aY4TEqzFlN5CGwugo0g6F
/XfqmRZVZwwOxKAr3ViUnzxS8rjvoytq4w7fFUaSpT3fJyffxSd5lMS4Tkx3bM57MwnpG9aJ4JM/
JG93jrVXq8+RGvBzxDX67JJ8A4wzcyzqzuzZzjPQ12kKIphobekDsDloBseAO1AX0jFEbrUEyhS2
3+Tcm2pkUxUnRBGraqLFBNX4aAA/LiI1bsGLp3RwOeQ1zFbXW3qcnhgnNSSjvJZOAdndbkSCvpLR
23MusSeq6lH0+c4+oEUY3QLVuNWnbSeXHWtROOI9KAqhE5SExhYyvixSSnZFqkjJjeKhcwyO1Iik
txpDHIp4uO92UiUHuJbQ5ESQCqk8mHH5wpwVfcQqnibAxwJfCs+gyOSkhLk6Nhn68uiEoeTske5o
Grpsat6CYbl5Rdc83ULQnsHBBAu9eOiTx53tJxG2L/fACkBxz2+5bfkGvH1Sjo+z2ImU9N9OutXv
LzF4HGWK5CxGwu5tiiDpf0a+Iwg7MBR0R+okng6N1emXHeWefe7ZaGBu0L1KDDguMNXSMlWEQd76
zW9qOw2dMvNwWxi/rTB1eGJiZLds1bxOnpZHlsiCi4WkfWctSRYGiQqMLWScgu5LknKsY8RBq+0V
DOHxwpO/XvKBNKyZX7FBD0403LJkUpIdLQlgYg58JdsLppvdyK2YjnaYYmRUYHx4yb+CONYPeimO
XlJDCrJ2oE4CEnn5FGUtmGNJ81L1B3b0x30FGH8Z7cxSEtSfdczyzthd/St4tOR8ucmD4jiJgApA
eARzokMCmXwx0D3rKJYbW5otBEtmoY7P+inVa5QXs6nJ4o2bIp6ACGyy8vgGxSjyym8mCFyRPRsX
8S+97+MpvF3vWHF3ergqBVivxuerX9IVDS3H612teIMHSrpwDvxE/toXTXGqqYKM4F6QWwPrmOku
rBN/7rCkwjzjz7y6h3FMRmBbgkhuRwvWt0C6/yCT1ot0FJbVQtbHptWUfJ+IjEINLfpbzaRQZUck
x/oWz+/pzKD3502sDO1fauL2pLm+YMsOxyBOUPAPTlUWX7mEStg7NhGb0BulCrdnVQpuSNcgAkXe
UxrIbSnfDlexmQCOKJ4cFbDkd9/mi2ViEJnvLoBT3ybfbqnEzJq+wa5YaBg8g521WoWSMkqMZqPN
+a92WjisJL5ZUZqQczGm5mwZdVSzZGUc4KFIZKGur8tqmG7K7/gyTU8khke0CQrwTUkhKWilXMK9
WAmQXA3zt6stjKIv7doMnnn6Y8re0z5Ral+fFKNZCaKN1WBOyzDTcC7SdNM5PgoygbFkoI8FSD9S
vAy85vnSNejmjthxLcyQOqUQ4KhI01gmyBonPrgK1/3RcMUoJsIZhgTDfzhPYsO5O8iVHJ5/Gl1t
ihNG6n+9Vld2WNQKk7FmE8nLcG0UPnJ7FINvV0QcH6KvG2MgpcJAusmrboD0WkWgiAdh0L4FmSjM
cp1HPBXdt5zxVKM5KTFXh9AZkoPagQn0NxxlACX7GIFQdL90sn1rXv7C6GPes4CMYG1R6ZeOdFyr
G7oiuGdNXA8zcEunj5GtnM4qYiuOpa5dg7XwgFnzyCBg+uUiDEpx1c9ggSYPYZEBCQh7GXwsQysd
Q4zW7vjjhG/2GlP0So8NSPF7ck7bVI3OHmNNtK4Ql+xqyppCPCvg5q4zGzqvimMX3P25MXkDmHh/
42p3xkgCqG+OEmEjPa2mhWx9/nR9FLUoz3qnZaasYVi5VZwIs63HetXAsbvtf+f+pLt8PhtHqUQK
z1qSOmQMDRuGReiR2HATU0TVOLSnYNfHn49rrHIw+Cc8ia0NiuWm/eZvttS9OKQz2xQstwzrXCTp
yZXg7GkitCCej1/Mh7MT6NaOe/hNDgp6tx+cF7ufFUZUE5VHjv7EtZxqPQOeU4MxManAzYp0bHP1
ickkVotM6DOw7Al6MAdy/dplrUDpGehMkNShN2rNd/IGEl1Y2JXcgbsh9ZFbUp4to6NtiGX/1z6V
GhfjQEVsAgLi3gPpnk12yXiyc1wgxcbCvGZrUvXXC8Y7xJO5CXbCk6ySkgLMkIkV0WidNZL9Dxpu
xCTVoddyJFTXjjYeNF9I7N7HS8bnh79ToL3CwAkR2slRlyC6nOF5IOa1vaUEH8BjDNUFiqd29JBk
RJ7jmzmOHb1nASolIUrIB93iK5dVlw6vi4Sekke9U/8jHHFJaUHevyWrF4BgDcLvrWtPa6cqkXbb
33t34kkwFa/4By2T0oEp35YiemvxfLseY5WqpLzm7eOjMq8FQqGiiPcajHL6M19hiEqakeW/1C6h
SQLMRLvOLoRPEWm3xAMXlMMW3tk/lYwTueqdPAmaWLFV2msmM+HmMoTtFIOn4CoIvLB/h0Eo81Nt
Bdb6OBwepGutqDYgKEhb/Vm9MVXRfXaXt7f9qZhqOB+0WnlSiinWfFjuAS5DVVaLsVqFEO8wLysi
JdW9Is+Ddeg9J+Lpe/70IhEDjw1JTCkGavKH7L51bbM6m5eWZCHMVkYQuj9NwbY6Yy6eJGkRoXms
r3q3nuIZbBLpYHIeD0DkQwYJkIq23+H8KqNF84SFCvrhUeTJAE2QX4nUcwDqbJxNWj/F1QVd4vMs
8h7+PLG7dhdTpg6KVTBwz4oBK5FEOKBp7ebsnkCIAnF77UwbPF68alkkHDCfkCpY85UQsCbeuM+2
Eg8nlGbk5V789OhU/FuyM67FgL04NHiueEi07v+H8fICa1eoAckGuSLZoYxGf/p+hMR38XPcUL16
AVcI0Lfa3qzUXjD4qXlphMyntiN11j0lyrw6HdzJcfuYvy6/WxNgzlw1Kuu+hCS5veachbebfPeI
ASCXupOqzosiRSYgs0MMnto1TxQVh++47jjblfA7v346oGvZPeEqbFKenOXsGHXxSLf18pBVbT44
ybiEIr/g1KM2EbWGXSTF/jawXqsL5ibSMdGbQumLM5OYQ4+ayEzEZ30ebMqoSP6Vn7RCq3ll4h5l
bE9eZIMY+HY7AO1mqCWV1zXG8VvpF/Q/vdQ3z/gM8LyeaJYc7QoAhahpvz6EQ1KKPHp9dlJDC/y6
l46n7aadKZFMR2jXY/4hHkA0qP5F5p8KweO++ccXeh2Sa9ceDJ7QqIVB1FGf/7jQcw6T/G0e1uUQ
k4xCpQ/MdtXxED97c+J5MewZUlQsTatUoYK08wMSxvouO1hHGpuIJCwtQs9w/06kaUNJ2+E6APY4
IXb/cypK++kaQLx97YN4KMqy7hSg5THnQIx/ugt6b4WjW0RSw/9snfFaFwKU+PYV1UkuuzaFbGSB
WTrXQNkt51hhWWWNaSxvSgy+NQe4gN92RSAhaS81TzhQTuTeOxElReL3eoT+Iv66wZXtWgXf8mCC
e/2wajQvXgRwsnxzm6n6L4XLZurJLGFzOt+m4wqLBegfcGkU031xonnXPz+E93s7SVaBpxoIOktE
VKwP3AoeOshJpErMaVQkFyeBN+hCnD9hm4WTOBM4D4ChORbDhSy+nc/XQRhiOLjux/WhefqZFPJG
599fCAtwR2csFWWi60O1mltY46OgQDYRnrLrBw+LPyWzH0L2MkiPT1tm5MrfQ5BVbfNB4Y5MbhSo
6Zxp2nslGy4f+zWHYYJCzdu5YbqDiX88Q27jf3eHzFIYm8sTcZqMokt0MFw9Mv7r4RAcvirbcS8K
02R/smSBrT9gf8TeOEiVZvFhTJ3Yix/EHVJx+dmdKsCiV5U87fCy4CaYdU+wYsPpiJfw6o3LSD7Q
T2V0uFJErL7L9cAB7SZOUS7cInQZOfmiopYQXYlAlFqdmcOGFgwx0oWYIj+gj5weR3HVgKDD0FTn
cb1yuF673wGZJehv7KFjCsHs/BPcFpWBi5N4jxnG4Wuen77CTllJr/ObYZdzyK1VN+rzYNj0PxVk
0+0P4jLWVsY7hSUgIlT2UDNg09kPY24AG+elSipLJwR+zFpIYj1AP4DzPY+U3b6MZYEgXmsj/MBs
rey03UrNmRsIUugVGh+nJVTh2TUM1zOgOFmNYY0e4vS+mVYrnO1WO3chP7i3O71Xvod/J4VYyWdS
bYlbq2WWcIprLgtbtS9qdV4u4kSQumE7loUfMg1qumf6/CoXZ4mGE2srX0CzBOjD1X7pMX8wbYNU
9eCO8mNAzBF926j58Mmrt7LwaEduim5hKzbAbTrlE5V4ng0z2bRcVgDQnFUj4RdU9g7K5p1sox7V
lW92nEmzqkLb1o8gE6Si8sQBUSbpVybr6bP6/1y19D3F7Fs/LMfEtMwOsxRjxEQkoxfcf6iLCpQK
nxjW5tXIj0GOqy70BehPxAGzcLBRK2oHiGNwxcJ6jEGxWD0P0AOC+UGi4BE22r5VTFCbdyfd2LEY
k4wcomv6VNFunRSQzB6mHsqDDxzBg+fzlDVs9zBxxZ3IqAcY+F2KdxpG6xRQK5XlbpCBBdU0XN49
i74gZmJQVdeJj0c2OJnHwPx8eYchnOVJ9AcN+nj4DPwYPeWZtCEy9CF+1TlMmYlKf93SNtRMl3J3
5mVWZBDlmgNfFYvo9BnvtdLbj+NLx5YlW3LVtamR00qNKWgUWXjmpAk53ZbOWUAUyi+n8zsdMs6p
Ae5gvNkJkd2xCUSkjIZ9OQn1qxk4qY2WdcWHXHS9VqMcCNGp6oJSc4JY/3XJPy8cHhjdi/KYQT/O
ym/jKN2VyxLLK2+D4T3dtGigu+fQZ9rYHbFUSBbTyQb9P+Ms7eTX49r/T7a6NgU1T8/yp54RlNci
/jDXa+v1umRQphW8l80yLKcCiY5QPni0MlpOdRraLmp/XsQcPhOc7qCF0AwLm5hxZSZFNiG2cWY0
4KTt+BcBrbM+H8TdEWsr2yqlQwTHlxsyNq28mYYwmeTwCpTLHKTmWiqdVPu+4qZilgXYGK6Gb/rn
WXVD+hrTCdPS6OzOfzAor5hkC1LfHXfLkeIbxAM94Gf4yW++zhFKtActLegoI5GqhFWuYr2OOYYw
lgLTf1CSZde4POtXixqca4Ehl23sqpwoNYSi+FeWlNRkPQY9z8VUJ5CrZjiAOykhVt+OkrhW1N07
/5jNKDfeM9VReSAuOVlXS+r01ksYEUfK08o7g+QFwfal4PKVI/BY2PFPCWQCIzAPUCpF9hJypBtU
xok8u1dJYY8Rfqxt8oO9DK6p+BVAuUx+fFckfe/0vjYGaWW6+bjYhnKSaVMnWET33w05WzwDSiJ+
qYLN3XugwxyFjjlwVCSS0nwfP90pK1h1xn6RB5XpZiDUv/4uEdp2soYZrYitZcE19UUUN8jZ6DSo
MySVj2gkhTWaz6qCXPRlF08rZ5E861LO8kiZGLpbEbWeqXvJoPINVAgIm71CpZjlcNSdwrG6hHtc
WXduLbteywQ7NTyp3t53rQVQCtpCvuyuGAmrNfC4zNI/7TiMnyFhxJkCs69iUnOHMHDA8sqGs8LK
wuBUoCMDQHzbKDX9fCUUgEDyDBfmWfZJ6/vD5vKRdCwsPyofcw9EP8cf0SqUjQfQTaEAGdiPojID
IKA4AyX6b2bm5te09PXxQqBBZBdCDNnRX6v9mvLCPQpn1YNnh7Y0eqm3elhHH6SoHYL8Ov0FvIXs
7QIks+FgzpgWQAjHw7jH/5e7Vcsr6gJgNpsAn/5NAc3+CQTbwJHJOoWUTbn+32dsEPt8J1eNw/6R
WEeW/qdMUd0PSOT2sz6rDYHllo4b2Fed9t2W9/y3p9s6+PnYIJ+KEnxbg5bnPqbcd7A/rb5HWYdW
TLr9f8th68jaf+bV43Bj88I/FwJCYlfBqVXCXNnN6MHq5hcBvQ947QCBMtzB7p6v1wSkMJGn+6la
GWkfnGcG1pJuKbrH6WXDVOEtCBLmLYqvW/stxjZh1fUKGXMo4m2XBpCGWmG7xpvBLrNjlIT/FU7H
f7EsR1+84XYA/Lol7ndhrE+6P4ZZGTrXqF4QDxf7U4DWTpINfRb2ZoxN69rsRHa5dsic/1qqcpDT
WWl9NqJjRHaq2vdKTVMuxD7E4akgVz5UE1J1awKXyUwB5OT6HHQt6TlHbzQjDgvAPhVySyVudGqg
VdxE2q/jO6pFeLbf2geU8KZmQV1olJV2w6nPe2xHzryAVDyzvwAtux/5e2KKiCLEF9weyLiIa0BX
OrFbTa5i4FpGAb1Zi2/pa2JjP9RaEjrjv8RePdpFKcHq4XOiXTN84+WnuHwYZ7S2047vDm28UXH5
KzNRFuxApIUO9glD9UbEHz1wOb+Y3Nuh6x5aE59TwYMwmPkOeiy8LYmA5EYeWxel1Y3aXsRwMDnY
2KomDpQHMST95bWibZacQY18dfoFH9CoI16A7+1h7qZuhqVuOqpHoBEjPPmrzt2GEcqgsToIo95O
ICjTl0XFVhqPPQv+HmrQnA6GIiNvCZYSTvKmX9cXG/A8+m7kMHUK+lYdsFaDtfmAA6INsouAsrtR
1CL/RvQQYdlv1zEhafP4SqHqE7PZBT7cDPeRD6AeKu8y5C/rd1gD29/owHZMwW1X+vFkfH1mS9ND
kII+oxmF4WQz2TtpNAfRAgFgwzxgVEDqSzakBV5bFcuKmHyWwIXsdnK01kOW0vYhZw0Uq34evEod
8s4Kikcez6DYDDfep+Kom+PMuKrMsc8O57KmwZY6gP3FSekv66+YtTs+gG+nbFjjWuSU4j3bADtJ
VpkNijVAEl9MqVncg0QvqU6zAf89DbATSV1yiP7N+4F/zqHhgE2Vslc/T9KWYDhUbD3A30NMx52Q
0E4UWt+j405dNvZ9JpaDV8kvP8xPV5nsS7+uIe6y9LMUnlg3yj+LfQvseKqy0aPXvHOYPqFLI5rs
qB1e1HPqK/DwspcsxLS0ibQlQDJzhT1L3x0YD5UiTCCtg3joV+BmXFG1eWFLJolx8tMvKJ1UIuU+
1HinJwsoDP1HvK3JDqr2o+xNbPY2Nsh19e2Koy3LN4FvcqmhpANsqdj7smxQWuBmN1wseGDlLezJ
Cbokqhc/+RHyuctzvo/rfpfqthZJX92H/Y8gqiwbMSKtRupcNZAYcHzUYXywSIkvk1D3KJaiMGs1
3n8nf6A0DSOvbjNEiFMRHDT2NFfYQ/z3tPCJPZ9wI+i8dv+fkCsTTVblixNaNJpY6bF7iDJJfb3K
0YHYCWy49pSW9rPkwzMr9PIh0P6NC3tNsijGSehxj9bEjX5qXpjbFZRq6vL4LEply4pHtKQPyhIe
oEO8daMhr5y1irofUDNSdh0zZIrLA9TWrp9S0Uo9uW1WqE3GJjoZGYGmW9enJa2yWzBvLr+6+CTl
VnoJ1zqaE/0XbCxh43nZjv1k4UNmKXrbMOT/ttS/jOlZ55fu6lgE3qxA1UBcW1PbTZAWmqs4ghhj
f35TF3+7XTsqUm0ODWwCUkhZPCxRchUMq8Eb3ET6+NAvGLvfrDyT4VDu1gOhMRWCTba0bbfnd8CT
rVOMYI9p6bi+zvLOS6iB70xtWhvksurGB/0WnhpJB2tP3HNORAzPe+Iy74T1te1a93SCCccvKAyf
VtODuEC22HK5VNL3BOnJawdlyK9AhhgjQzCNQBUy1lrfMo2xLsx34Z3voWtsaDckzTbvPWw/+YhS
2sxKeFtkIAA/poqvcGlI0wjDF6MlB19Crgel+de4QqAC446HaNUkUq/ZIAEEaH4l6EX+UEhgUoyp
KRo+UP+nNA44vtv6io/wpT/n0yTqOk+/bWg00I1PtygEtVTYOXmb+1wWuV8IBHsuZGA62BdNR0LZ
vXHL2DUZNnRg88uWJ+n9jCzt4gp4H34+ujrQFhPuEXeSaYLOAYNp/uoAR6S1yhv8BSvDZlR7rZ+v
ElVK0tVtBMxXliaVCvYerlEpIYwVdFL/27cUl4YOG7dTMc7IytoshvRqvCplKylQC5X+cezB37uS
1ry/p88L48T/2Yv3hckHUt+3kjS6bO65++Xvjebn2g608d3s2Y8LOZ64rYB5uTFcU3jWMIn+41EF
CYp36sSrBEPA9auDolQ6qjyLcJaLk09CpN57QTsUkdLfre+gbjs0MNj4y/zJwj+MlF95VksTAsaM
y8ZRitPCGl4x4qWwB8jZP7UQTzNMmJguVVx4/hDgyDheeOw6OyTrrbpsSY5P2zOewaNPLsNV/WVy
lckO+9gTsfwjKtyXvVhoISj1OPJ2jQHkMBvEH6BlWZpTOxWJgxdjSw6Yuk1idfbdFVVjqmBEIzWQ
VeKLFS+c5f8TGX06HewfnMQQYTVQbjHo5iCjk2VCY4whnYN4Shex5QGN3zLQHQWmFmpgUMHWoqBa
LQ06ioKrZscn6HNeVzY2YUfY4ZFSAjQ4L5EBBCtT231M2CaIBT67lyegdz7RZfN7FzfhYPtpoV6O
RL9SL6SHgiDKfxafrzyUdLJbos2dXQ4/D/ueQuhIieemu7F5XVBo6MWPH+08EwowClve+mD3LR67
tGloZULnIr9PPGegGoZlTCx1DaeJeL6pBFOMuVqYvB3/itrqwEhhWQ5Lks/9hikk7pYCXGeGn7lb
mPcjyV/t4R1YZGxXJSFGn5RIcRo1W79ABntJtIZRATHms/4vZJHCcoJkuZmwuysxNLtZB4tRYPCA
SUT4MwwlExd2CZmEp4EycJAfHU9Yb08p0+xxYYjPuyZPB8pP7hZsQwoGKZLJwvpjHk0ustCVZo5r
lPkCuZJ255TCS60ni0KQ5XXQLxZXm0pohKj9REbF97Jwj+rX/oNitMm2JLMI80TObVbPGCwObBGE
EIBiFh011/6rck8t/jXiCs3amrKTDCOgK6FRp46Pk/hZ7x1rhSyvqywWUsi2L/uq/6DJfrowUHDc
AgEdLytfdPeWK9OLUuQjFn0gPeXOhsy2uXnNac45iTX3dFRsJ8kIDzayUFFVj6pcuDLFIjcCSpON
LUhYZsvUFEL2amgvkqwUlAol8iz1nC4rK8Q+DZ7Dd+IoPB9WUaiNuctiSmrSVUogCdCaFUYHnb9Z
NaNiAJL8Z5HMDjABdMN8w9CSHqYY9Yh2yW111JbSd5IFYimt+jbiK6PfJL9zj1AYFPshaLy2h8TU
wWsnYUxUaqSYYZwNolzS2oIbHIcBxnbVLtS6IQ7Jv9z6t3aulI3UqeUfxNFoMBgr9nA08xUedIP5
zlYq1H+6ApAVJADg6I25QB7bBl20r/pdVjkzANdhmM0L/bHaTMD7dmE3x1N8AV7FpIiDjSJY0EgO
ekqz8PKuCpM25ABLEsNw8NSRADumINDHL67PPfNEEnQBmQEiZQqo+0Vo3ycBgsKyoiT9B6muZ2CQ
BOpwavbOyZm3TCvySomVygEevYBI8U0GfjmqYovPV1bZwFRtOb5VUQUcesLsvLSrRLzufk2uM/A6
V8+MHlgeLyjovGg2JUeXLeFDbVdtcloA6zq6xMxX1QNYfciit/5E1YsS2JIjG5H6Y8Ktn8+fAtCN
Ko7yfMAKWK9aZ2+Wy4OyedVoZupb5Tn0cITZeLKK4VLZ7AXqxPR5b7867g5ozkDaaQ/hNpFr+gx6
3cqViiq8DAcWgybcKTC7VG4p1dcOXhFSviHMxYgDA7NY1W9Zgs61InNeiL4a+poZfWJ+Mmqcitf8
RCSpkaoraJMo2LjOGDhHWz37XeIqW73lF3t3ETVErza+lL84jGm7OZmdaMF5eNh0oOMYtrUp7Dzl
4E5U8CuliwPk+Cw5xNbID0qN1ClOhA41JL3wO6aSNtSLOZQdY8McPOxawOsy9ypnwq/2I4pJOdCL
UuNtXZtGQyAOsxwCRf1buGQOP3JYH1b3SFHtTw03cYR812NeOATPrQsXhdBVd/b4dgpB1jGXaKt8
NMhxnpyQ2vRvRDyKyeLLLAs4njnv4lDgzbFTUqehBiA1YBDt+dhTlRISxG2B0gdj0RbltiCw8tRw
r0w/SADbdt/LzuFkIYB1t7iXduQe/q6YstXPTg0/FvF4oQvNnGL6XUuYVfHC4gGbTKgfHg2QDB6m
2O/MZqOA+352x5XFQpbRiEcUPr14SF1XP+H4WMnscOoJMYJ+lMix5oV7x5sFQ/k5+E8pt7BAYN5j
ZGVwIFtcJQqKMw0oXqYLrR15w6ipRk5rwQPzbXy0cVpeI0YXb9fP28ZdZkiorGSxpv4v6XfOviiV
HTsrwaozg+ZKgW/6PWTbYmqwlKNBhuCnjKxSSVEEYX0Vogr3HhNcdpZGyilD9965SkjqcLxwlwVW
fviRFHZNbm2LneGFkCE/fYnVBxi62SNvkNBrYxkIR68nmVBjQK0wMAFUndWKxe7suThZCSeguJkx
9+qWTkuwDnu2Ec4L4sTmMhbESvN/Jv7DZIEVmXn3tv4TO7i88q7YaWM+ytY7NgMW2gi49GeyWc9D
o34W6I/o+nn5byoWTizOMC82sWXnwcjHvjWMeb5qUe8vGWmYse+MzBZgkX3/Wk53NgRNm5LXjBux
Nb9MJTjITJPrxtJH3jSMHvl++I1M/sKH7mukhUZADF7xvfDjp9aEpLeBwESq6shPr7ZfsG37jFnU
WFidC0OOToTMBgma8VMEl7m0k6rz6+vkdPe9fnTswJH/ZUkI78v0pMmusZjAOIOQNb+BuwIavaxS
WGoiWG9pAKkMtF2Q0cZ0WgHkAJuXw0oD2jLDeySgOHFGCShOjcY6kwmiKNVB9+g7DwVVQ23fVS29
dcwkY7DjVW/SRyts3R1R7J0lVvnWZusIJ4gDiteFTUY9ukGkhq9lkCpEmhTsgftexzkS6zzlkeCn
34JqJwLdQvZWCk7phHkFe/GwANsioCxgr5A8gh1O4TgmxOdbz+dkQmdRclBBcnhYh6N+Vhnc65gJ
iqHx2DqKvJ7SwDThtTOJokRK4wkgK+e0LZYvi5Hsn93nRCLjOSZj8tYKBdZKjUo/ZKbatF8RC6UH
+lJDSJp3Cko+fzSJN43vfc8fgedVyXVODoLR2VLXp154imNEqrpBOm9Fm5Q4hTXNrQ4Cp1JGA2vL
kfCutSn7o2boorYU/TNoU3fZq9KTlc6EQ+7xiYTHPXRl4cXjZtk/ZF4EOCx+PecJGyUvuRcDjzAr
s3XDB0E31w+TmBkxghIKNBgIvzn3MoKiH7gCkZSSCx8FVin8WSgy6kMbYsSWXmhHWXBeS+zFKPcv
Ckl/+SoHAFesPfRqHzkIQJuwX58MSLmGfgAzC6Oi/NGbiX0lP0ztQLDa2ZPwF5k0OlD0nVJ8gGQj
zwJmazP7+AV/V6BdosGx5OKhBUPQkN3IczE/Srex3/WpF8i4ML5RW4ifGwClRZIL5MjyZ+88JXky
qy4+RoH2PIEyOam6wMPXIED86i0AEP/II3k8FQSs0Wb+DDjhoxBty8YWwJgObfrWabsahnowo0ue
Ins4OeoRNjzOfVobeKbme+02DjBYtIsweYMpKHrEUYxJGckze0Sb1ZdX8OVP9wyF2rWCwFANg2Eb
7jxXOTBuANcCkkwcIo5fodD7B3WF8IuXIU8/lCe24ckDdWAUD98uOm7XNzXs1mwdKXgVaXZjPgcC
dHdOSkP/x9dbAjupCLxzDoTaGxupqJDzPHyDeKcUU7LR3mxO/kwO4tH5l7LSrffRRZLafG6OVLgY
+BOwttrftBUKuHnLLPUSqKOJ1d8CAIrk2M7ECu5flwZJDDETVl12aG3gXJcrYfa/CWWLUUQL/2R1
ltVq6xT0AoT+AgbmTqEiTsBjJFu2HZbYb+FCtpaSk6wk9diXqMSOWZyYpvlKZBDEm8zR/0k82itO
XzsHEEwPtIUngUObXbcWyM7Uriypa508NCUl+896uRwqwepWMwvhkfXHvFxyKxUVF2A25Ds+CXHb
VTA24qJOywB/lhZhe3TlSItbfaoXuIfqG53qAK35o+D7zlTwIfYWAGHL9UIJJUBv0RGV1C4tLPLT
cW0HrjnGzPjFwAC1v7lssP1YVPSVYeIEOp+/8AvXnL2ICKzOCP30ooo2V2jbiQhgdBEskFk3W1Pe
fglV0lTc71w8X6y9+vSbI4pthRhcOpD/JIPPJkk36craSAQypXNQXUaT20gOgSU4jnTCBZa22+gZ
lfY1bFsXFjf/uT/PM39z4xum+NOrrkI1r7simjFHReLejHsqvH/lFRKJT1Z6wBa0Lq9qDF0Xr9ia
d3jRe/amxc3PKIllB4rB2UsxL8gIDRBR9miur8IauJBS7JKix0s+nuPuDCtNm4wM4jD0YG8VRB0O
YXDiKIIDjjXGC5TaYsLYwc0L1YguJpJ1woKjPbvWjwAdRyPEdusu4XbPGHxRloGLplTkR13gsvnb
DRPt+tl5fNi83zyaFUpt5HjuiDr2uOM++h9VW5c4wLzfMSKCbUGpschR09woVsVQm3dXKzUz916X
DhxHUZVnyNmMxHLmhR+v2it+9isBmBNmyqxPkfW7ZnQvM/MBO0+FbIWxVt7Sjk01T2wlDWn/KJQe
qEZY2JGySuLuk8HsBmhFPdD4LgQByp8PKd7kDOhecH4YuuN4ZHRNcgU8id1gZqfsWuRoe/syGG2j
vMb8HoKgZCPMTiNXlfN21AQ6rCFb0+i3B2cLOEJaQZXzsuxKRlQx6lsLGJDmWHt0b+ZoCNfLst/e
KosZFrFAVIhKqbtklEPAhwBbl3BTlRPwUGUVtHwgkz1twv8pfwnzveulHTpfrS2elhOryJmyIPPS
rLr0mdGrvufAW51kwn42tmVWCJVc5TcnRDUyrcMyQOyAMTHj0F6tcXKhlSGV3sxD9GTIvWj8P/hI
Ek/E1IOim1EA2KAY505hCUkq7h6Txp7OcAtFtz1m4lGC0MDyzZswyUv6IxXsa+Bw1gA812B3vDqm
7L1uc9aiMdD+7U+6wT8yNo7xzt3GI8QPWygBRM9pFeyew1VhjHqKJT3jf9Y6rfgWj9Op2LOuOkIR
hwjz/VZLuVSBmDI08jvVVD0TOEv74y386auS/1u6RUNGwE9KmKdhC/YUnopSrYVwSPAQ0+xf4AjD
yLRM8jXhrvbVKoIyfqjjY3h/avjJmBvdxEaOYgUUncvANLa3moEqokf+2brLaM+cUzhcgXsSThAf
p2Sd/0ZFl1a2WpHCapG0YdOTeiXuk55uLd+0b4ZMBlVMnjwJoduuxafYE8nCT72rNdU+ItJj/WVs
EeQfC7M7RbpNSBkfbepGfIxNH0LFpyQ9Egw8Udcq0ugFgUIaZOUjKLbnM3fkJJ7nOpbpj99XWm2+
wIIul99kdPPh8Dcursnen/O3ILByeTBp6O8kEn2iocXMmiObbyjkH7BFt+CbJDSPU8B9CQ2SZTpl
JcGDShuAfAcel9PeFZ4n9kef4jzi7nZDdHQPsv04Dzcd8kfCuI8XCXmrOtTZ9V5RI4J8QLuNuy7e
ayTryiRggs3TKPSSlW2CDRV5YCHffXCxO2lwyoGalkceOsigXgIIHRyrwp4qLzmdopyxjmvTaFjh
6MqNEWQ0xcbiFooCpZG8jZVp/FV79LVgamidw4Rm4vUgOdP0ettj5/8W5EUYwlrYclBzRStJyG03
YHVNINSnPtygA9EaOWVTdBZgqGYQG41bDbfuOfyv2fXkMla3iP2cb+kgJohfKQrn6HbMyDwoQ69A
ZF1YC+C8fL0cpkPVtcTs+9YdJjoMnXalwQxFxNayTFP9m0ao/WR+LLLIZrWg5bGeHYSzO3vK7V36
6MqCC5OyMRaaLq4Izc3tDixwdDe99COein1pxmsCe4drbEgrh3jBcNnhmT0oUUm8er6gcbPcbIOp
TUNWttMwd9NNkklrmGkkkylkB4fQjC4IZPHtKalg7Rnu4fH0nUqsc7/izRpSs1U1QBaw32r0flQw
2Q6ps/XIbxRnHRwPVcTTm4+fHb/GYu/NPdKePbducU8Q7uNXreZ+guJULctpwBT+A+SR1GfqCpto
FBWqa+WcpNrBmpZm5BerBKLHe+ZUtBXb+X5WeltQYfODEGFdv18h9oOtkugC95ey5+eh5dvP4nf8
Kb3inmr3ItE2N4FvXvEXYCf2s0gZ+F/NdaPwJxT2du/heYhzUuPyzvckKX/CN8SlDdzcZqRwCHiW
gddAPKb77sbwGttWwI2HrE1HVCIJH2+lMEsWfxj2UJtGrszyKW+YerX25U4ejpIW+PedfsGENziR
SsTaHIKLtXNERKZnSXE95cN03sBBzB31QL4rDYDE2w5k+RhftV60ZEQYpEqzZGuuHy+Y1UkWAf85
BNf46axOorZ0vXqJdvJfQajTKyV8Hyxh7qoED4YyWLlONKfW0SU//KXQ6GVHX5gwk5XiOmA4AOf1
i78/6Mh2lp8Zfupf6LdiWjQTAP+kU0UFKmuZbFL+ImVsDxw4c34zhHDiBHkx6X412JvoK/cxMtgU
/U5t4hFwaDE98T+Duc1QejzwEuaHMud4GF4eYnybUN4kpJEzAA4RJFsxFv2T/CfPaHYAeppK+MmF
eKziRTIK/xKA6o6HlNToOK6ojkBVs30fl12rM9Rpux8KFK9FqZhIgnPzoGV5jqjzPxsVpuDfwxig
YnI6AGZ/2A5Kgp7EXo1uLPurbv9dP/bVoMeflKDatFhLtf4wdDC1KglW94CfIoW1T3noVAYFPhpB
nqggVCH8ykHxBIQw2N4ot0uZUMQYszrUV8Vscx/7ngJaTIXkUUAyVJPNFbdyKFtUaA3CXLc3uCWU
Flbf+DIOOncLy4UG7SufshA9gQF1RThq+r+sjr+JyrkykxG7bBXUVEMxgOTbGsiSwPpzuuhhcU5a
55/ZyoG9nKTen2qkQJOhyigFIpfXrtU0wQJi12T/La5yK2hiMGFhZSUi7IcymVzXsHiHGroTXcNG
Pz+WYLvs5I5Ll5NmIuJdGh3OVF1VMg5I00Ou3Y0eBtZAGSGibg0xQ4oTkOEKivsmy2nIw2uJJyxw
49qkIVvvKfbJs9v7kXZmN2yGgTxQ8V9DE+RBrgxDS/Cm9Q/l8FBNMkJE+zz4hRMJNIl7mrtDzs0n
g8IWv/K0124EYt3dGQ3ibQMxt7v6WqEYBW933q8grvAJkVWZZloZcIJWLt9hkaCb54gyx0uoS3W7
5bEwgxu5CLn68jiPw3jFzwFLwZXQyGCxqm0mYeevZ8tGdgiM2sHE8PD9x1gn3tE1RQdeb5fuVX3I
PCt4+kY7W4qhHG/+eqNf72j96r3s+m+Rr2Kn1N2sq22p1e8V9yHqn3szxEutm+GIflbS5LczSKn4
ww7RG0H5VlALqR2YF9LuQrJGrVqYgkvROwQKtsWlubFQaCByrYTIel8kwFcgD5zRqtkDqVGaiS3e
lNhaEhsoGY9Iqsjd3WcU5eJDxDKXROoKAhNnv46VmZfsWJR8L//zPrl+tiH0DhwZzvhXDvbPyZdJ
Bioyl1tvRKsh0DHKadmG7/gDIq3Z4uXc4+Vp8bgGoczPaN2/vqyW8IUYCZHQYGXcXeNMTf2H3tLJ
wicZkW9BzKyTmbdUeuO4Ecz9ZF4BbQ6DO6/Sehm0OAhPytpu0Dy4KWs1RB84wFSJ/wphf19XgCqW
MmoO9zXW4iGGnbnBH3SUMTgLWX6ikogrmKw7XYO9T4122jDH5Pp4dtR13ARXNOhz6eSujZ2bJ6Ri
RAbXno0dOS1gavL3Kkqv5VH04WdWY5lmQJTDd2Spm3UWRrq6sJJT9QWBq9dhXQAi1/RMsAkxEm95
ArOgo5we5vxVR06psZTX2kooJDF/CookbiW402p+rPvQPgP2H80zPA7B+leoWWaNWnXM3KEPp6cY
IlHl2DnbNHDQ5Wpk2Qdau0n/gJgyZ37UnWsHBnEts4evVTMIIbmCf23gd25ECJ3Nl4NODrmvvcEj
Hlp+NJaTWYaUEL6LPBmnnIVB9ry/gaHUGyRCVKoHzM3BT10ugKl0pMLsP11fF5CeDHyljWm+zfZj
bwILc62Ree81Z/KSAQHlU1Qoc33iw3uo3S0DoLMqRVz7PUNbWjIBRFKNUMjmEnZszPuZm524uE5o
dwicxtWT5lOTmTbs3zYcC7j/tJ027r3viN3juT5atAj9x6FRBFdqHZrlqOzTVGnKXt0/oYnPoYI+
876Duf6EAlJGrfQzRQdcDFDq4L19aBEcuLYRnqUPfasVN3akZBk5wlOWXJ/qH4BaBREIaUt6Wj7R
T5HW6rXxtCb1ti3ku/M/1bpIiKt2otWz2WL3+nYwp6DNMtjgPK3+uvKxqd7OlrxE7Y7OX2CNwzL1
NIuxlZSpav0LMV6+7W7/dSPwXBZJloWgpbugkqA35/EOjxHICGJbbpUDckVL2+jVlJa9PLo19cXd
8Xb86OoYHBm/8mq0Ah5dHzG+qtAnOZ7KOE8XHeic3JDgZ9qZ4tdr1tQfJNnWY+f2RZhLdLye6oRz
v/OaovhdIAx5y5qvEf3Y9DhzMdRJX66k/M8TwvLbHvlspoo0x3wcr9qfBLHS3I5uj2PNK8hytD3U
Rc1opmj1tHntPMrk+O5c8WNgkefySArS8a/XRjul+FXE0fPGNivzQWF8UjFjLLxd8uvO7dnCslck
B9spVNUkP3xNo6BSYaTb809Ws2Hud2A97F0EfY/k0NCzVfgFg11lOVCH19icVFCb6NB82s7sMFgb
c8kePVzRxwmarGBJBsUFDNuDygW2B/JPq8CsGTjKtXYei0kzWtiJG5VrzOy5RiNqc6vqO5osyb7r
cxld12UGDjVvvB/oVF7m3PEg2DFWOXlNOyjcvMPVL0YEHp1lFfZiSGfThTL8qHERmsUrucTVnkW1
CjmSoL4vyV8/FBITUA0q6s6bIvR0/goPLGPKpggxNF/uaA3dTkjLt7uhFxPXeOJbCGgN8HWrkrBh
Hjqj6QYIrzLb8GHx7OflsA5eci5FiKbp3s3mKgYTQLhgkXoBApjAO1Y3vGMFkKSNt+gHDjATU55e
wUL4HgKDk0Ckt/ze697iZR05qNB9Mx1y2cgsTEvQp/GWpyO4x7FpacMFZM1sCh7JCFyAeSg8JuQV
+hoR+c5VYzPrrutc7ncMTLMNynRYrPtVGAGOkJgckt2wPgx+YBsZq9OuuQwiS0zONDoiVrZtRjKQ
M4A/0uTLMEJDcJdMFFqSJTFxJ5sk35j6KcN/VgWwkDLWOgraAH3dDOzg3Kwq1Rs+k9UKP8AgyPdo
amT2eA1v+0r3GgQuBMxpyLIoPu1bJ/ktHJU1RlHRsMHXNfiBb+qgSJpzg9YYW5dA26d/xDwJHdyC
/8gZwdEf1gwAsANbutNN2Rr+s5cz+52nYaHQ9scR/CHlNT9TUVhynxVjrWHHtWrf6Ed28UhaXHIS
xyGR633JqVmo4E/inl3rw904awW6h3KLxw3KtGA7ZuZH5T3cbQ+/h8F8LE0d0484v9UbYKoO65db
umyAtFf/mUMIy5ZsqHwfRCzySaoiIIaCGsZ7tX+glbgKRwCgcbwYD1jbRbGuVPrlEv/M1Nlz8SwX
NV/I5Hux4kFDlH2xId5NJEYYTdJtqLGMgN9x1YYFmXLzfx9JNe9fjhMLV5JLtk7flcoaMQU8//Tr
cllmrgRgucxaSTqGMMNfFz0H4HeGlBxSrbspIUZBHYrARfI2kv3pESKjGnyey3gSm8sxAIDPblYH
1FXk3pH+O2+9IFj7lFgipEJiCyp4h0wSXvPhB2rcW0D8lzFtXgdzna7HilHETXsk+gTMwBwGo0aa
QJcj1Gg+0NHDwfZBYSIf+CBvKyoaYgNsqxdjKKqk2/MvvFKzQkH1ql/fGDb+wm44ABTj7eWKMczj
PnRrbM4bdigLqTPLKYATflVXZKB5kD/raTvBCAY11tDG4l83oJtDUk9rnj8QAvTNe4NBBb1yuB10
XsI1lzCVSlJLc9e/iBGQIsfoIhKk8EpblUD6g1euY6uQo89fuH0jzo0+POifuOrnnWPUZePx5n/s
0n0V/1z5P7PnW670TlJ9mGqaVy3WZOLG5iNU9xGHgYszHw2/52V+qugWVnmqUJZUl9yHWInvIax9
d1118/i9bnP1OmCXdXITyW6YjORJMs/9galzxGe5oMBcY/ghLffcYm3AodUXoHjQPn0TYijIj7/C
OthZOuLZUIMODr+GNVMWwIpwepDg2WqIGl1Q0kktKHZec4YISusKJlu38TwfwSUGImhJvarATWms
83l2UwvGALQUxbT7XLe9u94FJwN0M0uMaaq5ZTXq5mH0TifcWU1cVuvTD2nXmly/vm55SAqxsQPJ
jy4Z7yBxSHUXllcTou8imJ9DTQ4mVbGwJ46cGvp6nKqP+YcQA3a3MLoAilf2PePj9N7R63hxfBqa
8wgkTraiowMkzt+9lPzgtIgv6glTSi5ixe9LbC/ttvfCgeFrH0RyFsxdt8eQNxs2pKgzPoIAg/ZW
WRncoK8x9jIg4mVKK22InQV01lGBjKfsb0m7M29yDuGLDe+uc9h1WOCn7SsGo410Zepto6mnoh7K
SLTQrRGAuW0DBLzARYtImc5GNpsQFLFM92z+W0exo9TRhWwvp3T5K2KPJcQmyuX5EWgdsoo6zP1L
0sFzCAIUDwBpEzg2knENzb1j4GOfXrAYsWhrhuEFcOlEpZma2KW0wT+ZYuCvTvVwZqw2V6xIdnNQ
4XBqQ/b1dRYMrHWR3Lm9sIge9ZyhVF05Rzd/IES2ZiuUGE9uhEJ8N9hKdERChsNFVeROThJhLlNk
ddtfQWpzFxL0tsOtovGTpYgtXnUdRkM9nwx3knyzBMArxy5khaucB5ikNOqK9cy6pOoYVGc5nkre
dQEOvv13h45iKlQmZbwu0XuM0GfeZWv+F7cZVjRii901hJ+bb3vx3tzG+sJPBqgMLpxG8j8QPKAe
goenSFxw00wkjLxNfB7IcAdv2A9XeI0HuegVq+9f3wZyi/0tLSAIpsXI5AMlPCVS+DUkObTVCwVR
rokAMHoi2AA62iiqroI5smi+ndYEaQiAipOSp6lkUbEz7YdAVTfyl4bqtU5Uzh5kfAn1Pof8/MRA
UnNOayDtC4JZpMzO7+Z3ITj+bR9EvcRGTQrtHCfjgWXbIJ0YFCzbcvYLJLwVWu4oI49tA18YDzy2
VagO+ML1aIwpN5/o23kuotZY+rbaCLJEqz7H6qDuk3VUuOdm7nYIdOgDtZ59Sy7iWZum6BDjXAI0
Ioe5tKH136Q2sEyUquP/ThVf7OqWzDpzaX+GCf6TZmCvHrpMyYteRfYGrxlGW0TOzZoqhyBpxvfV
Eb83OWmYQva0x+10mSy06CrjcPvNy6r3C+M0SKtNA8IFeARy3Q1ZCYQq/etXZJ+NSx7XcJIGXdSX
l5a7K6ldoN/yCHuSHtGhezodyuz0EhXo2zBuO5aMuMI+FQTnwaLK/DyHbST73fjAL9fjYBKcia06
wPQ2GJnUnlpEjJwMMQd9lnUG23bMm22qedP1cLz1DbOHSksa7wDtyHc0CwuFSxunA+GzgvKxC+h+
FQeHMTB8KtRtiCd03DSJYNLPBPY6qbwpCEI3Jqqj9vrVXyCCA/RR2juGbPfQopRmud88nfhkfUYV
YgLprPg8hUmyaZxrfoxAnqYody5AZD0bjLgJpn3e8XL0FB6OZn3Ygiib0DinZNmHrfH9NecHf8ZE
khjuNTaIsaWXrNjADN61dPSwi3TZzUr1Nal8/7vIU4lwcgctoerz1cvPJwe6r4wx8gjZAwrf743w
gl+R14OnLtjdP9ctqcarvL9ATLoG0OX7vJg/HOy1P3UtretuY+jaGFj646Cp2sOv3vgxDXXD3NIp
W5WkqctzbRfLlFBG9d6yHcha/KdwwmiLs/y9v9yf0GjnDZCKPhwh1gxpixtORhy6cDWpAXTOvxvB
qNikPNpgSP1qG3sKLrfHAbEpsTjOJiPRMFKVW586UkMvYR/rHqBTLr6yoA7XBI6iKYOuQgdicGtY
2fb+r7bBoUm1UUSK9DEueHZBDMx+1cbqfRHY8/R9TiOgsvHfYIzqWsVqJ9gDSMNt/jP+czx6xxiX
fASOt+pxJ8Jh3KOvcsncZbpTBAkyek7cpC0gdMSTmYtIZk41AYJelVtvUWN1SLqSQTYxvS457ORU
KK4PbAUxayiPuRijjAvkI2u1AYiAj7jupcMwa4kLbLu5CdDKClIuKN8Xi2yvSjuYgXwB5WjqsRXd
hhPqIkROBacwy/PTi5OLninH/IjM5t/dmG5fH9M4T1hSeblI7o58NoQuSFfylkZH1N8fjbh8Ek7q
wQX16uPHrPIkqpd2p/AqQ9SSMZNbsSGeaWUmcABrWWs+MqbhywTXi/+MPrEh/NNIXQ7pHIvLJXDl
NSj/JoRj/ug3KsPvY+6VIaf/SmfkSYFiK8SwIQ3LCQ7zeoGhZFWjgcr4OXzSVnNcVS75JItWIgWf
lTQbh73K39DfAbHDcXwG7H953wZFiQMrI2cjo5AxT381Uqup5MUQMaJv1Fwp4rfCAsHHLRtZKMpQ
4XpOtY3r2ti2RcEetlMzBMhQ470iRI9FohACxedqbo0T0IaRQcUVVlmmRT1Y409gVlWOQGffvmd2
Gyt8cRTsMIz7qc6P4RX4XFU23/XNtJ/R8AW/GOC0j7Na4tWJrk/tmTaVnfAnH5JSYB+zqIMZ0Its
OOuzXYl2jeCUyEsoiSEtzwX+JnlAMLyo0PpRMfP08R8M6HEGO1vGG4veqSK+7z5hBsDnun1Ku696
Lpgm0pXYKccvkgrl/YODV5wlGGHzBvd0aBobCdyb5qCFISI/jfZk9GT+Kg+JhRKd1S5rOcBGhkiv
qCfJeva5CEHvBS+QFEX443mHC/22GT+aVskSGhMdFyrtlARXxQ4al2wPxeBcvc1iGdPpXfi7/37k
GLGedv+S1CUFlYyppZfMIYaXbmFpE7EK5ZzFx/Voz1zgbK7UCT0vt+EhzDGBAvHtsUMfsON7wyRG
fPbpGlSXhlrB860I2j35KV0aH2Azk09Pdo+EI14uiJW6PgruFpJeZwIA3hG6aWOvOag785cbI8Bb
BO7zZ5TQxXxl5nIpCz9mCQq1BZQl1EaHrK3GZmg/1BC0mo267lhuqxO5Q0NNnEu+8DYJwVY151Nb
lKvQhy42bRclvmFse+W1s6y0v4V22w+L1f7SPAZwvXBH7w6OvsYmh7J+YVEviD0MllDmYYDX7dMu
3Zhqpf5leXaHfefJcwnM+GogxQ6kW2M7ZgcdXWAEJLrsyX98ucyVLiPJhwkdyOdfrc4HmaBTMnGv
N19g4rx/GQxMRkHmAdz5lzwVGGdgC52TpXaonjulD2ACPy7375FZoOuXyVjBzl7Bwe8QjMUYtzyc
4VLURHb11SdLXzCLDk4Ns6wcqEXZPSO6UqKNnkyjWzpk5iAjfBpbTy1cmaoln+7PCrIE0jvqKvVS
05AJn+oX28e2tNEhHQooVXKENmmAc71UJfmNLWqRtqOOxpARCtNsUt/YZsQyOcR9DEpEA/GmUk7I
cA3zjIhHXGmxPaIHFUoZrNBoel+ssd1xs/sMJyy5YIZZavuGETaslWGrQbFNWKLCxSmDE8i8bfrC
HPrSVKsDJR+x2BGrLZQik++3E1Xr/93G9r7IGT7Mo0CAE8RqTGCYlc73GitQbpBZNJ/xd0EbWpNE
UOdXfzHgjLL3E5CyYPr9xTLxzrQKvjTZzFqo4AwhYzmEOBfkevkOO5+UeSPMYhXKnI+ul31BqWcV
pxbP/z+T4Paw+xXgf3CNgokZ4U0ayTlftyav5+lew/CDYkqM6dbRLFg4OdywdrDBUC1J3oUrhvog
F84FcbyZB6QHx7a27qBe8BCpje0AGiFI0Zw1bY2yPGygkgDFgeaTo0QlNYampY77MMwHEawaGaYs
gkPwxfi/7Yjd4rXUVKLAaSZ0qFlG/rOX7aM04dTgnF6Jh0gUm6QomFF6GplJNNlbYFb3QSQ2u3sa
QfFUK8uC6nwgy3PIs1+9Fo3nWy8o4lXO4wS0oDBeYdGYNatGG4/vPLQwb37yUJ0BES/NH3/Qw4jH
YhSOSpQnnUa8HGjyZPYHlHsaH5dtxMN97350dyqtRHR8M57vZ89cIXzNfeJaRxfyQ66eCgFosB7x
IG9ng9peShvXjNO09HU1+OsygW3sx96XTS2SICDmqivo3/dL1E27mWL0ex8jJnzdKZFsnsCyJus6
9WQNr5a10BaEkGoP5MYe1WgOQFseykIM70rTQT0D7wVbzynaLu2jB/2WRnCkmR/9WfkyBUZLlGWF
M+YaIaieMfN38bMprRJB7kUgch/T5WYUrUrznt1if4st2gXiCRFGcMg8rEA5SOfwSePoJlnBIcQt
SkUoPyxy0mTPLgjeR6Afr23SeRE8KaDtiPr1c0cP4VQiedrBW3xJvkgLoHZDPLShJe/ej7mcZGWc
Lk5W22Vbreeo4dIs+hO6savafHzt9heEMKFh+LIQzSSDPZlWdmVNAzi3inPlQjadkhCTin9gAvoJ
0OTb5m0iaR1Xz4pGFl23t0vcgaOjdEF0TiPNy3rRCb939C7AqTl2EX6G9HIkc7Zumr02Ac1F62Xo
PWVCOn2+dL2if9L5coFEK8ppC8Eu+mYI5ldTxCPivBskIjlGjjOfUfTOZQTwdS123AZy1tvvF/HD
/QaPWP6KlM0yPvaRZc7yNc6pimij45+cqDF0rC71upKNr/c+tmU27eQkyDifcZghDmYv9QeF4+tR
M0wnrs/aGty2COxM8Yj6BBqYVGf25AvPwSdxxulifReKk7F8+PWFDDE1SNTXnAyr20fpUrMDagK1
rZ6mnA0jxMiv1JMu/bWKnMDrgF51Vx6erLqEbyOlNd1YzUxrFbz4YanI18OP8glq9jOhYXrO8DUq
hVHlRhe5FUKwCxuPTQ3Y2UiIV2RKOZn8pYBZq+Ly2BCT7ptzcfsd71wFxPCQQ3c4jgCIKMwocFqb
G/viIqNw9KunKh2+sNAyb7hQdldnBNPJRbnnO2kDOPbEyxN4kp4pTp8A9/8odOvZclycefFW3BBJ
2acLo+ScZ2SU7q4/Cvz4ZXSxskGTOZosqyZprgc3u7J53KWb6AlWV8lTH3j8h9pjdIosd9w/Av4p
xdCJ4q7Bta5Wr6qqUY5x0SnXkHlpMqOE0Ea6nun9qkCLyDLuH3Y61gkIxZ7zhYSvK+ViZWWRrs2D
lDMR1ViQ5ri0npdKu/pMPvXlqEi5Bj/0ahWKRwAPP+F92zSK6hIsi7oDnmbrTpweRXMyPQaUFImd
9lw/V3Tj+ofBjcOO0iujfA9G4At1nCgzGe4b5Cr25ENWJ+lr7HAsNvH5DVN+P/KBFg1OXjk0EPjk
SYRyRI+HsCof0gblr+6uixOX1p3V8PAyfXGxXYlS41sEi4UHs75Hnd9YLv7lYxhw/+rKRgGoMDno
DYlIszSzL1//zlX3h280HEPScVMWkyVp2qx5ZC0rE8Y/XDY+mspKogrF9Zt8Zfxga4SZyZDIJVFi
H6i3WwX0PNj0LLZNaMFRjNf0Xd0vZnAQiJA1Zzx1Pz3x3/U18B0MP9vfL3J06QVIyirRclXFia7e
MXcCmvA1zgXrqC2fOicGAn5FW3hZ3OzIrNrWqVcwDIvVulVEfV/suQY8psr9S/Wuu9DEu2RsaBes
Z+kmQvAnmYfvlEGwwxFuV203XLlNe0TDCVkl85IPdjXLy9yaroEd9ipkAsU2TjA5HvuboCElvsQt
0lDl1aZwxWxzPS8eCZjnRIVXZjfQ+UWQjEiRnuPP7hyrQbkEBt+G17NfNDRaXcfVPoOokwIjbxel
Cjp5ooR+1P0ulMSMcdF+n6TcadPDEvbc5hq5M5ZDIQRlFT9HRlnzBTXmhLlrCKAC4+PnOJeUIOo5
FEjwWsXx6RBkpyammVMenv0QK2IxnnIX2SY+SC7LOm8OvEic0ReY8UeEP8luegUJhbu7rgrFe9B6
rYxB5fhkRYz5GHkx6OBVfCA4Em0mD5Kv4GBqql4py96XQuTXXHtgkDTbS5XqAIkJrzYDSMPW6Vfq
aw6O2Rri/L5+g5pvbQ1NdqF4MmRdoJwOasNYk2v+SjpSnMla1Tr5hY+1bTwaR+B2DLiIQpLeFk0I
4kcf+alpNaL5JL3j4x35aw42Obln1zf0TN4YexcVQJRTP+SWUiYNLwX82CKeXjynZB4A3BVas66V
9AZZxNzD4g8xW5QoZ+tGZJ4bcELzB6OeFmwLkLdeh5xvdCi4133KOxNAYiYsTtYjXTvBYUT1OFdV
lJkjqdr4bWwSGQ4l7NfaLI/HIUG9dfcLxPYXeF8E3IvMt93cZ5snAs559yCTqPklcPWKhm8AMIZn
GVURn0oBM8qc58xx5V1zENiXTxEJAdrsGUoUPGSS9ewidG4wO7eXIyYK3MKxcqWqKLZqhC6Qd1Gf
CttyvoZ79iTk1FQhmm/CIT63eG8S01IWKaqMELXSyU6oU4QrOukvieQvBmEzWOKClr5xXTMM6tfw
skspxs3+qkyS3Rt3Me8FTiCzFoaz/Efu8/crSlMPSbs84DKJvm5Bg2bGKTngUwZSUnpUkn45eKWE
c7Dcc195ZUHUxCMaHAwquBH7sTCBmHp6oOmrvNKTcPuMahH9acX/cibsXYurivPgPC47kXjXjGiC
KTs2b22ltDDQQFI+hbvuCmIAG9l3ofwCoWiZPEywcMOhiWg96gNKX7Z1MSkNkYOcqDg7FR3Hwch7
M/RLWWxpZMnN2n/CS/Ro/ln+1jHCphA0yk+SdJHtNPhjTU4gw9zfUpPRbySTA8CN597mMHmnuouF
lhRgpNj3dFGimTmASCkhctHAbX5FqNVoFP82aclEIxZqBKECKCVmuDX5BvxOwxiA0eZlPJPgZmEo
TQPlUV0Q3C28giUBZ4ccbdq/1v14CqIp0stYpHSeNa/tdzPgZUxYljnQEXxS6b49sXmTnW2ZgHVJ
saNp7/5JyTLoaTKsUvXyY1lgm+kwZYmGv165SvapZc/tAoBQCgqvWdr5bAoPZ3k1wVzBfE4t8D4P
DH/cMT5O14/XKV+9h3P7dimnAgHhRVn5QM3p0vs+gbVAjCnyQCCmwTSj/CwDqDM5naySNxYPck86
zux6Sfdgr2Z8dHm73r9ZHzcliFIeE1Ry6oW/yFCX13z0y39JqtEdu/b0gJlberxGe1L5A1AICfET
Wg1/5oE98unN+ykRV669MGgcKffZK+eQN3ReYSt+yGqKcfWZnMKr8iJ8bc/sqMvpSp2vrUT174sg
VXyDP+b5EwkBKWQfDRaaQ2B585VwvzBBgnlZO810kS/uhDqzsjdOhSEeZh6wWzTk/kxJg2mDQ+Wi
kEvVL196JLGTK6jGRHdRod7bilo8ZKWamN1QjhFYP9249hda6/BcINusebmZ4reByCuLcejTzNaO
e/bMzzSD6+3Wo95FcNTVfE3keRxJBl8uyll+gYtxuqDvEDsLAdx8pplKpPbNrHN0dviT2Ip8CpJm
HslLZfqmgXsyVdL9pepC3gxqiXZO4snwDKKqS7B8rztftCzXAL2lt08NlHu5G3/r6jEWhC86+rcM
2+OYe+t3clKSoYXpYUyL0gaT85OLvQ665l+x/ToqzeLW45eyD5QyV8YMTwVTN5FdRIDRi7g7+Q5Q
BdyZWGigbh2WCEhxTFmbE+UYFpXWcq9WzozdtIRAfqlpps3W5bbnoZKEgoA7yYrxGlpD+2kxveYu
iOQf0HS7DhLaUmR74KExee0j0o0arzrmhtFdcYyb1HBwnqhObSb+wz9dQN1HeJZl+dBVNwvfcDvy
/m/LWg+LKmvXZMzytcCaqQVhPMnqf7GEkzsm28bclq4momvy/9ZCQnRFJbFq+gSM9TXyZEQxcpYI
jzdzQSF/gA3CzwCnnS/kv0hA5O91JLVeKn4dHxVDdIN1zgneSOiW11+EhVe+XQm55h0A6kJbLunR
yJJqtczTq72NHwdt1I6Cp9VRBRWB8r1wYJTuvC0LR/xx4lkwOudQujAYyqsAZNy4Mkh1bh8Fe5UH
Pq2vaYMyMSQVUb1P+IypyAaWL4WKRsGbTBMFsTxqvBkime4gLYo/Y8lySgTbfI3HUNOKhPQwPo78
dL3UeaJWlvryiLnmMnnOGL4OVwaukbPfNFpWXP/blMRICLkYbHPn3uMt+vXWoKt8oiq+XWUsWVsp
0sjjpLvZJ/6Gz38cd01Cev/hApInJlDPdmtrFvvu4kpnw6uggyHmIfGUvI0hdMsLuqgiWBA/lTVE
s+JVVGC0hMO+5pfZd/maaPRo61YKra0/gpAuokkTGu2XLhfDjuwUY0l3qLmRLT0DmeTTi17kO/VM
jJWhZZ9DXcZIYGSduibF+8yzTT9daD2uwRGgIQEZFU5pV01xd4adkrH4YIF5WnscSLSgR/mijfag
XR2RZCYZ3/s6hR5i9MUvUBzgThC/TJWY3YU12XfZDp6FntnhcAe+VtygQhJG/yBvN4XlykYVQW2x
kxHdRC6UNxnYa5H97UZ8O0IVzrdCYYGYprjxuEyDLotQB7UfRE91dPics0s3E69s4sppuj5UjEJR
8CskXPnl22WpIU3fFkN4JtPdwo0q7K9vgPodV1ctYBa1zSzp0Tz2iPXHBEZjr8J7APZhZtbBJW+I
gzzNxU644O0axTUlDuJCz5wD1V+g2x48NspgEt4ho4A/DNUiaf2L6JEnh1Kpti+HptPgXHpl0K82
LgE2BzJYs4rz43cD1ym8RxKYF876OeM2Xx0rccr47G9yUuuLPqOh8GLCDwU3wsyazcji32TzDSO6
JShAwwjfrXg0jaPCmCAy4VLUIvKOgvCbgx7inNdwi0VIUc6bu7A56ISKfZCMbq+KLSVdTMg9nSpR
H4Oy1vDwl5MV++3txj4Na/UihnNc97t0zUnQeZXMsbVl3Gkpl/7OMVEstnWLY9EDosM3eCs8RMb4
Uhq7/OaHd8A8OLYnrNlnBVvwlWwTLjiuQVGcFQKs981ugLH/SeMwaFjNGbf4chvQ9GxdayICsSjr
XqLyVGPl1SaBh2CK4eNIw9J34XkHpPsn/L5rAjSupGDLDw5wdYE0Ayt2vbpPsAm7GdzMDUEfm6BE
53UluuuwPnIOyEKoRU/fL/AMvqXq5LZ/ZWW7mk+ADrKH69aLXbJSer8tKi+49zdBKcVwsmr9pskN
sO4HduVoc+xEebfX43EEkUBhhdU+B0Avnft+Fwj+n+CH/yS73oFY8lJZCyvMSay6HKAV1f8tU/UY
4xi6CsCq2NbyqREM43lgo/rFKDAZ5ndJeOXefN454nrZB0LCWiBSt3ItHMCQHjf9tyO1fkctYUm1
ErMPiSBcRpa83T7lGejiB+kYXZ3Q56pIBmMzBTHtT/JVkGWcEmH3KA186znVYhel/r+BRSblpLxf
hm1w343BrVbVzCH7FB3wVBuTz7cjrZR6OzlzToG3MpsjljryrIn9eAJdEE509wPsMoAkpZANXspw
y/JPyzaE6f0hwKRoYI2r8gyISO53vnX+ZN/9oVbvDDaZrZqxF3ZwXL+PbKRW6XR25VC1Z2gP926I
zmfiWj0LMVsUcNmgQ78wji0SkNo/Mk/6HoQHe72SnnnBiMRf2oi9OuUPWerMz5xyhKE2vkFRlfYx
lH5uGmZrkIx7eFVzfELRo7nCniFMWMm7xWFsGP4J9X7F8UwBuZwdjOVC3mI+PLyNCKuXZtND9Bi9
1ZTFoPl1d8cCDkLYO6IuCYDQJ0qyO8vM0igj5MEXPSp7ErwL8xm9PEV2WlwmL62M+ifc003ocIUA
qX1BDQ3+1ldI0KRvwjd/5HVMD6WmPGoUx60eYJAKYV3G+Mh/GvrXR4xb9eEB/LOEhMSltDk4elhN
UjaxczokTMqucESqWB6h9j7vBbMvX5oO6FJzNsx1DaZyqDRLppRcCkss/rzuCmUiLAe6lUyFV0Vm
y+xTXshpLOjmy+OsIa68IpdMufWwGZNYIzmIGue8cI3iDrRFtGcvRkFUMMs5H28WHaZ7euTbwSKN
cWBNvSTIKBT+U2Cik0/6/aslKV7xjzmHpMxCH8xuorEkpH5dJyeIC4PCRm60+73f4LaW5UPdU/nR
iAxjLk5ZLdtz+qPWr7+f9fVM9CDVz8fnUDpPaFMWmSC9m6PC6mazhJix22kH1aKMI7nJCFmNfDct
H9o6NGbuZ2hUEQLBZgxWSRhuUhpEy/y9gRuREheFgPhDAMIZDhmOECbpVtXp1EYpqKS4ca/U4Uj0
Lftr5tBbNwPtdPcj6kAwr5Tcvb+YnBX9yV7DlXq0IcK9aG9719JDm1DJTwVJKkubauLiZiFGL6ji
mgoFmNTV8wXJ2KaDnDj404z2uLm+2W4rZ8wvEp4b+fV+652bmzy6Dp/9Ihg63gFrUmU2Q2bJ5G/U
d4FwppATz0UHbclsxM5+9o/q7HkFDmnD5JJAHSAbvGZjHdxARy8KzE31q6c4vfgus3wzpkS7Z6eW
Y5nQQ1n0xCXB0hN8k8Le1TvQIacxJTMGsgMpUUH+H0oUoNDhI8Do/Rllm2ogl/0tKl+F5X0ktmLn
duF7kXg62I19EJypWke6Vv2LgFNSuJgkxWO+ArAClaS5eEvvizV5TMNSde0X73HJNqycXjD9EU/d
j2yJhHX0Sza3vDbVuZKHjnab8jKTnHBASyryY7e+Be7szgifcYIStf3ynQHevipciwMRqm8aZYPj
LcWnJ2xKX+Few6k5gBaW3hno5JgoII1wx3DsvOVlXyiU6g2FDS0zvJ5Oveq98EwjuVVBvpV/snQE
9o6VfRVuGFSUBoZc/51nFYYI65rIkVUIXsbg4WUM6l/vP4ZZSl4P9swYzRqjxMiP9PtlzqMe3G81
BXLiMucprcMlSTCMU/eaU1xphdt8BOQ7x7GbbHRrBVYeZtj8hGVcA5H2pniVIwIEu5ypFYv/MzSX
BFcFTzKcP4ynhkTNXZfObHwnQVT6eQiCDIIhaKacedici+sy5L2XysyNm76JQAdIdZMZYcXqYFGC
8ckuw/l0bPz1yDeb6nNP6IgGyRY5KRR94C7ClIRg9lh+2VfGysK+jpkBQ37W1DChRaLkDZqv9MI0
KIwy72WyCbfnc1g347wTYB0YLq43QjwWL8FUw6/cVsSrFNsfZpY5lZG8uQ+EkeSDW3yXjG52vcn5
KPC6D2yiBXSxmWOGC90ldl78A85sZtCCODQq7nbkWJKA5a/eA84DlOuW8wCrOymPhuJQlfTT/r3u
B9oFNE4sYX0HjnLXiywQge/tDaZwcd5TGRCh+OBWSRD1PR/2vvT1n4wirPmXH0LzjAqHphMC4YBR
Eebc1LJvaqsfImzhYAZNn0+9+HuVJCHV9ftXMcpci2/JTEsgTV8b408p+ahcIAU8ceHEJKzi+Zul
X/f5wVAWVNXTIYe66aPol0s3Jd2N5rKwm2KXztwVOqVottSFfnZ9qXgiDPbWZ4VyQXWdXCOiiAiv
I1xcxu7nFRfvsfmlFAla0JKKSt7XbRadOaJ1zkJoUCK2w5zmTFYPwn1iURkrSyA5bEHWvq6uQczJ
SF5lE5LCf+tCzLBD5IesRjC8SUmH5/FWo0vdK4TT9JfHkHvuOWBlqweU+1UxN2PP8gabxSovolzi
lHyFY7cnGblpaPFPHUusU0mZW3Fhw8SE8UzN/kFv9r17+H4nP1gUQxQqs24l1QlzDoBSNqABXSdm
85spCcIh9xnIzsE5SlTPLQIZFCH0QD6viia1dU17MCjHdLRxSH6S35HbvyFiNkBVR49wCfn6QDMo
2tYE3d2c0e6SqCFfCEJ1zigqdHuDRDlG/CAxo6cPz1GVY97L2BjPT0ZCyZIlMpdgLwgBb4aqXfY8
u6ZXSF5hsqAMTkFn94rJ4RTKrFghgQ6uTYAsgxrYAblRWf8NHcEqi8a5SGlk+zqJNnEO6jesf0vJ
Gzza6Voi/1Lwcu0QakM38Lm8w3qh/ruk8qBgkT9Bt54TmRV5BI5zxWXdq9zqH4QMD1LwBNAd1rs/
Tx5sRlD2zxnDQ6gQA0nKa/4M7uf3Q0YDydPyPqQJLm/yqjxDyxHga9EfAuIIxLKstgL6GvjoyAOg
PEfkGqbBLmXmV+GwUrFelZyLdXX0fR8aGxdixmHzC5nLBDdwcafyH15lpzulPSlb8yp1KKE7GBIs
6NUB470tw6qEu0D/eSI638xdAyRFTwbTORirt83lH4kYOdoDleBNdb5+frJJWQL3WRh93t9irq5s
+AHihQ5p3ggtzFGB1R+IpbkEFk3t4zWuMMqJ0+iVcHCGjrcTIICCQPI85A/PHBwD2mWx6tPWfRc8
Vk9ZhLxehUHCFxe5gqi8v3csAq7RluvC8u4ngbuZ5MmexoaiVm0zVNCdIq7Jy7reSmHgtTlZq7gk
V1xEmKyjMuOwdKWY4GJNgpbw/1QImGg5oPJVMz0LDVS1xPtEpJw6oDhp6PwkK5X/xkBlqY4gnpSu
pHKRF/acIb7MTuvo2EF/qmyBwB78Sut+dOeRB//km7r6eLmvfEte39L/4dkRzDaplwDr58bupwMZ
IYHWigmOD9r1TWkmuAnC8n9d8yho9ujgiBo8YRIFp2kdTeHh9Nvorr52ze6cmHQYNNGNJPibSFNJ
U0ySFRF3Bi/n0qq5Lqsn1jroNfsqR+hWWNXwZBRcGzWc11gHPnBiHT3tMPmsQLAjlmbyD9ZZWnxJ
3HQqD2kTJCa1wMbiwBvsfTH36xYq7N5sgUzHi9m8TE0aE/ioaLswEgssHEiU7tnwd+YeldPsW0pG
sVa9ddC02grXKGiLxiRDZca+jclN/phmh1oQ/IRo+H5nygalmx0if+CACNgzevYQrQ8fqgaohqlN
XAOjnhgOADT4sEbA4aGvy1GOU7iTyoueqFYE7r9iJIL/K3gCoKeiVwV2X4Pq0ubtJ18ccQhI+T9K
nYmdKS12T7wYTPeT3eIfOlB5l/t+85DNeN/7bqwZ+OSyxxlK8vXVz/AjQ6+I//eh8HKoQ6Wa5AvG
pCaBGbZhylAIgHViX6vW1m+8ooDsLsdeCJWepfjMvHRNmR5NPZNHXa9ZxYa581pb+iRmsZnxSeFB
Yxeohz72zSe2dge7cy6RhKi9pwjy8nOV3XiMja0znnvgqPUNvJwslPrpzngdPknuy0JGJonP9+dI
jH2NV8C61+OjJYo8Qe1aySXiKWZlFXBU4pZ4GuZtmtdRrC2qtv+NaKM7UxmIh3oo1xu5b7gqBZzd
KvFtWFDXcj5BpsCF24VBkvSiZVr2rpmkFszDpt7tC5xZIWGQXzIaN6Is5FiDqD/LjNRBzZamfJje
GaRtM9EcaHP62H1diJWbPLnF1ZRqY1yYx/7ag10IcBlB4+s1tBPE9CMlV9O1L/4ci5cqN8NL+DDF
gXDQ9n8IigKvvbmHIDNcy3iw92wp5eWJTBk8/RAJqbX+RyCmdB4ElnJwfUc11k76NbubbTwGowmc
qajz8EtXHH+2qEGVwOtSnJ5Ku2d/0WK6maywILQOU1E7MDPIZ3fHA/aD0XiKswduKkBbcBAksKBl
cHnAW9oB8/0/vzOJXv99o8WWiEDdvfnoj3GKJgHQIBTmI6FfK3jHnDYzVYL07vPdRLpu0j0kW7yw
fMRqaDSckX0vdTajppPuCs1t3udDNRoxKX7bC0kDHXAhzzNNIWIsRJNX7DsAcbRIIkAb763Gg/lC
ws0QLFkBm7z2h7DNPx4xdAzbAsDMA6qK4oySsLHkdSvfXLCT4Vg68fUzsCL4Hg+3cr91LY7K/PeU
C0Axw7APGNxFlyUDafxHq3OjPumTwlEF3sK2UMBfs7RcAKPGPUgQ7SdHkmOO+HVCqVk3l4BS7KgR
sQb68fR0H3lokBAnpzBzfrXJajlaDbnbE+4YqgGwSgmtv0MAfI6o0DIXanl7rSVMlInU2p8w8jaD
2nujMb/xA4yCEpiHsyAJe/hTLHJevBNMwEznsGDFXLfYIXv6FE5qq5EulOiYcCva+qqojnN47Zon
QPfu1Q69V6k17HV5pazYOKfEE5Qo63F8YN9UlVwaFXodaU99BbNvajNsGKeIwC1OPPV791nJ7rpk
Q4cyStZZgeTz9602rNyD5hZqKnAEOZJFk3FUTmtKYZCnyy02pxVh3U+ptPVVXEu0XWwhQBgMg+Ef
yTQ5DWgR58RQ3pG0E2ock7SRchGTRqvqZXOG+y8UNKLOShjMqKkjDjL6jbrrsc+ufsFOPGdHapMg
jIRi2xcc0bHzWz+AELiYMuKSjVarB9yU3YAcZ5A1WS3shZCRkA3JmA2VnqoUqfQ/tTYgCI/83zVg
aw7v574MkCmqK6gwt/5aR5kFPbQ/FB1H4RNa27QOpIGdFeyqHc1W+3mUjT0x9hjhWdrQ/oadThH5
BMU/cIkcYXbVAtn9xQNJEd/KKMfBBhCG+0n5KZ3GcSPudEd2HyXHCXhUfXyOFFvbXN4b81bcPmgm
+bvutN/TpWMR/LCIZ1XhEDQNs3Jkimu9mxk0DJvK6fovImzW7vKSujbDCScwvADtGBzvrls3s39N
zEWFwzeJUrvx42p9Jj9mQf/dcS6WmJDU0vgmqS5x9MbGXHdHuIp78rqQv1wVCvFbeC8zwq+makxE
XpZLvH9KfEQ3MsIWJstlr5n4zPQFxAv/LFnBY/b2ngS9r29gGI/SqMh5XSVBtRbqEleVEMI5wDts
1rvcrS9oWZLF+93aZDRdonLXCv494g/KlA4zb8N3zamD3Cjx5rJoY5yeXMp8+bwP/4esPqhUTwVM
78uvx7o2rmkDVO+SijPWYhrvQIpX8KhbMFmJB7nl2Kfu3eqKucwt2CdzyTtHpgHV7MegvmPr8L/p
wUUwSR5XeYiLuHrqNJ1z959FbNEOej9Lg24w8z6S/yLt0vpuKhaRIgrLKp/lJIZPWqpa8dd/xPUB
ZAGYkia4rPk5Hbzrq7a+9nzlQV5X4lHSF8+ETVCfLJnyfcsX5kXdHRvYmyxNiUlgKjfwZVQ1zTmm
Qh1ovnVOHbP0MBazLlNKS2gs61T1DAFJiFGJ3x4Dx8agfC5EkeR4YufMXoUO6GGkfJtDT12ZpvDf
QRCf5e8Mz4VBS/HDtO8ONyrDDcVYd3zcWQ6/glxRGWZr5bTRr8gZVf0GbHmg6URKeW1sGb47oWYB
K/1bQS6F+A0oI7e8zVm5CQx9Csv+STc2M/zYt5RkSq1Amr/tU0/K4gTuj0dThRwyvraJiMKK7gvw
WCFMPCMI86CxXnPdsL1dezsqMh6e/Z5fSJh0u+TWUufuBHqfgaaulojFiEaPf1JDgVrWoQXxfvZN
E7bYcguTXUZNr2U2pA5Z/nhBViUzWiQX5tRI6mvp7G9kB7pUEQrV+ugec7zRarPvONX7HPnYtnRb
5ucpXp6krtG7aICJ6lzoESAOHundeexjdA4uTsWa+jtDVXremZrfMsJo1tgOIupZwVRSLBa8Hib+
5AZaSm85Rx7RLinHTOej16uyTe21hV7As8ek91y5Y0RSyiaOSsc6UfMvaMDRKXlzWtoKz8xsguPN
l+VHTPvzEm/bJ69HW9KU0Ynabihk1Aw/DvOMFmD+Pg5TqL1ydWgVpd53dqpacuH66Ia5Gjpt/Smf
KbCl970/A/M3TO1tvIekQN4iNBhNxtORZkY7/7N+RTObPByih8B6Dvr3N7K4YQlvgOVFOAwVIZp9
u0OZCJGvkCzfJ7GHX37Qrtpj8o03otobfRW9L/sTHPZpjU5/wSs1/QgVdqIJwwoELnUj5xE98MvU
QAB9DV1ETfMcmG5Jfme56x4IPbxMJUpl2eFhxNrv23li2D8uZVunPaIv1QjxS6MXMF1SK45o3MkA
tbEbVAECgs5wBnB+ENDZNFbEUa12N7lwOOd5ewLtfs/M2Qh4nUyYPikTl6J/FiJmn7bOeqXmU+Ra
uKobRYlCHpYyQmlvRG6YnujOfq0gDEYEc7KyDgmaPFKM1eM+YNaoQgCCrXgLTLIn7fneSZZxKsfR
hET37XsLfHrsA474onmMdqU//tOHunNn0MWL5Bji8eiohg5bMWzmZuYpL894oFvRxrrXVNtnaHC8
hLsFdAuT7N/57Eo2OcGJQ7VU01Juclb2E7AuUCaFv4ldwDtlsX9wA2cI8bWoomngAvsTuFOuX5Y7
oNIWqK862q17ibc03J/RNxtmmYCY0WAGMQoZrVGyce6SKbBHsX1PtlSIyzuvs9v0K1c/mSfZq5mA
NQczQaUzRLpulZDPcGjrCrao4GZ6CifR70FzKb6C/jS4hMz7rmYMHsm943n7k9UqmBGqMyiEEYe0
EaUpSctCfdQ9Q60yYNQzxCU+9VecDuY7YblQY2jOZcmhZ0KTb7SD9i8RjGLp+mEtaaG0VFmgZYtA
oYhXjWUX6JKixWKWL/nSMvUfLM0YQaEy30jMvZINHDvJMu01pyaRnlozG3t2xhd9bF6QE4fWlT/C
/Zak7HhRH4tm6s3BRJGdRyKZ+sqnIdB2orLbEoX1ogdZ39DITK6deA10od8ia8jqxBq6mva8XBI6
9TQnwtl2jjwurm0Ppmslx2ghZk418/Q/xrvR/E7kjbrAtlkutldiipmQfrpR5c5dyefhipdbnnRA
yhVvlcE7K7fwQNhxbks0SYGbEJZqLBjdfJNRyV6TVfWfkpcFbS3nDlY26ryyOtzrzPhDfzXqafQC
KCz/i8VUAbHW6uXraJGuZt/+QCdo5iQT+RRAETlF7FdTNDvPqSWZJnZsi+hkJ/tQ8zXNoJK4qh2+
X8XPQfRcKLTX66meF7XEKx2v6R1joPk+Z6upoB7s/WPCrmONj/B6zV1guTID4JZFfKRgQ0Yw/4dO
v8GFR+LsGGurCr8ZriUlH4ndxKZd8qObnpZDsmeC4gIQm7Z0FOWTsR8KHy4FDdvnt9dqQyou02cH
io8Ow1ld5QbvG5qMFcbUwZbUEk/72ZAzn6jDbC9wl23jkCpnvqx1L3YT4Eh1DO2NErg7mldeji2G
7UlpxPLvHo3VzqrkOPMdYIHo8RaHTv5YcPBhebG9Lg53anV2WGPRnB7vGw21wfvQkG10qcEC28Mj
nr6MU5CDeWJRDowuKjRh5bwpwbSUyI5ioDSxLnscmeHF6BD3ZZNB/1PhsFgaHlpz4r3wfejgY94r
l1GaR3c14jtzcUSO7a0C9dayTuEAwLZwvZ0VWhuN26sume3JHejRstVjcwidGXQdjPUr/WrlfLbP
zzeQh9If3qV6l+QkfNB30+A2HtXDFZioV1lOiqfO0lD18OFXcWYeTKoFHYMyHiMqiEll+joKNQsd
c/Ykeaivb8HQU7wc5GhIMZKYwjX3VxMupJ6F06Msap0Abthbg8jQImS60hOUdkJw7lZs3Ey4QiMv
mNfQosez4JE1KBevwlMw6iwCSXkomU+1FNE4mLQUk8z+1x8/+r9rbRjv+XfMWnyN8+X+e1oN04Kq
8cZsZwf0WFaVE5JMnqPGOEtilRBzVHLmuWyqbEiDdUdVh/MPPiOTLsSTTz93xTZIgM96QXUiOkf0
wMm8F72fOeraRCs5Y+ABWxpgfJHW6lqV2y7acjJJhgLs36yKynM0H5FG/fnmzmoXjOF4SvKL2JVX
G3RzxzU/zqO9gsuiPCzJUamyGoLG5Be/Jdbk8IN6Id9aFflzjfyMbOITc7ywjyHxD3Ir13Yn3Sye
2eZHUMTBK9w74RZHZhIrMclpOanLE61+XGOjC3srExeK6YE/IC9XLCp9DenXLldvi3MYuMwuC0rc
DcfGBRIz31BbcVUkzBZD2iAKIzaIW1FzAGLxKfA/ZUmkY2UM6elAA9pWwIYve/ecFUVg6of6P6Un
rGVOGvYveunXzko2OQoFTLhbsQnI4ZMzPgIaXFplUENPeMEhzjbQJe8OPLvwreHC9tatd8DGu/gU
X3OIuWYYf3WM+6zH/MShLTtzZrfN4Lijwgvk4N3tEnT9APXYLeAPRpQwVCwpnX9doobioT1jhLZm
PpkhQ5dTRrg1uvfLzFn2dXhnb+HXW+ppNp+Pe1IlrpxM8eOKS7RmCbSZ4kcKkjo1OkUuyrqRBOR8
BHzSjx9jFeQVySil8lh5s6gMywxfi7Xh6GO0LaapuGIdWgfEcaYOavkW+oUUqPu5eAhdzDYN4mGr
4HhIISJrY2aH+kovstDJ3PY5JD8DVIKpotFdZjSwOxpDcJawsDFHAjB2SnWNswanJl6l7P4QqI+9
d9Yyy43kx/TQjEFviNg6ipl8adwQ51PyrS/uduTAypTy6FJRK6b3w8JgxBg4KLCU6AIkXAFhzblD
K7qY9PPBDFSDImn2wZtKj/STUqLInZB9GvjUrcWBh4Igc33YO4AUXy790DW/Bs7fxaIwB9EEKSCo
IJk6LI7C0agpMXq/tL3Bd3SC09/TTjhS6qguQrWMqpwAKsZggezSVDBMhmeWzL1oEBYY9E2Kt+wQ
w0E1JjBRtA904FKf/VQ78hHMMfTLHVJ8kJITgooHM4zy5V6G4A2iA03k/iJv7mlwhpRj6fgOtAn3
Rc6bTzy9ynJPuYJT4xQx+CUoSY0O9aPop4vw0YIoMQV8res70uj510r5LkyMvRmzkO8lt2/XDpd2
ewSUICM15pprK1Y3zYK8G4uqJGxBS6SExOGqEYqyoeryXrAzyS22mYkBY+JmSR3GspwTTR1rqNTx
Ehi0qpeRUMSLIp4A0IOHniKLIocUO2WPH+TvTx4b4Wn2g4G2la87BrGbboNbNY1/4C+SVgkvPFkQ
54QlgbTfu5dL05/ByHSRu3PfEj40/aPclDCQok9Dlmmd58TRHA8aeCKtm/utmGuITSqkXZDBRS//
/FFAqcwzs4f1QaT5C2xehkpr8LKx5FfB3MaMCSYyE64UDiN9fDcTuSgTpD0o55o26iL0bV/dty0K
PQM/f/lxJMnwwTzwXBAVbf4qcy6NB48sVHiIWrK0mx9vzVsCw26hX+p8KLvTGXkmQtgFpGqiLoON
M29goqXO9LWfqShbFTU/LQKg565W8MDuFYsCLLc4KGD+GqE4SGw5sT0f63hV009IaYhtjOwbdw4r
xQ6lJzhmYPLvBbAAsl44HKetbuziIPH+nBs40UWoDXmQ0fYPiyowx2RtJ7iIE7EvymmDb9zhDhXR
6VvyTt01APQLmwv5SZFxtL74gEqRiZMao1oR6fRl+tR0eqKNl8qWsBm9GWj5yMto53UWONro/bW7
IOHKK2nu/RYdHF6V/XdcktWTUtyqrZZh6cqjUUUdEARA0r/+twMGspgy0OJ+4n3/yVWWmKWsk9j5
hIqGamNb6QplmKG2qBYQ9Zvg//dKfv4N6KFZk10h+6An4O/UB7efoM2Vq1JMmfe7okSVxgHej5y7
4XzIEZYnFeGXk82J4KkctunT/jM6uPb5Icxcc3qxmbQFOBrSbrhXkSxuZ4dn1Y9otYMtLfFZKQGX
iG66jLS7ME967V2w3B4oIE1WuiWeAuYZVzNdPqERamPlB5wKufodBECoGVse1k9PXXhmL072IZCL
UZpvblltGf1GkJ5ooyCNJj+Jrob2U8BqMEAO+acGRS2gV6gQJFpHZ1DiS00VzvsQG032gY7nE9w2
pe2Jwo+ixdrN1DFvvySKzfFKt0McOrFM6IpN9F+OgnELm4F1KW/ZAgYop/5E8FwzFJn7cRgaw9nv
jsgg9Da086C+HXyCZ7cNIFdwwmCTfRhRx7a4iwOSIvR+dDuwMmwDCQlOHnfxHon5AaedZ5t8V++5
j2WR1KZSh3p1IrTlu3X/CNI0aMfGRoBbEqGW/veTnjGTzAEUHnLIsIsQXcLyvOL3gSlW3YzHCOhm
lGUoFg8XEI6JMzb1hC2ellT5kARfT4SXX0bPrMB0CzJKIMgvbRKgiDNTi6sriGw+VNGQWqIni4f8
dYmSj4s1y4TuQgqxfihweYb7wbnbUE9YZSu+GxqnViT3NyLOLUmLCCg4ml4i9mi7BezNPkNKziCv
5UzNdNgmQ3YpuzVMubsaskIyum1kTRmzhCxrNwk0V5vIYJH+BuEgXxvQVqNfXqMYV8Fjo4Pg2kwi
veEpsw0/3BvkF2Yr0LwFZyUaTMxo8941Cvv4SHsNUKr1SMhoBOuTxw80OIlncCTb5JC2lbk/4BUl
bAtyYh2ombkXcl4CXcf7Ny9uHPbZf8suCYW+L/QV+S8Yn14CUjXLD+JQTHZNJw+yPatcjtzWK6id
uGOsDMV/5TP14SgR1P7cCseYCbyyKCEfGANQO414pfx3GHn4Fadc0wUB4UWxq2vWgmK0x3Nmb2SA
1QDIk87yMbkxRY72MYxRRreVpDLGt3osaHiLJgEP4gtStzZu70PuqyAEDyFRCqgBIsm8S0AKHAMR
FnEXOrTgOgbH7Egwrq869s9Rqa/xhtPHXzOqpVncaAQg5wRwaUsmUKO+9d+O3VosVtYlADL2JBh4
CD+/0t6RY7cfCiAyrybFnOqUPDBlfO5pBU4xbQq7YH/koaD1KVctqB9GJVQ7E9yM3D+WCk98mtXt
Rv8GzltW45P3+30dcPVvsfnpKfZml/F7GDQtb52XyqSGganU3QcSzymL8HYgUfSMqo30Ursys7En
kw1WFAYEbUbrqn6WJOvd9QJa/B+oh5IGGNNiUkV1f2k+TheXv3nVsDhNyXzpz/xRZrZhIiw1SwPd
aRasTg/aao6oIoZS+5zmX2O0s9SP4FUIytGth/s4lqGwAwWtw+7gc8yaRjE/SNj1jAH6WPhBn68T
0v5YUMiTK7Ve0vYDkehCa+7KxC5jAKieskpdSTZMiVFV/RZ7gksVgPh34w6tWkb9iA7IJrDRnT9S
ssuSVkoRBk9LDqtx6ejMf0VD4NvYf+zhGIN2sUnUk6N1m0dEKQ9R2M9JL21sQFVkltfMXV+d7uP9
uUThERHBsfB1zG6rX2whVPlLvFVIulzGYwSpW4AR355287+PRv+ru4suX2lDxHP5k2gYuV1nXmaw
Gs6rpXXXarAOh+xBzBZbzlqLu675CuX71jNDSd6rzgZoqSX7axtfHKb5olTW1OKaNpwRsahD1wyg
e3I0OkCY8CaTGVlBrnUNUgZ8y7BoZiFvqrZpDjqbJfMHqm5/SlyRjFeI4l4aoCGwQP5qtoQzSOHr
XqFcf5fa5CbnSik16jBRbKiLo8y+pFC7E6QEQ6L6QWAotNFMFPxr29HIvtxEC/dG+kWhgzrztBYH
HXIxwkmV2eKUP+lNM5Lh52iqw5TZKnDTfDIHVoV9s9fnABkQd8iBiRo3D1YS3FJ6QCi5dGPfJBzm
OIxxzD8uGtq29jf4wjKMoi06vAGkkgu63RkR7c+wE80+X+X9htD0kqKF/KIJMxyNAmM5NGEe2b2I
QYpkQbbsU2OCp/mdKaFxHCSjmbke37di3KWrXLERtKRw9w+U+1WN/Jxy5lSi02GLimZd+QZVBHM2
ZlNg3X8TjSvv+H/rtswrGgEdrk9gq0pmGY0L5ugKa1qj17fOycZSk/Z8SMg3tDBOqDQHlD6OpJxa
gw5yLswlyEDlmSvLLupMjEt29/qYFNIZCCImAUxLomdxsBEHr2EOz61cfX6ouS21RysvkKx1i9KP
zACVOkmIwEhedtA4cyzWEktdutEb2MKi0kZtsLS905Q9v0qhC2P54pG/y14ZGswuBKEL9q5fjvQg
vbxWvCFcTFdmeLoiQdKgMYnXMJh6c0UpQ9CDQuLUJWN/KFdeFVtciNdNkfliZWyUy7lv/+lkQORC
hltB9LFBOWA/4HQ8707KhO0J8GU4a9vjPrfDbSSf21x+GN5edjEalAwLk+lh3MCuQ7xdmTEg+W3O
TyHVL1j8QLcFCh6FqY6jAl2KOwuf7bXQ04auWwni707YdEJhak2V7NsXK/gAlyzCMRZn7lahIKXC
thVd9hjOQVuX3rec99SvKfIibsk972sNeALOpczNSyUMKF1FBq1Pilp6hM2B2WCqFtPBaRNeKY8N
hZoC3NLHwfMc1m4Us3A5RDzT2C8n2HOz9q/YmTG2DqO2aN5WRdpG3H2SnmoaZa//HAMPpLAJzHCb
tK57zRkv3OQh3YQKDG3ZAIcQaGiKFEwUw4UKUUKBec2ZEwPFPZF3N8F7uo228w20Wm5aUNcrEwB+
KwGcl6+982S+I9mG9yu+9UAwwdvncY+FusF76QKLjZl40MWeQgvhhm1bEC6/ikubrdN0HeIpqhJX
RDzLN52TAJ7A+mAi+r9I+ibk4yqj5yk4A7qxAl2NaQUbniqP+m8NWOtQoEmrvB4s9UTDwE4P++hI
5uuq9WbZCgcsNZCmI8yRS5Py/rA07XT7ulSRnoSQh1AP4p/z7YxC47oNFn+XIY/XXIPvjlyaarQ4
eRosjKshEOcl4QEXJppd+EveMXDzhQpJBO1UxLPPRIJMijtduQqs63OfzLngSsRNNZyXJvX4j1c0
mu4fEEtKiyQUjcOHUaugnF8EQrfS/DDO15kiRIGJ2ZJnKa+SaW6TLBmEnYoFMHc28LoQ1g+xysc7
YtSZtBNFMNBtpRX/bSmoLAoufseR7xSTHLoYwVFaEINJxcwUtbf8T/zwFJYC4OQG5OBUNjOwumry
xEF1BKCatJ5BJXFLg9uvqww9g5Nt5jLkoinBLWFWM9vLg0K1sLPH7up3VvUqDrpRfcPJfK+EMMD9
ShydgRovReq+fjugXyHnfkPoglmVk3vV+MRnZmjZKqVg/f55kk161gD3DuFEiix690kv5pxIqaX6
JxGAk6l55rPKEE7iGTvg9pRR43QqKzK0ibdQM7dHYC71aCMTGt/KDnhBlLrIj7yR2g8AYOw8kbjS
mB6GP0GZ0sPdjYwAPPj57mT+sXSPPVpvI6TskYNtmofbcWqIt5oMwq4UEJXEF2ICpcp4gRffBHC5
uoB6FUfofOR9pe0LuaWo0GeuZRWyOyczGMJLjldZ1uUYGj/i21WuQETqHqvE6B1/S5A/6E0PKj+p
uF2957OY6qR4uUVkOb4Y+zdFYJ1IjMV1GQcdFq7+k97DJSFCNFt8+fQ7/uMo8Dvxp1iasnwSIZgg
UOJclQX8+90jdYnhBOMQ5kk+jTv1WiIM04HqScA1fYu8e2Rg8dZ7rHssDwSiJlltKYNWM3lrsXyP
gVV9vH8+ryXzndeeFqykkEVaCcDyzGvfWxzxBzTlPzVl7xIww10xNtq3lxHy+AgpA5tFmemgntZq
0InFQ45UQek1Z2+lGHh7GrlcAMT3kfRyRbtUM2C7J3RrNyiTlgXHsX2mqA4vcXGmBgyqWMa5gTDM
waWwVV2xWqEz1mjbbmTgGi7WuLldkTwBhTxNod4f83A2Sva1GCt+eizwLYsYctEKxkS1I7jJHQaX
wvoAJYBySLejlQqbQ8IhzhbYfokTzm2Icj2Y1l4uWTp5ZZp6diXXGFFCyfOWbDXKkukoJUgnGCpV
suDe+s9sR4hcisVzrWkdJswpPmmGPgWVK4Olen76bNiD8yZ5t1ppIInPnUTDkFofZ6i1w4R7jgoM
EpM4UuZiKnhvrXGDrwlJE8V4OxUn/M35GN52WuuF85HlOy7fgMAmXPgi/5HSTmr//5mHEBugXtEj
8JfCztMLI9pPo3x8PXKg5EXXHCmrUeOIBWUkWkOhRrP+U1c1vFMLLNTkzY2y+okyhvm5DPSjtpzD
myPGHJJ/FMlkdI2JhbsTH7ZNWZFqVLJqbLF/U+SOMuN53iZQcIcMcdVWtTLw3znHmQxTJ4evDWmP
moSDltL+vjkidlHeNtrYeF77Do7NxTt081LO1VqxcktXbus5w70biwxKOYM5q5K6UBIRJUhwf0h8
TCa5jlMxLeULtlM7uJZ+3xHfB9f+vHsNh7NrGl9t4xoQOoEcz8PD9zTOZTSKn6It/Gnuc0CqyAQF
Ri5nPzXOKZzGp9JuMaGwEx0k+uNFGAlw3pahigiWiUEdL+sBDYVOCjuf1AZDytDAgKIqo9tK8Ndg
CnuK0v67pEGWZlJdQWZ0h/FNoZJ9tjBLLQ6sm4yGiAPYtZsZgRVJE33UlVAM4W7+Y5xbnOCDSZKo
inzuZtq3V2C2sIx8uDl3XlOvwNds78ntPzsoecn+DBDlaDJK2atyR14Cq1sneGpoj5lzUmYnYXZJ
oprIAU8lBSqMcDs9lqMUug91QMwZ+kQVHRjhi5TAlRp86ftWX+U+0O1c6lUzdHC3xvL8PDLQmq/z
s1LDMce5hIsi738SBIESWpwFraxq6MpNrt0KLy27WJtYPrOqUMq3f+TKUZ0R69KDvfZzJsI5gHD4
uqtj0JxEfZYOCdiE8ed4ypB7LN+x0pxfd8kTbkqPz15L7OOvG2DTfuH2RbWLls9qkaDFmxjlt649
nDI8+eeD5RH2kfTisYufU7tk3SRi8R0Qykc9GvVpt6FI+ys2N7PL8slNhB3NJJ9g1KknUWHDxDHj
gK0zPBdefXoawRJNcgUViGVcjIcF1aRhWTzbOSPPIYuhA6QhPn3LOdXbWD4FnvVcU/LycOELg8xe
sx6TXTlnU1Hrrhph3dWkNGVFQi3RMh6V3ipVsIZg8uzfJjYL7hYidQiwrMPAVDpCDsfZPHLDkMmN
Lw2PaLZVvR4vUdWwq8hcyVVVmYCAOjhN8kI6gQj1H3nrleilujsErdnVWetRISOMpBELBv1m2x8z
KA78CgL0w+vg9hILoLmi7h7PnGcyAaKdE54SGldmAnUz3k/ApIIwmqZcAbZQzV81Y8NjBRck4a1I
0ADn28bM6qwvI4SimqAwY7AYRfNDv9IOVqCO0Ds+XdswapHeEWldFeCAEqkOgPX4ZF98V8OcbwHW
aY1TNEtNDbAEkRXBTCi5si9vLKqTmTxurovSY9HyiVUJfSbYJCPrC2MggObqU72eft3G1UqrqWZ0
5yol2xU6v/9qufupknv9IRYliRcn9xEHsjBOU+HfdWHOL+fcGqv9rgmoKzA2wI4ams8+MsgL/LYC
8NUvDx3aYWEagXDeLtnN7BvlEVqqurQMW2B9BfU7oJD00GClJqKm2uItpsDNmC7BppxOQ1npisfa
VBVt7VdFcp3snw6uektJoG6Egweh/Te7UWJBLrqW6PW8Ez3NpBaYyk4qXSgTZ8wgvcevPDiuVenS
1cJ4/661saYYIDMGA9pHsHvZoHWHzTfirDqcCvI32CDNN23RbaE33Bl6omYNKeEhjVfRaPg188N4
8Yqt9ITxXM4YX9gcpIBIhZsQPPVfHkHVYtCaxP5oOzQNr85vR6FPtZPdiPHM1ku2tNnIDXAqdth1
xvw+LkQO0hAMVFcArXy+H6WuMtM1bytlNGWR7D4S42kvqNIOAztcAe+w9mRIityUHuACLyA/+ROW
wIn2ubv0OqNzN8CQ8rnICt43SlIn6kfZaSezwW7PkLY0xTXCqVUkf04GY1kAwYFRnKeGBraDpSxi
+ipyGVPi3OktaIL8W63QeEeCsIlNUdI6yAgTE+3wjoAngU7vIo8mIsmGexaLWBJelnhRhSc4yJYr
kTm1WC/ltch62OijchpOdBtuO7RMHDYR0nGv2glYfomVW533HXOqUpew34Pr3NCVs6tNyiUpW4lc
GH54+2EM3UILX8Mb928fqUPZp4vqaVJlXtcR1mN2101dkzxppcIMEWns6TGdE5I3CtRCoMxywf4v
hQ5fPa7QHTWjrd7J/P9uFKAvKZv6OKA6oNaf5Gc2A8kBKbt+g0DT0nta4A3Bs2ZKV1DF/1eUChQc
06yC3/QZXY6n3rtr2Cd6Jqb197+SGw2+4wGd8HHkNa1ORVojOcJGwTY1WD6aHIyfonQG+zYNBj40
qgn4edtgxP/vimISf9aJXpK3bme1clf7eOwX84+bPmBpfXprOuMh5FrOqe6ZgbRGUUSnlGe92Ewf
gE902Fcy/JzQRYQukwmNMRoSCA/wgr1Pob70bb1a041LxNJVAm6rd/x8P+QO8eoC50OhyO0lQceH
B/ObLcklNElvNP5dzIAnCwIwC35cF6JH6ONHd0+lMok84tFD0Sjt0c0K5V9JTVSZfC1B546ME1co
wREx/S+rL427gm5gSKQIdUnIlauyX+7B8xvmz/wVySeYjOaB5up2oncKPgVpQLgd7yqWdasmI2L7
7TfRNII7fAi7Jx0BTq7Xx27HOM3NFZEBjDW4ugZK1pIHzHFoO4JmNs6VzdUGAJmwWmlhRnhGb/IQ
3Qu5l6k1Etta+/kOiETgVo7QjHiAdiJoedHrAvofGJQnvXUlG5qauDngPpBUZYamuWISbAQ7PBDk
ISlaT4nhW5HjJsWImoyqrhVQmWg9ptPK85FJ6amAyFKBjdNVI+pxuq/szqbAH1mBDTKuNehZqAKc
liCi4ooHLNc2Sy0IqTk+NgQjiPM/iR+s8xhEyMIDHZrpu3Na3hjUHAkC8cz9hQGcQTR2tcjP7vqv
qY7B5S1WPa7djjp8ylsYhtse905r0eAalyKzNkcrY2urshWjnsr4/o7ZOrc1l0SByP5hF84ovOik
l1/PYkj9g6ElkWGYUF6V26veZcF+W2mkCShmhEA9v2geFRS2PB7F3xXhp1vuE4pMB7CMFtWXdN64
l3D77A0gBs4c9i+n5rBYOyvFVvziHyfK/vIUbFSvb8dPVykSHGJCvAtmN1OEGV0pufg/NPN6VPGn
9iJAD85NIiWnKk6wnbpdS3o/MFLvzFP5surrY74EGo90YfxtQD6Ijq7bADlsjoBSw/9zfxCbRiJ3
kAA5g+eW0ll+u4ZQXVxcpcN/+Ztx7zFLzuOluSCHLXMR7rIbjYrYgSkO4yrLKnFC32Iu6tsnYBJ7
UnXhZEgrvIUUsSi8WjiErndZ6vCETWUf9FvdKe3kBaOg4foU9iEivgMHZfBuQhpps4O9iWnYsKUL
HkpOPvLEQgMRuqbrwTEp1n6nn7/95GTsA/arwW9zP5/2m6ffAEl2i4hJJh4/uL4NOM8ncFPmWXdA
HPxOE9YM8TK8jNr2CyIe1w/y/9KsjpPs+iICJnSx5Kguywg0bYrvo0p6P08UvFyJz14BbpGM0RkR
DzST+fQer2To7p2CYjWG0VSOwtkEVyu46vfMrOl+2zEyoWoKPkaWCsgLBLUPROOldNAyqR/vehOD
r3GPZefGt979oXG/5CFTjHZOPdbXKiaavo2jPjIU6F71Tr7EdKWZUNVu6lhzN4D9rlWDNwkEEHSx
8Y8zsHN6UrShPgPOG6yXzy0SxzBl65HrLbDYO3jaL+L0+WcB8oFHJffuNP4CIGfS0QPD615Y2Cnp
Kxz8Cmpxi89UDLR6iPedD6F2W+v2d+fwFNiQhIq4VQVbllDr4pxM3mUdPs0XpKxJTarXzMdzmuGE
Kj6OXZm/uTxfP+/aq3fqieKEe154FjBMkf9OJce0IKsIrrfvYH03o7SlkyWvb2McvSch5FOqskhg
0XCTk/fK8hEKzpb2YBLfM1u+PEsbHAD4nfHtowcDkIf8WZqqG5iyKPwFUsLREqtIF00V7Hyu7as7
EqoY2tiattCMsPbOAkybj/8ya099MkfsxJAn+NUiwnv6zS63fOyCb8DiDB6LbuIKM0+mocIP1UoT
UEcHfk/6kPg2WwZks8O1m9ALPTjRQuxfuBnSY2/ad1ElJRhk73VKEVRJks9guVhRDRsqSoJXyOuH
O6gSvTMCGJ/Pm5pwLENcaX32x7vsyQNwfr7q9mXrP3UKFx4sYIDmneIxOqs33o2WnsRpKAPz2+1F
ZKtMpnXr0nnIYuI8ruUq+IkcFBhO4iKzNUc6PDkZrx3tRS8ejazwXNmc+Bu2VMQL+HuIibAJkc+I
qjXLa2RP5J5nGPiArZX2YU+7yoheKBmeCv1X6UGrWKoTMDMNzHt3I1vi/5erElL5A690iFUURZ6C
dI/qfBYI7DrEZHYRvSvOekUUDT9iOnkoqs0+Szz/VZD9Gwislc5gr4oD0HAsVykcmVWeGDwJldJv
hjAqhrj+4n57JNpkiJo3xB+72jwNCqc8m3aBVBHeaM9qWnPLI4yH3iCbM+URHIbODedXYtGqOnoR
p6gi2Fy9MbaBichzjFf+tRDHaHYlgNDW8ufMZ7x+iF9WxWxC5S3j5gpFsmDbhxqUUBzy743ICJ9W
riQ4/9zOEeDxRjEh8OdX4PO9TVFRnlPkve3uwrd6D4gNnh6GMD+l5uWOoDrWlkiwvnkooXltM2wC
fCWNdi6QQDWojo2oBUYahqwApbUUe/9i8IreiLzrbyLVT2kSTJ6kEtGK4MrDk9vE5r50w7257HHL
lqxqQfLUPIDzmNlL80Rbg2UWlxJsSRwTdya3ocZfLNkHAw8Hd1Di4s8iG3GwUL0NRlVd13Y4Pmwi
h2JfpeY/mtdQWsdSl33p2aRC6OEC/9NxEQPXHMdrTT4rir61PovQkws/N9lSe5QjszJenBuZ9nCr
dtSfg4aOUhXnCp9oUVQnwD1rkdeMMH7F9/DSmhQu/7B+Fr0YnKcoJm3w0K3z/VUdA3OhN4AZ9RIL
RvN5AQAytkFwc2ynRnd7m6gMKSVWs3sKD9iQxfAZq18BBbzBgvhTXA/Y8hMUqF79/gigKorutLh6
IS1ukVVxQ047edvJYFv4rb1vCUXkqi/PfNJlySGwFnUrUaVej4rbw8pbcMqt1PYLOEw+cRTQxXQ9
4ubQhbvcWSLpJeMs5F04RT8dY24JBUfZohFUZQgJYSig+x/CWLSxyJNtMP1AHg0snYO9UEHgcxSH
qEPnLnF8C5Dwe0IIbLuGarFB6NdCvOXGtfASWiQugP8IDZ8oH0oVOpa9m5FIav/qpiyCi4LLLoPt
gW9xWwHfmQU6pZLyRyyTNJ+u0LHkBardoVWJcZqRz2qB7gSScHpeXdb+mqEcF1AOPRUJQdEKqIp4
xRJiFCvRT3xOEaNsdbvmEtzo2AkrYoUuNXusz/OPLLJE3RkVGaeDwBAbEksnKHj72pduCUF5BJci
y9Q0erzsaRBkwjs3Vx+gxtckcTIPo9hySc28MnU8y7y79iqBvVySEc/sRMrW39XGNlef91y3zewW
AiqbNlpG7PoeQ9mQjbF1PiwvlX+DlXabDi64HpophJ6RzHItmJmE8oVMwnn01/LBhJSt+uybUR0d
OIGuOPQMdUEdab/tgN8FcX52rs3kEc4nQD30rYCM2yU+uR+MQ0hcA6pGO1dM0JG4ofHxibn3GGzH
DvBACBT9n28XjQUF6IVv6h9jgM9vZ+5UJhDYydAzHuEnk+Sj9WdTMLNjV/Ok8Gxp6vzDulPCnysj
LsBHsqbF2QrtIVcpuqcle12j6AVXiTVmHo+12FQSIuJy/jE/kVMrcKjH7Ris/id2Tp0g6yX+28xg
ppHqPYgGhiFIIIQ6MANBWnIDbIn0YY/HnZCmbQxHZa0/mc0TKgLJZ+F0s+v+6xM+fxR3029/KZny
CjbhCRLr7HZlTlqnsv9Est19j+kam4DWhCD5SJJPujOtE/9dQ6cHs8v+EzuN3Gghw90aZA6qdYUu
AHgGEQZMGKbZNPWPgY/46A8ru5N9dr+bU2BSTtlHUoM3vT7CstPilCgoaw09aRHwvjrHiv1HZwOF
8TMGMycNjF16NsJ/wLmfXkX4dp4I+5qpsn4c+dNy6r30JqIpHScGHkIq1zWh5b6mUfXPhUnJ5CHA
fwKLUazhFGZMtYvHa4GblLJbd8ywrx/i0ST4KTic4o0Qq7u6+DsTSjCmX4jgEXLrKq/OA9rcqK+v
FBM+JP3hR7xPYJp+9HXASkL3FfXWJup82sMgJU0/+H0IJHkl8QtMcDVDq5zFvxEFQ2C9y7KAgtZl
8XiZRjyahWVLXTLuU/SZ9CqAgUwi6Nh4nmC+4o55hzjrvQI9N8CsUvslwP6WwH2mVpvbD4us5bnY
VMHO5wqThSDqJlCoI/Yntuv9ia6+XeoANb4FBpWT4q6JnrYT/6Hsyh0Bqy/q9XvZYtVR7E3c1iC3
RJ+DjZjDyzBN3uBLE/dExUpA8m7yqNgG88z6x5UxZ68HYbt3CcbzH8Wr7gHFyofKnDtAsNYZwP8+
p4ydWSVpY3HzRa4+mhLNvbHJRUZvYkBkHQAx0nKDYAjJGNaRsRYpLrKn8dfEOzNHg+9Y1yD1aKsI
DU9MOHRjHlHBLdx1i5bk1JmHVCqjB5OFt5Whs3ybPZLj3KRGG/xWCuiFsOgx+HjFQR9vw+0z/2eP
yWVrwljZFuYQwhHtuWNj88UQuNFv3pbtwYHky2MlwZ/Oxb4phZWsK/Y4XttkCH6M4SSvbB08NWb6
oQYXx1U9rX8ta/2cEDMCQcwDgQJFQlPXvKE18QU9HQAFEiqLfAVnOR0RXrEAM+ARCz8A800KKNjQ
41OA8zvDZVQvcZBiR3T+BxMQmY3x4DrGkp2mSBJlp/gp0naDRD2ElK5ft3/u3rz7wiekH7YF3e/r
ssFKXi8XShnQz+HhjMjSMgUu8PnojlITiLdxAn0kJQJL0lRSCVPmV0fBA7l7z57unKUOBUKkYaSr
bKywhLzQJVVz/uWPi9fHImrgUksiGbgBoqyw0bjJQmDlN8FtHsbmAg0oUOGpI0f70Ui9ghWi4MUr
DT/tlCr8grmi0xsG59PLikQfH85UEuHBd2AhdfOfg+ic+80AoJpajo5kHq1Dsb0R7XtZooheuNjD
85X0ckzqZJ/10cYV+jeVo246nzwGtLIjT5JuL1EjhyEy8bMvJMcF6tHHehxFz2P27kjnxJ+MW3GP
9cOUi4U8u/Z9UARFTKvUtQrDwEAAvB+Oi5Qo99BgePfMLKK8i7jjniGTTZWAuGfEutzMayx1f0yS
hqfBGunW/uvMsEnP8qmJwrRkguMYgwMhLqRBJHphv4EI/97edN8qBdmwnN1rgWFyjlET7G18h2WI
uywCG3F199ZgGsgSh7MYxI0VBygXqBVjfN52BIXtOZPcFXqNU+cTW2PahUqUeQgTE53heMciFIlc
nfK95Qn3yplWupGnxqIH80NHlxIBAIVb0jvleD4LLvubvIGPjlynWFLePL7+bJWOn7hqvtnNUn0Z
MZSmpfTg0CkzJy6/LTUuHvj2xAnNm7oiIAWh36lT+xu5gRmSGJzR8V05Qia/yfauDgB2IjbfnLbC
yWDbIE2J5IdJQpmBaFHBq4YqDa9DGc+cRyFR0Mw+9436LE5r6WtpKAsIDdR5IXGe1QLcegXS3M+b
vakGMrqo0WMz7rfuPusksDY8WZrgtx/2akz6vVCBNoHh+8MU4QTrCENhgdxF7int2GmCfpE0ICY5
fy8F+HI7oR9uszKmrBM4anW3aO3A/DqD56ewGI40yqltj4bTXE15o7U81uk30G8gTl9kMaJEuFyC
mLU3m5oDmfNaL++J3CbBX/nopAEDd0MJ2mA5hSC7MIu0+HM1KsulPpwUdjXV5Ue7ImedA5B1Lf9o
7pu+UgVjX7r2+TzLMhL9LJiMkrsLZxHsK/p0EOW3s4fKDW8vY5p5Y7zzcYmKoD4j/XOulzzgEP+a
8/yP8gwE/WSnB1usQKXieUsbXQtrV+EISFMY+Yuz2rY+zMGxfUNa5pDwv9g1zpfY3tZqRJS0XpY4
rJmV1RNsQ8zUpKqt5BrrFbK/mWiU3LRVmmBPbhAsaVabzHlZ6QAa48xTPInjKfNMrL/rPenfZ5Di
PR2sTEQ7L9JRoAaIQA9hKBi58KgyniARn5lKrOcgLL5GeerXguR7c6iaorxbYeZAFIU3Q1dACR7/
eQYbXnHU7Q+eKYkQIJom6PfYrn8q851FkGA03Hw187nLtzU7ORu6Q/1bKWkCSPKEDuCUNKxJQIKN
0SljzamGryj1P5LD6Y4IJ55AHnSOivxTHI3JN0TVbHSXSVc2lMinOzClf0LmwXXV+dj2CCC8n8V6
CMCUGaAruNTgHznK3SSz21dp+Foj0czG5JB1cLsUJpOSu0aT5sGAMbix5y9/BgtZd+ijvwZgxjnt
V6qE88zsD2siRYWzeU82nHyaDDA3dwjj87OSiTydQbAzpMfM6Clzpy4RRLr2kd2ys83gcJxCEzDW
ZRSCPt+zFsdfuERZ0/lawE7mQWAxJ/Nxiow2QKp0Cpg31vyasbtQLamjINEvm1I7FlbkFvzYVcYi
JjMLlOggImtlI2In/8a8t4LrVwTEDoMAajpwJL24Fs6sx3sSSdBkUHRjUy/pgtFhXsOeoP4T+0gM
z2f4KLkHnErLQdErbgNB8kOyBaJdF09lAqIdMRGljtKgTdc3FTtwAtjKbqsh8pfJnOM+w8K3DIEP
NUjex1zDBfX+h71uBN5Zn4PIT+yR1JKnZPD8dVRFS0/D4AZCzUrx2D7/sVWHlaBk1LhCtYEHwl6j
FmoV3Uf3+kAwKRK5LsNdvMXWHwPj+9wxTdgtpuMAy2RZwgEX4++Buhe9ARI4+gS17oRgH1ERlZ8g
Lnxfd6mYasjcTtkqMoboLnuzQuORMKJP53JeXGu845w7CnPxeNRND5qL5UNwVXgZlHV1azVsPxFv
3PZgQn6mrw38L527ZXY59Qi78DoEM0ll12UmzCJ6nb8uJjo8UmRJEmOvPFuiulr+fjGP82Fv22xf
4+zr8eo1lGVZ7d44OBjX0gS5ewM3vW0TYe9N4+qz4i04xnV+0S3a/Cjowz3wGFM29kWk3gl5CJEQ
nOOs6fMJkdJXXIzAop0mBLPeA1YwMMlrXuJC+G2joYNA4TwHu5Q4udY9TpeRxQ2NYqZThvPAbxFC
sfvBfwSqNGjSYZR8vtj/gZ1AK8UsDV6JrKKP9hhjfBKFwMnp3Xnn8gEJFQBneYdNMAqQe9NrnAi0
9iuDu+UJLaubhss3L8oRKhEUUsC52FkeUkQrBkuybMPY5ki5SGg5TIpuilusiRcMw8sjoavRNHKy
Z++qgJldFrUpwNHU21j4FYxMZs1PDSFobBYOATyWXWX3uVCvkJdrQpMKsnMimX3voiJnauA7Lx41
aloWM8xCcqWcf1kBiPePU6VYBPc0f8fvjSxSwokIJ7XM6jHjWNKivWIeHEqvJrut02Ja1bWz8qGw
uZCoAHE0qWpahrzgku9p4kLRWtu3dQvVkH0SbtJrjCKlMtFnJ8wEX0MFI5jaOHdnh0qlbdh49/GD
9iXUxkgfHLtBCDRDk847OiMoxhrmYmdQzqtI16jChk3AM+RMi9cZT/PsLYJRblMaCjatciHKM/PL
Xp4IfYUFqep2MP8hbADPUtaXSPlgjM1wc08o6EleTwFdrcsPNlGPoHzWsrilsQeXisRo1ss7j+F1
MWyjJWl+hjHr/fJmRhVys+J1kg/1tZN4t7+L0OVkPL4s56dbfPHqY7wPFTK5GQGQmLRcNU5orAt3
/wazitlCFgZGEhgvhpwLSTT8pdT+xBxsiwpyOrJYUISL8TlFVHV5s8iVt0JRD/p47mZpFqTnJaXI
BPWG4ZqgvSzKXNLH1ihp9KEtWl2N9isAWcRMRrhJWTpXf2PIwLkSPLRHDft+JMnQ8xaSpvUWmX/s
n8VUAdCvzxMHTE0DF2sno/OHBu8EZU9kfOzF72sVwM3Hf2z2PyWlW7z6rq4Y/PToZFg9043cvZvJ
QGdAa8tZAw8VKC483vUwZFmit9WMfLNsX/5/RmtRhl+bmyxBYTGGbSPvlYBWDli0CM0CqiNmtk+z
8YQuNOKvVSSEJxmvy7CZC2XuGgsCYn5Bw77rzj2J8OHSH9cThS45/Pg5XwHTX73EMpoUqE/NWrjd
QzlZYeDmYVWXoxtR+5U05qX3PLfXFS7yizi+Zz+rDaqohQSUVLrsvH3A0VFrWRUOtHGdhoABH3sN
2Zo3VVCgdmeqMPRVTD95HApJyTkjSJHijFUsoWEsswdUy/Tf7CsYlT643NvGkTF7t/oGTdoRsB1a
1Epk5fdlfneeg5pSuIWFHkMFbM0/hUcWd5vgOFWEOjMC2H9hM8MGTyVtM4yfSgzKC6lSsAcTFBgQ
hCixBBrTrBq+uFrudK+hovGJoXKUm8/kTHWr5fIgHGdWu7TGx2bKT1PA/DY4qUEN3ba4ACoJYEla
xM6bwgyBFkQic/+Gpe6D0iTylHwbmn20xqRB9vGGDOKL9Xlg/emkaL2IIVWGAJ0BMusVZz04iuqL
35l9iFrT6Sd6Yk9dFNDblseuJmlnhqlZNFEUKvp/8IDJIj8rUEkdTJcwlowBx/azMwYwSV2/HMeV
Yw5ZRI1lMYAviLaIUJ/f6et5Vuwo68QOqqY9l357BZn4jDtML2+vzb9H0OZVO9hSu6PsiVmLBARe
0sasI3A0Y3gJXzER0jdL1u0slNfDZnctR10uEjbKWqUJ1HOFJ974dwnAtwRmkqz1MQdQZEGTlxOV
TE/2WExrHPxaVfCgvfF8R/UeVHA3tWmbE4AEfwWTIrV0u8aBbFyIqi5XRER5tKfDpr1rFrrYzjyJ
VLQyh51lweN4jk8NSlZ5CyKF0zjSn+KFF+nFYBl5SFXo/zXOvyi1ysArJqjhkkKF2HdRNdDkO+AA
sdQfvgfBZl1GticCnPH6rVYDJc5tYk3HHjV30PTjedHDMBOXt2PKglqTdmXl9MOVF+LHU3vLfFVR
8pPgEqkcAw8peZ3CSvBDM8rkXBKBCp6Y3dgEXZCSXgW/KYePuR8uZck5jYDuutWr4P98oB32kIh/
bzK5FvVPOUeQ0RC3opCjrAz0sleKeG3tt9gtxhQrk3d89Xg02NQqk1jNHFR/Zu6hXizgXBs8xqiI
Fg9EVbVon8Za29uCx+X3bCgeChgwPTsIqDsMAiQS04hpDZQDQpjDd6brcy5FTTy+qmaD78Npi1ez
yw6CQCqU8wNqQidGsoE/cR8jpO6pGTJDgGMzTMwgjnsMrMzV7HhnlCyEl5KPvLbtI2gDgNIqa3wY
Dz6RX0HQLXnNQpMVj9EKUHrsKM0YzPM5nDF6IQGHdrbzmttNkJm45HzuJZrEw+MWq/Pquhv9tVAv
dM27hj9ACksf9YZeGiwfpGHnnt6NRFAW2rT0+rujb631PbnfDojboxZ8/E/Po/IoF1bvgnEHz2/J
qIHwpxt3GmpdqEwCyfFzFxWBvYMVcKUk+b/r9yxuDrllAwQS64IofBrWhQxwNS3rmM1/rKlfiF6a
sZMhiuDD7lsWfOnapdvzmhbixD94+cclHL1HoJuQ8UQqQ/9hfVCakCw3TBG2ELEAL6HnPO+ZvZOE
G2a2jxuK/sPLF4G68E6xHofsuWTdTmegGde/HkMPfczCfhMYJvkAuwiyXaNsJjD8Ww7nrK/csSfE
S0BCpk3Ek3OMOV3JfemrJ2Ba/6s3kWXn65Qpqm3kVQf4Hxbj9xmAfPYmyU+xLsRkdEMwW2glhygq
YUtetZo0Eaa33/GND3QyKx2WYnyeS1HA68tHejgnl2J+yxKPSrF7H7ABnOopT+oUZdj+N9xmtg5G
bATpo9hnVOv++ZpRA2+K9MGnl6B1fHlHgHEskHnWftxXfYWaAUG7TWBm/2M+Tx+bQmwVkybcYZZf
/F0zRuFX4WqXONg99uWXoaJIbvwYvpXtHPxHB/W03lburqukNIbZVoXRjU2Rg7xcFQQ8jZwOpakE
ruYWftjDoUpilTOga+udQxN1rUXyzbxZwGdjYsWrQwAxxCFjgXZ6uE1oK5ZYoYOvbRUL6dHQ64/e
s8T6AGc9KCnOrvRROkbhBMVrEnkyu7xx06ulXklsPJvf14Vn5lGI1ZR/I5QWELSYGnOfJAAMXW6r
muME4MvlYj1NMs4eCoNUCQ5yN56FupU8X3aUuwTiH4GLC6znsRm1kA+2pcPJ5/6XQnrtSqB2oJOV
OwzpykyisFHBzjh2qkNGg3S9h7/ZOrTZv5bMTdKtVreLvtqlL8Hzr1GzkimIGBcUbp0pxruIHSOL
2T8NfxGFpcMWp3HdMb+rsBUUKUuqUZkrUTQygfggh3Di5cX47TV8pWgS/yIQu4PD2mTuZw8MQ2dp
u7FjSIPeAa0S+xKwaERX6iGQ1no7Yr+IE1cLg/YPYrlN06h7lCQ0XUmrk817oRXeKJwPIRuJzUEH
w29UcCZPIY9BgUiCyEG7H57qcHtHGmFMOrTtsGaOuDrZrfudrC6csuJQ48/B3pjFVecYEZR8t0h3
72MLp+hC+hUJXnXN+bW5ZHN5gf83uqK/BCkp18KGKPSysvS90sCK6A9LCi5nq9jATxfaYRqeYXm6
LQOWtLWfftBeOvRak9ZUldFErdezmtKoYbnDO0rL3lHYf1DmF2afNoUfHxm2nsz3xc0g1sZq4qNr
sg0vGoYC9xI1jmltt2OEfybZX5DfK3WTvcRyvZ/dGzWGHy8rlZvrgKbgAxg4mE7VrNhtaG6bSk1e
n8zaF2jIwCmnZ2H0+7jNc8sT5c0Kk4f78AqiGmGAaGdqiRalyuQjT44BxQ6w0feK6f3dWyuDp4s0
NDVgYqnwIYWeLZrWB/PnPFuyDDu/A6NtSwl0BBqgml3bFHT27N3dehcBiUD6RyZtxJZjeE1MCKuS
GRhU8fTUJbHcqBP0xsA7qRWLWb1WnvBkbSCHMSuDPS5wRMLZ3SKJ5D6o3Vgd/oxlgWMZgU85XsuI
Tv9EnKe5unFhk5NcWBB3X1djLDTqmmq1bUCCDiIlRGYkp/oA0x2uX2HZFSA2LqzGm/3v+y2rIOMC
vkF/T26cbEoiSqa/Z8U3NbAmxbgo9bVhxPIQvEr+Jb7/Q0wi3kPP12QnKZPDKwZp6rEi0gbogvS9
dkJPcLq5MPDXURn5zFx0NK23Rs55OSai05riKzcdcKddB2aMIevWhJ/R2ACU681uW6oRNxRXvLFz
u0vr+U3Rg1nk9cwTviuYXvcEKUxdTwF8S1JHWN7BJFnNVdWXnTSqs/rb4T+tBL4uSCaq8l+xPjXu
5OHiqoh5ZkOglVIeMCx6Icx+FLFrSaspr7YO8aOXKL3oZpwnc3+RzqDTTyEvgEhntuELjVm1XnHa
yU3j54/2eTvkjBmkmLPlMI6/XcW8vgDztS2fCs60z8m4d+lS03HBtOu/yB0tsWvTQzL643XIcW8L
mh/Aknbd1n02umwG9OSje/KH20lKhk3wjFLZUsrbpKXOWScFw40mTvgkVrpBj6Viv9LAa71NUYrm
UenObQIjkcjHZwCY1QnjIbHMTrIKVp2Znov79BfhF5RRDr//n361wVQITLYUNFWFNAAKFeAvGJfe
/unrwrgtT7pxE76EP9hqhKjgN38eeNH9rQVqtOMem2GyUshMmeAu3rYOiwkjpFFHXFksD8Yys1KA
oFdn5MPza0dJCtZQA3QMbfWbhT7kvI3fymj+xsQ1Qf8OL0JwVbSnfHYxhW8bjA8bGDObsVaxQlIu
ZgGJs1zJZ9ljK6vbkeFAkTYLnWkL9CxhybJeWJ7i7JFp3KWZT6JVC57PfsVRHo3EhjeOxQUIV9qt
BqQtEPURxvXX0VMxOGDuy95yidSxhECBSwd5YPUo7wzCq94BN1n5mTvxgapHOwMuBLmdNKjT66of
nkjQ79oFLks4iOfHicD6SoQmF9dhxqolPKEDm2cbDjTDev3KZPwKPoOSH2Y31Wp2YwuLh7NjKuWG
KrpjjgvlF/AGrPJJyCZM8Ub8PD//0XsLqLkibw8djgWmzgzJ+6+F/DV3wkFyJrUYCuQheUtLU2rr
N/0BeJSe/oa1txcnswBBm7+8CiLnEnn1alm969uGw69MO/9fcY6sWdWKZzkEav8hLwCBpS6JXS5W
YGsbot+k7sYifnTtivkXOrwrVEMoeU4XyGdYPf+N8ZwfwNPB2RhcpZQcwDbF2v+eQts//TWexVtI
gdu5C29ieeA1YvpedMOXb2p8CGKnPia6tavOZiAvA+Y/vSuChxFhX/bFEZbPZcGg5Ku/lTPvkM3c
mwD3oq6sk5HMlrdAmQckhslZUtL+QDfVyuJVxzIWdLJjiu3fflLdDkZv+ZkHP0RIouRxisPcLFDU
wCKKWLeAKCCLpoy7D3DYel7OQrlpT+TTSPdRMI+bX3yM/vmLiEKvbEXk+SQQJqVY+ODyWaDB/sYq
Jzi6Zf3RlzNLpSsyRhj9ucgo9C1VflY9Oh2icOHLoowl3fljxp+leTkc2JQParYgFPr17FWtSyRy
3xFfLDIWogtwQyyFR/mME36LH/AQ+9iV4UGEgSnUtTuwZIDk07lmFFXJEnsVDOy1AapDuWJTg8Ag
rx13VOvyxHQ7GFt1N2PiTQ5FFjSqq7f5g6XthSJlxOlXFzjROH1F8yhMJg4KGt8HENJl4Wz29rsW
W8XaHH3aBTTSF6tPNSKbzdJ/AY1zP2R9BVXNS8Hlx/aoOmzAuidvhluSpg39VgdT9H9txp+6y674
lJkPSu1Aks5LfNrVsfGZqa2Wf5URzPV3+Vpvs5P5wOr4gkDPy/O/39Sdl1ruH8d2E7NV2iaxQvii
BLZ9G4NsWteBYyFjWEaOqXPqkgVH2vZvlLuSwFNqA5rLsKye2nKEnGBITjPtvw6cEM/2sbdHnAsA
Or5CBRDpfmvDNjLtY0Kl3W+i0BT6DXdauc5J4m6JPJkvCwI5R7wbtqmVqlsKEwISHmhFweU7Y8Lp
Lo2ok9x3Dwuqtz/3AVH9+P/NXo6NpMo2Y+3dipaYF9SWIKd6MVP4d9c/cquf+626fc1LP+vz0foM
d1maSXTz3HA5r/k/I+4Q2oXppslmCDACWNe/5VKABXMLjRArqSOGCHH68+LRBZtfiS0BI0XPUH0U
cagBK7thqyj5n9uPq27FMz0LIoCp7ZNo89EBhvfAiZ0tIv65lAsrXWxuCpUp0F+/qeYV3c9Ittpq
K18WGa9E8SsjToVsWQDRERmq62Ezc8Q6tnqhvn09I8k3pphAAoldwn2Wk+GQZQnlskCPODim9168
4MIQ0Obo2SJ3wQLKPIe+Xg1Tp6+Y1XdF8Lgne6FhCLCZU9BQLjfgDOJSJiwsTD85S6b5w4Ji+Om+
EOXXYd5iTFJpt0HDVH5n3g0mdQfu/IHUMlkOgF1jVCHREYGDipo+ENHURs45A9subFhIRm4vwDko
VZMVtH0JFQOl8pyfWb13cx8dN1XUovCAbRXvPyesLmo2DPA/d4soeGIn/WlxAJs5lLzazGGh8Ex5
YXYMqoGa9TKHrbbN7igiO24b4XwG8aCy9wfcXvvLItDPno+AtvKvWJWtp8299w3RR0MYXqWiBd74
cG6hL1HH3F9uN3H0xPEJfV2MC5Ej2m4YuA/Y6wrhm7J3RI39HmoarWgg07uXquUy4XRGKuglVlo4
L0Wek1+jTKk3y+r5NtMskjzmoLVqE5np78MFIiFv1JHNCCKegb9bjE1f01BwDVFYF9V4sK4GQ7XZ
3S2Ddhp1a6VXexNNTWSXKyJb0hADGW4TlUz26z+ogmFr2YRvo0ueCixUhX4gnaLsNTN32pkGdHaC
cBXpl3HJelXZKEhiBOuJVKI9W7plZBIlRmomNyn+AvoS7vDSTr5PcKrUmguAsX77W9kxYoR5cJtL
7Ldo04lz0mc27aoyluGkzd4ifrE6Uu4qNhZ8Z449xKepdvKtGPVWKhw6RBgI7CpzJdMI23hx6SZ8
qbSkfFXZ2M6CyJLU4wTkNf0h7CaJOfFF8ggtWfQnGg8hk74jJLh1HkJel2UvTFgucMlTPKk9bEzG
Cfc0Eh3o4RwaJtueo9FjTFfEiMIhcST9X/oaw7eHE0W8F+/d85u+TaS/qhbe6NMNK+iXo/fNoZSf
C0fqSLBglklmDh5kq9gDuk9cPgPydeZXW8ZnOyam6sxG17QYNpqNtIWW7Bmx8VgsXfMprJwT1Nt7
++dWaHjJCArpoMgD4LSK8Hrb/unHBIg5KLYPHf9Yu7FfHlap6MMQYHbsh22tRSh48J3jbGG0S8ua
zCJBaT2UCyZUR526E6chzBsr2j1wOZ/V+vC2tYJB+izUyn9f3nsVz7bz4u6EdMKxZpwiD0C9kVnF
A19aWqGgr58PfpLR/Qe1P8eiQ2oMdx0ibqyqpRK6Q7i16tD/3/9+NMKGw/Pr15TL5H2lLe1IPytU
VOuVNYNyOt1k/oYNkts+M0aeg4OYp+qaK+KPFqiQCDNX/WI76Xzef/D0KPxrAiP9kzZrftpxypKM
y8yEsrGs8RH7k3B0/qQQr4n0NU2u2j4NxCkSV/wYepVvGLxFnMoffkNnxOWM/R3uFl7cnNa//7Ds
iNQc2jI2DDIcOh9rFqH2GaxJQ5nvYmEGxwcgEDJdWn258f2mvzp3vxr4kQBe9ideuC8jUddAcKOz
XyCAuxKTTzwtb18BGyJN2EJd0R1peLwGnmfOYszazgJGcBRKLeJ3gkgqBxemTZv5eo6E7Ft7MQPG
p2i8WKVwlAJSwGBeFOS38Al6qzAt7OO+d/9123bvBEYCdqhqsrnj7PLh+mtxsTs8giWxP+KAtG/+
dqxSE7iDkFJYTHN14VCnSRIWhmOtdJCMFWU0B+cGUV5lxmGHZU6NKd8Njqc/McoFDwrA561L7l9r
1m/7GUE99NEkBumimPwHVugySUf7YUvS9i0JxDiKPHZuoxDkVd179J39rgjB20JsKXCxX2UPqetE
6ZExYV+Xdjp/dtwfuVot0N2u1z5/D1sAwX6V0Ef5ZQ2LZ8fPYGqhqQOu4j42lwv7XTm83sfsiM8s
IZ0SV/uVVErznnEsPbu5GgAyvnO1pU2jHmfJh1TtuqKLWwqdJ3kavxo8W07ybvBRq0JCYEPJ6duN
DjwU6InoWL9LLkoGzGw1F47FP3qoOQnQFCXeoQoeK2fuJpPvu3uKeM3joQDOFcmc7KqStREnTYB8
zmYTLFxnCm0gYvh0aujLuFFAKxIWIL/sSZKkQ3JMSNEkUsE46z3JPJ7nyqJDOTIfQiGxCEEhPk7N
jPhVG2FdxpM7utzulMDpLO42/oqN1dfawV3Vd2uJS3zw6eLUmoD5F02GZuq1S94DJu57oKJl2R3K
JyUUveE6t/qeCz5blkpIvil76Zgaz/T3Wsrkx0z3GMngJWT3gC7JdC07A7Ds3THVZdjil9t6nqcw
xZ3U3XiY7ZSV+b9VyuEdLR4VRzBBqPLBKdd8a+/+Y4ZXDEEoeuGCK28A5Ux7S6SenMw9b1t5NNtl
uf/9CMLc+KNpS9eC+S/daIlwKOq1jCa99lm0mLXL2AgJSKerEG2Ii9wIlnvV0t5na5gw8if219DP
40bdUnj+udVFLuSp9pt/2a0rxkxbuCwRc9N2TEpM4Lryo+1EW75knWdbtWbpHqfv4+p72KW8eagb
z0RraG73OYxc1zv4HL+04IOtYjAZkKRUb9cXCnWLrkSZ1mB2du63cle4faBDNoqmQFZZQYCiRpe2
9E3lnMeTr2CGfofNwrHBK56K2odRrbSz4wSIRyxYxzYywJ3M9jDYdfgPA4M/3v6DpK6+AO0Tljl3
HmFHmgAhPTYiSulwutWcd9Jg4fasSCde2TTFPFo2jssqj2CUkdWrJsCVzIFo6FBbrSjAHB0UpcfO
1tyMO14lLPHHDwkxZiKafO/iFbbBCU7B/EO+vsZmxLpnX6H6HJ5q33gRT/Lo/FSIR0nNdObQatG+
aE8irQuU4kwO3kiGf4MomTU9LjN4zWvq3TVnJH3ho2JkQbTV0+uY9TGobCu3fu4K61+6/GMLYdCl
049DMCKRv0xH5eGK2lYdNhOe5MROdfBR8RY331W8v2pBlpqHRVZC2jVRjV11ocHMmjVk6N/tCzAq
gri0LQuQmtt4cziqwZCibjmjWhGp6CqelWBSc5DvaMt5ppVSh8ERa81T+lOuuKzbFfV29DsaMAH/
JqAJN3d2RdT62ruvf5TpZ+e336fmQbD49rBLWkEq1jfiJC6kAsSTd1DEnNhjkRbtSfSaDYdvpVgq
FD3ZdHNzJq6VfsM1z8RgU4CXjgaF5ktTI4FhsItDyUQQKzwt/RWkuYYNmYWrxxziHHLVt+VoGzqI
TZ+uswK2f4ruz2SzOH6DDtiRPyoLIuZQlRF3U4D3CWuSX0n7xp/MNXt8Sw/HtbZEXcS1JikIf7fn
3/uezETijvsjHArcYKDGWtjaYR4gzCFzpDo+/oRvQX/LJI2MPm0/u1zU1CrHFDHkNX7O0vz3f7xc
73mqqjukb9LJDl9ZH34xpvTW+CasZXH7ikZjzxrfqA9BIYKet61JH+KSZKVsoSjHPjOGBdAGy3lo
7MglQI+TjQA58zjPfoOTUk5LSI88+QmBSH6qKa7zoyWJNYXTLH1kbA0A2SqfITUHwx7GqDZf2h30
hrw0GzG3vYrBqt/R801rFgKk1kpdobXGaclvgunBJFr6XtUI9ddoxwcgjfo27CQyirI49Cf5nKQf
/d1H+zilQfZRrZdAM4hlgOqGxS/kzYwdfI8hZwotJQhlArAXBXl2KnQAB13sFnmqAars+FE7y+Q/
iIVzsFWPlKeGwZ85S6qaPxZ6EpzCtefEXLy8yf4C7Imud+zDyiPD4KkzRloead8Fw9UkXb0ArmEB
AU1I+aSyWgUE8tOAQ2v4kdn8ycHGY48U4PXxD/Am9EeDmEK4omMCWANccbrHKcewnBFojwSG9XFN
z3/P7ZUR8L+48ZwYgJ5lLFlwZoVejHZYosMH7e/vhH/M+a1kpwWSJm32Pb5iC4LwQavtKX1SFCjg
rdLk0ZobVPSOHwoPioyE9i0RpUQ+VsfJKgtU5ATZ199sHnoWchpmVIPE2rkWWjMC0lVkmGo6hblV
js/pruT+zzpSpBqdxKJG5htKsW6X1FNQXtCiXgPy2A3r8afkv0z0MU9ZUA3eBJM+qYDcSX5RLvg3
ByaCUGZDzPlnDswV++l1XWUaGAZdV+epyPx7jJXEJH4/DjBRXKBuTAcp3ILrEOYcLveAnYG+XYbn
nH8NR6BJbqWsaroPEtfYaWcu9m55dsqSevZWO3pt8G7igTJ3NlhEcyaWlF20nyZwtrfK8vKVBjs/
c3/C+MQNglTGo8BUJXKRZgHc4P5T3grbH7EJpA8nBnGGXvXxYLEwjxM//RehSxKsaDCEepw9h7Vf
dfhFPTOwzoqQBKf0w1HrFUpV6REjGJMDIJIGE7S82RL7LxzOFrqNfzKpA6jxTVJgx3Lvm38PcOPm
WoHaQQuZ4nf//fk4DVcxjheljiSDp47QRgLVBxlepC7JQXx5Hk+hhsF9GO7EMBTLQ19VyLYbV2Cp
zOHvJ11sAhqEnqsiKjpn6ui8ewIcyUVNDQUrDdQk6nnbuwM49ZN+f4iLCyl/EWoDwI6cvn4An9yf
P3CBwBTKo6+bPedBMlN6NM2xzXB7Rr/UzNqwmo4Qds+VrS33rsy5H8A/lNE/t1xY1gqBEbHSiFD0
yw9HFAXYGv2QZnzeh6NPqbc0t7wZ14OTEVcwfu0RP5SE351yxkSTL2P32izpE+nLmLOAWNMYOWaN
LdG2B5Y/tZ1kvzhFSrF78IAsIYT2u2V9CyK6xpL5kVpjIY+SWOgKMGaw4VclRlKv/12l8+0vCctS
pi4CfWdmsCHn7CtkKUvzB4gy2GCLlxTm8PSSCR+AG3bDzTH9bokME6zJBN8klX9gOHdySUZsR3iP
O75Trn9BpL1k6mh2CJDqPhz5J+C99CsYj0RuSMujSqmWqnTsW/O44epHiThcjj3hYI20a1+fKxqr
EFKN70d0m5Rz/s+qJx4YiiynVx2LuP7st2KR0xx5Qlf9vRA9bLx8LVxCc6JRHvopHx3UGtsjAkel
8A7/z9Cj2A6pghKp1yGUAGlUQlfyAuyVW/6OapStT/EO6tjYfFBuQTwDPDETWE3ixxTPBtm/fIL2
mgDGQPq+kNNhD/DtbSxHoEEwf8j+a+pobbC1V/JroORf8mO1k1IkhYLPeMLY2YjfaM4M2PW557WE
3cRWqa9X1gsnpvIPdR/WBuDG2HY5jnjH5vSbQjGpW8U3hJ6B++g4FS8wi77RoxEeeBXaJMVL8tH5
0CXhw5XS49DI+hF9Wj13qYxcCNojPstiQYAcl7EB0flFh4gNbN1e47IwfPFRJRTLoCVxnQejopUY
1kqksvL3TnAFyhHstz1cNbko1OPtrNIet0Fkkp05q89hxPbqDaJA1ekqhTsHWkiK0GgQYkYLLpkz
5mmPYeImg6TTx10fWae6RLLEQIdwtuEtL7BRDLr7x44q20bwPPBTOJ9KH9fWSqbcdZNExAcj3fhJ
6ObmyB1phe3tQImEElgpvhrCBz8uzJbAQC+u3KhXwVA8HbZOyBZNQEvD3HBhNPPpEgqXObTgE/b1
UfTrudqyAfjUZU3z+MdlRid6so5PYEHgXu/SwPKNhTRH8S4XkrSzw8BcNoJIVLeieybKYPf+KlDp
1sEK2OH5lBJtgDhvaAWy149f3FanZgQYbK/dgsjym/MsM25o1ZwOFh1h036g+RxFZqlzxMOt1geN
NybAz3ipFpzn2sGz51ylWqSljtAkvrFzhdshx5jRDtplkUVn/QdDZH71909JKqoMMFniCBANihPO
no7IPlbZgcWijPFkjU1G2tZzSYqfiyCTPMVG1Qrw8iRu83930+lyk7QYP/51AqIiAeLvV2PCg4Ss
0lYsr1yy8AzUa4K5XLNFL+RmLQ2mGQHDXBGT5bnhax1GuQjyTl8FUQdGNhzgLHUilHr/yGb6F1gV
Vtak4KCVS2ihiMaTb0epOz8BEqoRqEttWAiCaydKleXi2l6TuSxfydCNn38GmG4Itu8BE1SuVopz
efNsPraMe2hu4k0IgBiRMUhrIiLZS5D4qbwOiLiMkrqNjndzjGMLp+GRFqaRUPdijb6UeV7z0KES
TMrrwCFv0jKNRteg3ASUNTP2y8mrv3avjBuKsCgnKWmd4IO29xD2heklSE9cKJL2N3PaIE09eY0+
prYUzaY0iNNWrmJHfpxKcT54fIRPRwaQPNV6TTlslMYtRWiWDYVoZ720TQcPPnA2n5ipV+hxABnJ
aUI6yIPh7qUSr/UfCurdaehe0gN5mTJOYxCLLJ5JoKl4355BxHLF7l6Ya6SldpaZi12Orp+lrtfh
Z6fSSecL6bB0OLhgRXE/DXBvcah5cG5y1XaIYMWra82eiPrcIkKeaby4XpRX7EbjQD37vo3dpse0
Gsn7CLqKosOPBGV8J82VytZDqbSsHqkmoXrDEbID1JatAYcNPHXPGyL+DgVgFDrv9Sp0hzO1VIqm
NhQkZAgM2XI3aDoNZRNB8ZoV0NhzioNncnhnPyAPFFW9Mv4B4mPDbs6d1mlAx78mTRvJhQriZsWY
DI07kl1ZvaoMugGtTRTATk7oXaE7TiuawKTDzjNAs6TOy1NA/4buIkuN9K9aFlbHYs0t10spesro
jnppXLLXqIqT3kzRg/uifUnpWE2tfyhmCV2aPGbzfAw9uPR3lw1sCUlFhkFELJ9Xg/KX/xmxS/Pc
NyMMjdX1KjlvZCMTqfjYVpZyym6UoN8wgWhfXqGY28p3NDtYuCzO/9YMe8ovHzeDyaa2PQqnJOf1
Zb5ylga5q2jDAuZDn2X4X9FAnKBaW1E7ljhSI83dNSoQByRrOMFXrr83RdhoRrAbrl1bp0ncNYVO
79YySEj/30ZZVGqG+gEfvMq6soBvLTZLnfaZdSwDbw+H0215P8T+OlYEAkgHmEVYVVNrApHijjNf
6FYDDhehTrKJGchLuHiAkDLou9FDo8KJ6hYNACjtfa/tQ9FPoFwT78a4x49MtljpTLUfV15XfvM0
su9ZHunajl5zN5XKwdhA8L9Aze/PJe3FfXgsr8kBJjIuvt/OQQh0XQh2izemT7MlvCYNQKYYskEX
cyqwcbnVwz9V/g8XbGhtGVMCdgjMD0gqqrBjD7IAc2qr9V/uKXzzpiW7jz5185DjIKhMVJFNcCnh
QMzLoMs4sPtECMg+EVVITmlsEak5TliGG1xjyhhZOCy27kT2GYIUxfajzeXHTrsRWsZpScxdTZoV
cSaRGFgJS6mtcd9iXRk3I4QSx1FzwzE971LYU+v6VQxDhXYG42aEuXIlqSwoZ0MivZ05kMH66FO7
Iyn8mkksTYtMbpcZ+Ia6J45XME0vTYzjqqEZcr8baI3wmQuph5JLor5SlvH+fd+FUIzrRxejD3pG
tghh1IeyiL0KCwHcQhUpW/i6ifH5VVQ21/YQjrH6PuuPHwNO3ie7/Zgcq5ZL82aCyEAeDPM+EmWC
nCwSXST8PDS+3gM+i6PlFZ91kNxDDCFPIxAKShQn+UrLBVhyc/mslszMtYTLAXcRctJDDuhIyiQ0
mIMNXc5bn2fWDK9843HQocezHJfPjwkiPhybLb5OWPA/yF6wKD7cjlk6fluYNibBz9sb96OP/EgH
whji/qzVlxD0r2Itk879e+ahUEHWRcUdVifRZylkD1zC2DUzzRXRl9Fdp91bF9cYeme2ujfmboOQ
QS+j/yG+9q6VtcDYnPUygM8gqULMAazs7Q6CMMhPgfKeBqmGCCXMKupHPmLgBrTyUEJqwYhWYK4k
xrunrK+VZTqXlQQOIr2TO9LydBJYr/mV5luitaRYcP0SiGiDx1g3BYIc/UUqyTpd+DUhtK4tD6xY
EWgupNLgbyL4E3ethGX8nygRQFgYobzSafWqJEgSVad7u8e8WN+rHnN+JiMjZ2rY85prXeIe5eq5
ntDeEwFG/Mm/PnFcq00N8mmbn8QJwJMYU/2SQqyxQOYDKGneKv+JyDoj6V0t089fFDs11AMOjovt
nFHHXtImW9pIYqGa9QuMoO561PJWtZqSBpgGO8cWUoOL0ZlzgWmvDJPv75gJZE4my8UBdKD58OWu
j1ynaYugA41y55Ikh8xzfJlyK+gdsikMR9e4wLixAShFKnowAuyTHxwX1p4tQaO8gTu1af8XVIvp
ld7Sk921Q1qIKHge47RlhL29nwdUu81MvY3mUjB7xVsbTLv07qkBsSkmoqifgeCnzzEE45dCWmIg
OX9YYLFkDfi22zwtwbEKoiU7pBlLcaiKd6VMYHbRgB48KMH00WDeTMBJ3DgLFRAMgP1heRHWjVTu
PeJ781dy4ufy8tWWhPLBOADoFYhZXP6p0g8fxm/ORfQjLXwllzfnUBR/lUHuefd7kAYbbYCYsuQq
TJ/UCDaV8xFiFTLWVv/uWlkj1b6HxU95RZEsYB/6hBvWJeMo+HbHlFAczz2ua7KPx0vugGKlhe5a
ypXycZSAwRglwlPSmAeajSaY1HFw2MxcTpMAG6zdEc3ub1z/IZ8z6f049ViOcByEb5eTsQMwJt1Q
3sOI/jApalYkL6tXQYgTkOEUL2VE48UdibbZBT7SjZzCWL/7crRGtaqcJwsLwmi0Dv0HU8H47Zyx
xfzMeyRBCbV+J536A97Y24WfFDA30v0wjspIvdFFWHxqdxnPoesmkAgitcgsIpfsgdgKZPeBQ2Mz
UZreIN9G5MbzbShaz815s9V71IGinY6p3tFCelEQA7ZiiGAaNoB2g3lWcdxQIYfxOaKzT9Txw88S
1Jv+LBccn5dFnppgAQI8clE+YaO5LfmNarDlXdP+cYbufERTsgQGumKd9JMLXEHMql5qiZYXU0mm
EiDYVTP1rjnZl0sbx+OWSX3FGrWaPmlff1WxLS78fXJm+3TUSAd6jWRxQdjlQXHh9NQvhGS2iMdi
Dgl6lwJ0BicxLWKmefM2423W9KuBL5ZkUbNqliYn09mjz5Rrrb1FuO8/ohU8PaY7sAeSM9mcBQuQ
j8KfGaYdnMdNqz490XPrp4CKvuqL4wLV35o3QESiXVkIDqLW7wPHDeDwcFHAtazMzillW74kiCr2
q9RlgoO9ZZ35EeqP+cBLLJfRoMacKyeAqtPwaTFvtwiAxO0slv+WLdGHdJvFvS9v6CUzZREppogR
rDVvTYFJPs2yzcA9s7c5KqFZ1loypE6W8NeKyEwSOOc2r0jIONEQM7Car7LLF9mUSJttFlALPM0g
TvIcrtj6h9gqhvmmFF4fI0wcKgd3kZjL15dQAb88VZbLdtj+QTVtLnb+VO/Q4zO4FD/wLQvR3hB9
VocPmSbXky3K80iOwad/xdkDpf4gzpBoj6y0odGjtGUZM0LtXy798ndHvFRimE/qaRV1dNpCcfKC
/OXOTR94um1fPqAn8SCwp1AaofCinaXBPM+JRuXn4tE5CFqNPrQ0pBQJMfdSuRDNfur80NrlJIZ8
p0h4H6EHT7JDnNVyLtw+H7JDxsBVJtdxo0xpAI+sJG/7PNa07FHB7bA8dWh1kmgFNu+ljWGN5uyw
7Pw9dVh7Oktmq9e6B7KM3FoV8qmMUyIfcRuRuzUoHRZyUFUFnzhImg4dLzT1I8yCuG8jeW7IS7/5
mkYMK3m0TiXBlmTtqNPlegZJNSYfLolc6ziW+NoiP5kkByLJL32yZt2QO1TaJGWcvwBEFuilq2la
A94cwLBshKNJJ1rV8mFjo+YpMbq0SutJxlt6WsHRkm1Ajf0EPKqqNXK5KC1w0CSgXPbFExRiQ0tF
SW8kdjHFeEjFqKefUVSu7uDDi9REQ17lFrNrTL/swK2SUidZ04XB6qmGicfjqDBe1yo70toPksv9
xU1BpaXxVhhty9Wbrq3TwzgGRl4W2j0H/8ScTcrNDLFt+/SoNOTWnSHDLgL/gUIiCsTeXTPid5iH
PjskkuTLAqgAM50xnW83DE7Z/CfXxu2zus6AXCLQUkgqGnVWbx2Te5IZ/xZ3bx+V+c50V4sJPSHb
tDRxCyIngJbOmi0EHM20THAlCgYg0Mo1kCBOVMyXM+zsw8TLz4b8NmyPXevjSR5chnKnnjBtFFDl
bGYO+zjET35cVVyyhUrwjuIHXugFWdOqaQMmM2r77hw1fP/IWHACZHe9Uf+HSwWEkDvkFZzMY/+S
48LdG+veezg1CuytyFX3iKAYnU1TMAdvbn+E+tbP7u9mX0P7kg7nLF7lMU+eAfox4hv46I35ezZC
5M9A5pbE1zVPZQKpCps40YScs1P8tDVN66au/V/VaGM5IG0NrbnTQ1NieqTiT2tQNF4DlJjQFwu1
7yJKngfAItzZyLkbnEtq80PXIln9VmMj7gJ5YPRgbbHWRYRXStgS3EkpXSAEqeFFQ/ABxhhEkQfh
TTH0Run4K6RYep6Z0vMHwqClUSGnfOfebyj0nbS109Vqdw1lKTBghyZ69zKHzRwWi0F1AFpJxX5C
qeX/ZI92slGgBZid01pZWJ9SGxYQ2UcETA0YlP/X/uchzaZcZIDhZOM82fORTdaE1ZMqF0eTTwtQ
HFMv5rSG/gV7u/hJxzwrXnI7xoK/M63aENI+GsExTfFpdxdp7TPXwG+lPC4rDquCHDLNZpeaGUM5
TGgrWhDAV/svduOOG36XsTuT2vYxAEpLUElSpMOfm1DRTHGHFEVbm1eI5HcNTgg5iaz8tnLFJfdh
36Vfej56+WDMSq7VmPf1vxiy4dQKMeMt5cVbvupb2HfG791zoUQxC6f3XPTMs3OHPgsW2uXnoZ/D
7C4pR/JLpm9yLEbcIskJtM97bsIzp/SdNzQWhCKQsHahVqz5grjfi/FNFsiXkatBRdzFnrWNTnfU
KACOdJHSv0nIu0funpxpLe4hu903UtxQqXeOUkiV/nGRq57SlFfr274x7XHXg0hu46iUsOaYDvXd
UPa3gy0lRsezP8k455uhF0gFQI/GSLmDgKB6QuAJ/1QkQE6kl3EnhRNr//rTkNzy02MTG/3EN2Mf
EI0XI5ABHpGzc3RkZb9YN1u3i4OmZKzuoftBTsTZvhu2n33qpJ5X0a1n4GDXYmg2emAXHkhAQWbK
Pz8bL9ZVqcCUqsgurPQHLn8G6aF+2I/whZwTJwT4cKjECsoCg8MdcTBZ/x0+PjaTEnv6uA168vlM
1J5/uxsyzF8hA7HEXFsHpY6s+LbgE3glm3FK/ECB2UdmGLTplKd8+Ll+g7cz7Su4Ftq65x0z5I7k
Qy83eZfu7UutV7/CDVM4NMO5Pafwbs6f6fCUoMuIjm3L10EP8ymAV8y7FebAVxUoYCwVQZy2ve5i
St21EVLwRyktD1Kf6mcy8233p9G+JoM9/xb6Aweb7LvCfIpYZ0GlcugMBeEK7DAUo9suTpPww585
G3PB7uxGuajM/ohufy6xqHcSU/jwjWPBQezvxBKaF7QDJ75gh+4U059LexC/OPTL4F2TSnyHt27X
Xlv79cSo//N15x37mBqu7/qPHj5m0xZCDh+rnlL1qTo7WJH+3oeSRDwLZaltQ+3OEYDPu+bW4Awe
Yqxi0QrN5t1dD3Y5OmnadYDx/MVp42oG+ekESVpvSrcMMHJRKvOtkFhGJM0jQQLByF1pJHRjg/c/
9hU1UqTe6Y838CxcqucrCimphSJtIzEIZBeIHLyJsxC7TFEN+WCE1PlwmLaSNHYKVA15DcN4aX7B
PCjKU8bHghhVDQZjN0ITp89WrVO9PPcNmHf8WHL+GcNEQyX63gPQWZgXYADB4JePVRTtxTetylCT
Vq0LkN7/qtgWdpoRpMta3MVqmfb4HHiKf4ejE+9ZQZkpZpR2a0dytTgaQeB1isbxrBUy2xCq5q5b
OUJN3zWb3pJWKXanCaevGGFQXAt2Bj4b8CQVPFShOHVNieH/cGY0p+smYLOUBfcPXeF/vP7wYrbA
vYlOYF8+bDdBZbBlBMfKblNecRjYbjEZaYdkjLE7AouLyAEe60hpHrhJGkaZEqsQ6ChaJBjngrNM
+2pGCzG4mjLOyepaX322i02KVuH0AIafRkNaCvnb2qxLZ8cWrAo7kRFxP0oiWRg8bwizc9uq4htv
5/NP4k8J0abGoiapaBSzmQO964+ZnZwD048CJLuhCSWUDvmGo7ICkPQ8SbCyigCeEzjAlZX6mITY
uT8treX8zv1uwMyCNorQOyQZ/TLVAX7mUUO1DxJW8t1M0lXgJ2VJKlbuZwqIgm9K5s1UTJkfyJNz
qKUAT2PZ91VqRQAgFLXgxqxLzcUvMo9O8VFxkhJpUNuebDbX7N0T7pm6C4JwmBNCyVfzrcWjwON1
8U1jvuL0WCvxtdfWJYbJe6xPecdG1XntYNydQb7GGdTaaYup/sknUnfuu3HHVho1OsNCn/6ll7Lq
iLLoMxNGpFk66Oaj2kLZcjfHXeyl6g11LSR5vaygHhxqHSReGaN50TY9Odzl0nFhL0+C3/dAltWv
/9HKX183z0x0CoeJl1yTivdLHXNkZUxGiUFnSrZVYKC/KpyuadZF/XSh3vay/QdN8RvVYz528/Js
Vb9GjQlHxNWzSIhYRk8jvSeco7nvdgD3d2qUah1Bxa7CLRbxaP5VBY+LokNudDG2kjq74hHEgmVN
nVl5ewg3Q5fnaqI8rpyI6ofrVkminZDgH6+0x6BoO8WRb8Dkz9exDnHCshg9BGI6SuUMjZoOnBeD
gJsPIM2E9z2RB3ZA5JnEHruiNqJQoBHY4mZXfOwReRcLPzdoI/Hm838QqYxOnpNB4AIIq4Pj1FRB
/uVF3qIToFTgm5EZ4mcIxgrnuRBwVUwufb0gavaDq9WrikPnL2+TMbWdZAq9a01tYkwCJXqUNfGJ
UppQkrRarhOXeQ28s4XpIyocGhR9E1mCDSHaIsfym4AOvdDyLLjK9mpF/l7qwNlP+bEF1Tg7srFK
sve8ZD1N54lRUtKXUakeWuwMUo4vKD0OyziMqYbNOAs+UqjPlVjkLcomSTpt3LgxDyO7V+wULTMj
XcZOis0kQO5zrJF9sN5JjkhGygn0GP+BZpVT133LJGYHbfNQ8et6WKyeXhWRaHoXLMpN/FyvHqa6
vJXcs3EBY5EM/N+31dYVFmbXm9s0X52o7XfpRwXwZMOqHTKoH7am1dsDNlUBSABD42Q0KPAf3cHs
9oSQUC6gk4eVonHsX2slqP6uTaopgR31JQ9RjhRRd2Ntf+af231XgGk8Kca5+HS65n2AXdAAoL5g
zWnXCG+z3HFxqUNvcgCoL0ve2uRqsWPHC6UJYyYTKIazoVq9jhDMqIXvvKh+g/Aqglajx07D4I+O
rIRKwBt9CViL7cdrsx6hCypUUm8qN8vK/xjg7iqlmT5vqsekwKs919VGTv5PEsThSM84kwiyL9zD
/jLJiaOiOEw8PXAIoGvX+y7NYRcp6uhTKabgDPQ68yzB7flM0Q/P57r3e5bwFFH+JskfkvR18fpv
NJQyuImwjtdcetr5zI/i79JTtZSa/ItVHgpg0IQ6/MaxBvkDsK+0DhxYN7NlO//Y9xIrrvfvEi0k
aWvONep9kFi9wNFLtpRexgiHcrtGtX3vOQrpiTOjcP2dvGe1PmQK0zeYaODI8XD0KJ41vOBC6nYj
YtL0ZDpuuvLJmaTPm+7HPSu+GGQvrku31Lna3ilSKOv+TRhjiFgW/VYg82LzSmJCkag2fXJVmOkT
/FIccPaKyEycqdnqpAo49Hc9/L7YaT5V7FilYY4m3tmmhn5+SsgpRA8KFKXw/xRtTNlmUicnCHXB
aYnOm+aJS7Ws9MJ6UBtyQfOHG1/ZlMBj8ZRBhe7mu2yNFjPWrs6PQg+MKha+eD6Z/iD4YrRM8yQN
OVPwGfZgtOTIat6+mQE09BgJQuk2l3to0xk6WwU5UnJ5kplVuDY9CUT7QQnjLA7lAir2UTrD5i8e
F5tmbzmlR8MNqO6ib8wgm6Q5puT5uSK0u2+x0Si8HRmdWy6Yql+FkmsnTOirHyLvuhwCnRn9yZDw
XV8rD2/4raEHktENtbvCEsRlVtekfNTXbcNM0lSszvf0qb2CxiWzUpw6fQwi0b6sWPclsyARAbKO
8cD/8HQULUkmjOJW6FS1StZWmdasYhODL7K05KpyRvRtEWzWa9StZcV3oJ6+qURu/PR6ANuUv48i
+AieKmt5NhceO8/gZJYhVKM9hrYEV07CUbF3WXDqra/R6PGZuaoTicnJUSjzx1RiOQfaoPTLyUIn
gxof635ggHZZLV/slcVVf2PT2hOzzcxhRhomkf1Gr/nFRnkuOxGfW+8zWVrn9MQeYVY1lBULRs57
6VA/i/A9LbBsIxH4bAXHlnCQoXAqJum5MT/TW7pr0Ax7gPfMkk7NtN5k2QC9ilJPu3DJbKMms5px
iXHzW79GadbC4SQ5C5BYakLhx4H+y2BaSSOV2qkVGuepsarjEMlLK0/UVD3k3JXRKfhepfmMyZb/
M7IA+lH6aPTjkZpAfI92c87RRMgSXrHjpwYuxJSp9jXwNh/hrEx3gt+9PlWPrf28lPE2WXc6eFOD
fxIYunn4P4EcXZV6Q48ULjgSZ2ijR4s0F0w1s5gSXMmX6nGcx0T6Y3ElyApJSjLzwuuDNjP8P8wg
lQ33K7yFXJVFnE1Hvyug6Xsr7/2CZNLLsxpvdMiM9Ld3JsucApknIGaz/0n3hhepIhCI+M9IQZYi
iLnLIneoPAd9vuAFtxMd885ZYmcwgZM+mFcW19xU0iWbXAnPiuNVbHdzcBopUf3GLA/IAdqs9tiu
exR30r71P1EaKPDw1+lF58HJ9hSiK/G4t4KXtmpITxRBDLNxHdp/mEAHgBVO4npe9dcFMQSIyKNN
8O1yNwLE1obXCaAsKCECXHCQdqnFwCC2UpAgU3ZCRXaiamO/N6hx5k4FCdvVijQK/qdbncxmB85+
NlfkPdx4J7igjO7alw9zo5bsVilK4nplY6bIlw+cGJ1T01f6FnUPPmrP8HV8KX7SB7EivcnnXjKX
asmAWXnStbnI3I4yzJ8GVj9dkW4gd942crjr2wgFTJyOQkK+fHMnYBkfu5+yibEePpzu3iqbakPa
1iqT9qocAz8PZHCMTGcW48HxUTqJpvLm8liskdPeBZac1WPsKLCf6f+USTlzoDzjFMtI/dS6+0nk
ws0F+V72prPTUrk6rOoj7UX3EpxTt7gqtSL3E/nVkaPe0CHUHfVUDbTLCWkOUIrLqwn3apGjQiY+
uRzQgLI7qQxFgqC+OcJjGLC129JKCV7w7DZSGrBPFnGsfE1y81W43Xk2ei8KBlFU/rtAfC4fhGzp
fq5grmYrKcPsVZ8gYK7OTDCXm0mPoWQuvqTN7zc9j8iMHy14CQz1TSKoln4GhCHYS8/PtCsKWGIY
t2fX7bjetaNCOKh4C1SAKn9LYRUon276GV79UXO+KitTiPiGKXY7PIz/y5TFirtE/xjKrczpaT/l
qgGUMJDnHWPJj0FSU1l0/JPzx5skpeOxoncy71BLnP1vzogcu/WXaSNW1LM9/HFKrvbC7ytVWsF1
bLzkC5RcEjrM4FdLm3SYrSZdFXFJepytS0A/9EvGQRwGGWPX431OA7n4kIJ+hm5ZgIPvpGEEFkC5
qkqIUQihpKptWaQ6BLnZOPW+YyxvdtYZkdO7nbSF2x8a/4U+2uFLons92/yEkxD252ZWLQwwZhvq
l6XGys0eErKSk4TMEABplxw9BhIzwiyrX1RXiWYT+zA5U22XUZF83gEAhdjwyjFQET+XoC+Dx8Oz
jQpM8feVxVGPWYRAdblQrBamLj4bMrrlv56vpOpPrOPojQiMB8a47fzwYMObFyCsywMdIu8cSRWh
EAFxHCHKhlqdVGjOlXHnHvKhVtM800s/MA8vkm/tBx3zO4b5PkBza92UaApZmWeSwiyi7hjIXXDj
g71l2MaRmd/w+0bMCEQ1NrrxmjecFP31T0GApu1fXKwj2ttlc2MPhlebHpb+PtgiRJ2hd/oU7rqf
gT/V4EKUM2LoBnZiLN56OeucWV7Lvex9lTBp2Md6ZaZuTgmEWauDBAfSnT7WG1glJN1I/QCW6m61
tvXtFCVqx+i7Qa8yka7lwNJQwmQh43Flq5RJ0BoHihlYhuOTAE26I+JLlHwSQ5xDrwz1GP1uw4zB
85Vnz6eJZk+QUpUhW6yxSBOJLVDSMJ5/FGLm9F0Yp3UH5k1BozQ1+DKQAGvQueqPYZI2wyNZohKc
xb9VPLljmBPBdLrzgj09mqS+bAnBlYMPTS7msCfX9aGeDB5do1+xVuSo5IRZWY4PzGCxxmO+cWbK
Now7toAIyyjnu+XK7i1U2CeEhQdRKO4v4ASqGEmauJPhMYR2Db+4bYfxsjtm0XLrf9spnyTDFAul
cj+OnKigPGaV6fbbaLP97hZm4vpQgG0DFiaXpozRiJqKAZJB5TldiOzIcNeFES0av18du9lEQVzz
QoL3OQuXbRD4REhby4lrQ2a/XQnH9yJC2BaEYtjpm4lE7tRQsq7jZnpKdhhD4AumPIEHGcw2BfD5
OESPGESQEPKbcSuTCL2Vv2sSEbR5BDkuLRELTeEApOaUdmcSki0xRwS5JDqyFx2aq7xCxmYzvluy
WIlrcM0cUqEh5i/ChWdPGIN7WaGpnzzElFkiKZLHbf3yBYjzRijiCdTOl6XiqsGoQBCSoBzLdvaz
Es0+hpcDe8Ns92AJmCjp3DV/1RQbqDRKmbqCboai8g9cv9yD4WIgL3yfjAOBiPHa/4Muk5dlaWZJ
zd3pACGibrr8w7iUfddPWPJS98b2JKBjKa1nzfE2Q0ZCpxlUx6Sl9wSdkEJ1CD6a2rBGO8PPXaZB
gMXX5jqd5uB1rqxiVOCUnrncOJ53XRIN8OFWexZ7gVqAFfbFgu+L1kZRqdcXHYWNZrLjqY5ztFws
uT1D4XJ40JJj98GI/G2hgGSMgBZSdDiK/OGcHv0NpWIg8qyAUWB6xu5nh8hTaGbfvduvoQ75QjHt
ouppEpnv9e2G/82sWdGtRxXvJhPLaWf4xxG5HM95Llqybsa8OyPZAMEEn4l6B43R2q3cJwTUJtcm
3alAaW6m3hZz6RWUBRFxCye7N7nCavSAlJfzpeK8vukWpM80knar/a0OzTf/8lykXVgt2XYLJ+e4
P51BxoasWCqC2fX0oiqG+LaveoWG7IbAZ3Gv/r8ZH9NB3C+jjoe5QR3FQaDy1CGIhr4EVMrzrkPC
3ACYS9ujBpDH6fPEWnJEaTylyUz441UAjamJdAyY2++iBWwOvcge70bABBTiG5Kqgu+66uzU0/BJ
B4OZcUaVigcUPIRG+2ZfU5dQpgo/viWaiKDLMUQaDXJisrpkgKl7KloKTHYqkknCJS1aXOZl9AU7
0MrZixPRPjEEpEWC0g/fMWiBAXZT7PCpu7jm6AL/lO6SV1y2wA+onoDXi3anrBpSKDm4d+c8r8XR
NrN+wolQxYAgyaP80nkcnPmJ+391BSrfIrgTiQWoLz9kN1KxPWFTqv0L4FIiRzJTHBoZB7jniC6G
JVU00uzooktHS+NSvP9G2ApGI9F/JrUWpotzrdaK7I4ce7g2cdPRl8hPwiFpG6jrPK3ySbGBwOWi
TIMBLuaxc5ruxgg2VRATIW9Ow/QmUE2d5iebjKUSGR65+qk+tf/zXcQ6aEiG5q8pVQ2MSE8xh0hh
uTZb6+OpkTgRni19w6Ownm6Y59aJBEZ25XV0sqIl5WfkaPNGZ5ULyY8/LQHgZC1DhbKfdaojSXin
PhSENKaeLruAAeM66i6j7ECaOTfbDid04g0vot5OhcHTBI9tSy00XP1VqrFzOvfKrYyX3lzgpjFr
xfbLBHgIOQlV6c2/sXsrnqNlyq6Poue9i2kn5/v3+gcLcCm2V6hn//OUV8iSHxu1+ZVy2laASRgF
qSPns2+y1hmfMR8O0mlY9fN/QIISItTh7XmHDV+y0ghsmqrgx8qGGJiXS7IOcxBnwhWYzxSj43Uo
+aIUVA7p3NXBluoQpXpnOc97w5z05NJGuPMm9QaofD0snkDBQXIrD94zMIFc1pfvt5bpXukMntgG
kZgY5M2dfOW3fGvxMGHw9A21xeCGsKSbAAG7d6yA7pkVreYMUFT6mo3YG7yBlhj4GYEfxcotv99q
zvrpqEp+/hNU5Vjfj8g5pTr6HYHc3P/Of66G2+gbO+NdOFVFkFailTKAXszKu33+g2sk8ZFXGUiU
9RGgqjVwY2QeX8W1R/ezg4TPHFb/0x9sjN+WMGpbKCmrr9so3q7WhRjiU60/jDVL5V3D+e8PC4jB
CamtLOgG+bwP7zT9SCR7wxcMLpLg/MCnXxY0t2Q94sYRBLmY5EQAH7JgdctD7qVmVR8ax/ipJzUJ
nIl95Zw6F4NPV92VjsPGX2vRdRGqnaqzu36rlopmOMnt7oiOKDDbVbZZF5f7pFlW+Dy3YVVtyC1X
gvRKpezKQFhvQOpa3/oOEd+A/By2h2uZAFvN9BoYpZp3LEFXJ+TdHOZOGNTXYOgLss8YODpxlWHM
GceoGQBB/EI8Qwy6Iy4GASsNBQn6zZm3zjMaxMm/vdGf9n4QUkLJujtDvIR/HLZPb75odlyjcPhO
/XPKLKGkokcgjmckq2dtxGDfddUXv+Fy7oP0k66EHrlbOhBPdX34xLJKHNQ89Fe3914n07Qt1Bcp
HDQp0iJrzREodLmNbSogYwAKp+0VuqA6YJLHi48sfd0BofSUybXzGf2S0ZgMVj98poNAAj0BfOGY
HTLB5ASdce47aMgSniH+tcACpdvucn19lvjpUOVrZrX3mubzwQjaTK4moUGOgwVsOLbhMjDKWXed
rzGDRoKUIaB4LqGRMYz7WXRe+O02b/jzWp9czY407zJlODGXZbFR4D1wqZIX/D8/TP/BvNlTq+rO
x7psUDa7Ck+idU7A18MFOfe267N36XRkN1rasBDDAXtCDV7sdmCoCacNX9GROL0wP/+adUOwzoC0
cmducmaFaThcJinhMS1lHqe9BZT4qQGm3gtI7oV0cirP7TPv4YLfrOhhaXls6brXqF/KIZLqNab1
KFCXYPmcHPaiyE6zwJi0p2Q1NqpMgEJyoGW7zfkGqgxmo4fGsWNJpWB5kccpS5mbn6Q3I2xHwV4I
NsLut2BC3qEYwZC/2bgHeiTsAzPi9ECU5iEKbrejMeqjy34rVnnC2RZjOJP90V5C5hhQGp+6t9KH
8fildiXrIjrRTjXCZOhjSGul6fPuE+KR1ciMRFRnGRQMZ7zmqZudKL9u7o5/cPGWzdkT38+vbwAh
4DL5rreacEqH+/X/lfRMizrZUZrKGIFlkB4sb47efny33ykk4hXQyhfYDH4IPPpvePT88RucbsC4
uRhg6Cg0J9vF+mL7SL0LDGd8lenCb3VSMHSM3xEmnmwXVxYRTf8tqMfG3XchWQBnMotfNcqgOKy9
KHMqDLWLLucapd56G5CeWgccAPn7agt8Ji0GMpxwVpGzNUOhXf24f4bpY0hVZQ7Dys8kx7oqhrUh
46gUpcIFRlpjlxvQqLBfmvYUQtisiRTxUi/gMsKUi8QrtyQxFgvCtWOO6XJzQ89YX0jYKKH4MQYc
rcLFRyy8uPq47Q4axFh5DLeBlgMF6bSH6901DAv1AATYjwrGvSaP1xyNlPqem9t3ZYOuBhuLEBU6
rRc56aBk8rsEDQ986Nvk6iE/7N7Zz2qSXbyDu+QVLhW+uDW8Rbw4afa0KcQx9J91GQspOJhPeaCR
jLHvYCDbaInWZvXWMt9ZNvTO8PKd3RwIhjL7Lhl4OmNChRLmPviV2NI/IN40TPKWHSoLgoF8FieM
CLMJVqz+k2t3Lk9mj5hIsKQ1gyIfaQzwG87GpJCYNRG/ZuL8EJbpCecLyQUIebOW2hApY1zWu9SP
R3HoI6GTlQLWlIZZ8qr7wwLgTion4rMKsr4DieYF7lozAzev7eFqnH8n7it+qHjHjO+RNzm2M0AH
6+NxrtUzMW5w147DeJ9xmTnCzDefBI5OWHfcadvIXd4FaZaf1fWK6cyCfzSbyoLiWqmDqPrIJrRo
H65WTyRu9m25umO7wTs2oIV62z0wbBDKdeLvD9dQASRhqvwUysTbLO3VilNcEfS3KTDps7Vay1A4
ScoKVvXFK1XOxMmduYY+ikP22GWo9+xUtY4mRtjUpdqd0SiTZif9jtWm4JLXItxoU4M4qBBDDRd4
n5Va1iyDv8pikccmT0qmYtka/JahnNUCSc9YLHi33Epp2ffuxtdLKQGQDY7htGCImR2NdChxHc0Y
fTgtSP9kI9hdg0gtGipMOzv33MO5yzy6EPeRcdAp7KZkQvq5vguXpPxO9K1wv2hdV6HxjShkGWWq
E/uhQOfdrAAtWdQCQC3hiI7jxdmiHMmalGOmQlCchRadzJlhibt+lHJKEhnjXSLZkxbALjJSRHBQ
mjlqKIB7nRFhvah2rs3iMB4GM5EyyO1ZrsxqJqB+OwamPBJHpOscIdkRBfkHVJf/fmCVhhleXXZP
24/6HvbGNJXd65m4hCX5HUrTBW49900Ziky9muhw4ujX1G8PpUchPbrhI/Y9EsT3o/4nw/ZshMUK
vw/ays2EhjeMiFVUkNWLizyZQP9yafnB+UBH588u8g3MUaIN6lJWfgaRAYjme4hvGs/IS5ee6487
YVY485QkhCQ2Yo5JuMn9zqyS5+oJQxqA6PWuVoheFgMZwrBgDYYTfaQje2bqEIIooh/bnvRzCZRD
cKZdTPpx6fV8K5HM+il5WpLk/9BYcT1bTNl/o9F/5MkaDxj9Gk64grJY78OaXsfeuQowqJ2yGBLv
JPTPyhGmoona53bTwtPC0GCMGmjPQB+pX/SJqU2A4y6msuwxJvcLSdjTKecWviSroRK5KxC79iWA
JPvlXr9TUp1VIN4xL3QpQpe932x9av5bKfNWMTarAf84416DbMalXWMEwsu1gQkOft5HH32GeIcj
yHJKuVqCxQZsAaM+xQY9czUS3eHi/GV/jYIKWyB583G3Eg47bumoFhPdjQCZv0o3Zhns9iiF21XK
Omir2R9IKW1iavHH80SzT3Vd4f4i/lelQxzKtFQv5xzjL36Inb4XpqmtRkCpVQKJlH6Ae3F8sUWy
6N3Z9Elvxx2mtnZV7I2/+dvcnIHAqHzffbPZTkfPrLTUfnCj5IelJxpu7ubUcJS9rk3MBhSu/fL2
2llAqNwckMYNYhqU62XUE629pdNO3pRibw1CX99YZ3JHKrmJHLM4Vis9Yq78zebni9PXpPc+hhVN
86r1TsBh0vuKj8FpalTPN+qmGX3dkNeDO0z+ViArqIjLbd0tPkLOqyyBoliIJbQZuKTguc1Rm55e
s/8oYcsO5+eQuZzCe0ngWKRpRAO895TeeUDjNplepy+5ck3XwJmp4ltvQlInKoFeUF4WbjlBguWJ
GVPZdxkqliVxJpTf1B5iN21U8e9uLjR6/Q7fk0gPYwNgrqJKQVNGwU0QX39Oa45IgwNjmUxfp+fo
oHw5ox0kC0vqFpfHUxzJWuHdjt+uN+tXPW10+Dl3K1Fpd1I7D6DGCwz456XtdPvYqsWnWslrJ6Sy
MZOg5HrP3VI0LbkxZpark2ceg6NoMiPqEvGhDuYu/vErpQVraV9FdKecwlUo97tvVNOMLb4vydKd
oaCDMSzfF+g5m4bPdCKehWaeMEnWlpgn/engS9dkxtYUSS9+EEfaiccFFqi9lhJb0sQoTLIJZN2M
Bxw6gtSAYm2i7Ijlh9ZzB8DH7Q+EcH/IsK0thNgrmolOsMcXPU9yAduF5acuCoLfWoZ6BXtKo1wh
2TgFWDtAWbtzVkrfntWY3uR64BxvBINAp3/6s4Mo0aOxL4fqP0HyVzroCiTseWk61wPYosoSYI6x
r47EqlrPZBJPWQ7wXoxtgRHg+skHZEmd+39APLGYSQYk4FawJiD94LNcfrL2rMlvLHg0yS1qBBG8
EFXx3NC8TochXHRU979T0378pzyOyWOE4AASlUE++mmMFxvlUFAnphioIwXkv4N7tN1TGDzioHpl
aDmkKxINpl9VBMR0RWLSjRslI8RX8VF8MNi4oD7S0WRoo8w0IIJKg4jZJZkhMOMtWkijTXQ4QbR4
incgHyX35aiGUAS1W/b0IxOS/VJvbDsxTdyl2qcQV8KK+u0OXFq6kotghBr56uzd8MQFuY8VWN/Y
PrU8QXMtpjBFNGDy7eFCXbaUOaZOGswNEIGeRnIiEzmChm3wzGc9Z+XP15qv2hypq0iLOPhZ9LVJ
INHkZIrv7TkiH1eDY7+bXj9CH49dQ5QGfxQq9cvy0MTs4/hgF0TUeFqaR746NWFPeMOKJ+MLNAG0
9QblDx4SpPVXQ1+AgPPoKMnvlWJmateY1vMQfB6DuBxGr50vuHh76IF4IOUsvvSHCCeKBrIJnT9r
W3P0b8PqBrZQCua0f9rBoRaie69nUXknLtz65QzYvqgCXrUd4deq6P7/AK7Iz6i97d4b970YCLKz
ThDfIRWtUXpHR03/QkVYoLkEZrxgaf4Les5XyJBV/hQMoUWazmDLv10BvCoSC5Z86hhMBgeqoZGu
gB1LCc1o6XNvKFWYUj7eljMpLhG8mbj1uYw/T42coSMVCX9Clyz6c/Smf4ipmM3ggMJG+6+FAn1k
JFw8tH/wX7WfUyDDiNK3eEmaAiRSD0H59Vp5JuTHF3abJZkYrDDw3NSdR8ILWX8aN6iI1Q4Ht3BS
a2rYOiXdZD+vqQbpba1DbeZSOhkIFtS0I0voJxqrazQ+qxXQXAd9v7Mog26IaFYB1tnI70Q3OxuQ
SHVfHDyDb330EqUzKqD7m7IF6v1QmJpahLtZU7dzRdB3dHEgUE/C8NV6lQPWc7iaJbUo5qnIvVvK
QzhJOh2YCnftNvIASQoFLrLRIaionRocju5njiGD0uqAHWaUVbLedaaEYxdeWpjKx41IcZ+8zvJg
pkVbFOUFKsx+iQ6q33wO0xE6Q8M+W6tlaAqf7kRE+bcn6aICaCkHy0NAeT9RrwZjts47ic1Sdp8i
cf6Tem+oziO4S/seGi+caD4FaXt1ziGXZrBwlA8Rr3S83pd+0idG0orzIrmf0GknW5UGsVSGn3NK
xPRDhNdDCsx8iLwOXfQhupapqM3BG+/w/QwtzSajV6fgdkgaT2NmbERO9Z82vcqM9Pht8vr0fslS
SGT+1/GwEk4BDhxY0OSkNAJ1uuL2zXnYFacSt/TAsxzluQoxKc8+Pyx6Iwh9J4sIUcbTjAzhYBGg
iUhCV1FUfdG6u4yEBqgn7clySyvBJLfS6vpav6gLbFHq3NxoS6gPFB2ABpJfl8G3Sx5ZC28YC0Ez
BdosCqRxj5/aniGAgYaWOmziTPco72QgOveQMk2givkiGx4Zj/fn9BNpTrRYIPBM+aAmCrAtGB3d
KbDnnXRAE5OyukQ7o8sMzPKLkOwSY3u0B6/wUao1H3EJALXDcZFMQ2CBbVs1boi478VW/NPwlrcD
BLBdtuHnVDp6mwO4TmdleJOYznAPqjXWZBX3vyo+Jt2sua0tyfIzAhEWj6sqh0xdeWMY1Y1SXIud
oOzlFG6cBpQ7FqK96+g33rBsGtRsqM+wxW1tajGpMg+7fSR97ZesiCm9zIAdf7rTczsS7IG8x1dI
X680XDBsEo5e/fE4ghp0buNRteXtvqoK0dCl6AxYa41uSl5mOJzuph+QWpHY/nB233tfVVPyhfq9
E7OkHmxhxGOU+3IZjszcXVOvLqgZhvUGjh+V9BhEYuwOM/dAGVikNXD/IMdQx4GKccitCkscdn/w
odMyXo9ZGFq0SlRb+vhUdWgBn92Ngnmhu2iJ3j1MSdrQGF/Bp+9cUz2ltU53CHNf1RPHULKDdZJA
VPOF2dhx1V04w0Kcl5YSska++dP4Ih7DVv7acmY1qE/ODl9V9W7oLdqPPovVmtZeScGcjPEVaHDH
Ha0fJiZ0iDoBYeBy03t7LVwPEFsDbHBLD/sOV9mQQk46BeHcKnypyI71WT1swcROVgfL8Dy7IdSh
L/l/UUzC8EC2iThcbV7xdmyUkT2sKnzKY4PRiy8bT764KUzdPzk6U9GEBkBV61fAxhm3jT1jQdm0
T5kTwQNhlqkYKgDR/Kwoe9fz1QrMm3hBF/o8bx0mfxemcUJY6ifXSIaQ3jiJCZfcj0X/oYvF5tWy
0Xn16brpJXV2bxG+aM6mA72FuDkJEbf+zBO1JL5Na/JvKGbUO75o8LN3LPiPlJ866leoSpOl8795
RrzgMEjvInknGmI/czzQvuw2ZZ6U0IU+qkhV1PltgRTx5oYppAm4aUQAk0mIuCv9/DHMOeYRITV0
F1RiJ+TV56DLtdavqM0v4LhbiDuiaZUJ5wn8fJAglUg2FcSs7wjB3dKz2YGRFc2tgbTdtYutvuRr
QhSd+QAahsBXtOp98xnxx70Xb3ix1BMPj+iriKb+44hU9sDQr48qPDEGbFlBuCxoLR5f4/ezEFpB
Q+V+nD+gHwWLlEOC1kYkpr7WNPwleorbO00uxosEZXta7FhoqOcqtJw8DmP6IxOrA2Xb1LmPV03Q
bgP/MMB3JmJuRLRKg2t8HzP4dSQZuFTZ7NLbVMtsyoz2Z+J1M3h1jZvk8D6dl0spIghOfE+6m/jB
BBIv+lOWy5kVnz/Y+oksncC7w5s5lYOuKZfseObtNoXOCVhNQXf+Ts938YBo4pDxKXRza1e6LXo7
vQgfs0zuHKcMbAuiCfqZ2qesGO7JnyxEYpcuRcY0TagHvtWzE6XtEKuff67fwUmPdi60r5VgEPhR
fvuhpkSh0lId+GFYj+2HEz8VB+lMPKS5NoBdj2kYtXu2VmrDX+VmQ6wpvQ+ZpPA6atMpO7Dic8n4
+EvoUI/XXpK3XcaXeaHCSo1P/qIcoofkkQh+r6eFJlhHuDuDcYl0EX2P28d/M1RgmbGaa+/SqVOz
gfhiQYGwAPUDB+bsW46QZ3DLNzv0vzj+Fihov0rtXu3t5zccT62O25gUXw+6snm68LnuxljVRi02
e1Ng9SuxXBcjSSptQsHVrRdpoYaokULZSMEsdH9R8xsDgHrg088XQgMtjBKmKORgwOv+aSuzgZkA
b/zsfiZe5nu5Zb3oYzd/AQkxbPQilDRtKEFWXp97HqVBFRRJD8MocIffTRtLApIe/UcteLruXcHG
c9pUWVGA3Mwv+hoCaWeJB/SoNGQ+vlBDXJfeIf7i4CWZw7lyyWW3J4Oe1SmkY9Gsl5CHL1RRVu5c
INK7oONBFqxDupBIZG2ULE5tFBQYfnNrQbDyICLGc/ui0U2dpxqyx4aOfmOlJ6yElPazVKCpRGhD
9QXFQzB+lDItxfnP3is7xLnoAgs+XBPTLWubxKokER1luodf3Op6Re2ODem/chtKl8p1fLlYHptK
EXAfOViQytV/qajgMdJXPeuq0RL57ZW78URRf8bMIOXN4FGsB1gLEkkZvx/c12FkxJ2DUROQRxFS
sbevbma//MbvKr8upqhQvYXyg+EemQl7TtZpNj+tA2HG4NkzS1LqktjWR8i/sXnp+uU18gnmyQh4
L4UrJFU22lv6hM06uggQYMUU9iZ7pzTlgXvrG8f7ySPl7uj2n46zwQESi0NVt5M2X+/4PSTyB1eX
V4ze8OLm0vDsv/r2VEEiF9Kg9m21fWddsqG46LLm4LED9+4pAOGxogGNq9VMqjvFgSpGvk23W306
TwYX1ZLlEAh6q/GmZajtPp1akuwVyDODGuQ1QVur7M8zR4v03NTq0loN6X5s9IaHKKGvYydYR+Vd
axw/kNv+kCYq29yYyzTxMCUnJEouYfJ3DSiHQxlm+lFqb00n2j/MdgS0nsd0OeC8RF0NwJUbGup9
I+kcF9xjCJ2BcD/KuMAUrz7hMJDycBkAEHz9HYpVsHD+1j5rWsX7wnV0XAvVO/rAEridDFl1iwGb
hCc3K3qoIQGeU7wqDSBtUEXbcXzY3iufcZPS5FE7y5CeJl2Zdlqtzi64C8QTflbZciew+JWS4LQS
bG6u5TTCjmyN+TLnWVysNkfrdcvC1vUioejoWUNKltIw/GipIB4Ou7PO/5Ryz/rYbzlUr4mOnpIG
7XrFq8qHjHIV8R582WrxRJ70yZwknwxaBCaJI6jVbC4f+MYrqojN3HbwdoABk699rbeH58cCvEQh
ShMxfrONDm6KuZ9TvYXryK20w1IObXKcZlOWQHJ0O0DIlTA+IHn99hWn/F7VCsr5jdHCuGPyQCs8
Jbmg30wIacwgyf8FIiJD/fVDTW0CllKSH6AN2YaiM3M1USrMx/ne7OVpueSSFM4TB2yiAt+cLTzT
bNtxYnou+/fv21futeobtesRiDfVq+cPljD/lp4WxzKiHK43msDUixiZp8MAHCDxFZJlxPzI4qhe
mzzGUwYoQTMFV7KefK3+q4XMtnFOCrPBUsPPak/2AU+cQCWQ+Ks+hKv4f9i3X610M3ur65rQvrwP
LjAEjl8E6bb+p6vlwyzUK6st+/N/lhZlpyscZhPgycBgD542Qqqy+/jVTvHILcjjax96z/JANekN
282dooG3mWbZ4NapYEQfWOGwqbNcmvdFnXMZqkNTS7Bx6Fmx+OvIln4LjBOuRe2BQ4yvSrlrTDLA
LSVp6lJ5KzRTN2i8JJ7Ad+MkQBHIWDodPqyvsdXaLrm2d9oSzyIBJ/N+5m66mFGx7VOXq42/c5bE
Gmp+8rhvSQoGmu8VsrTZfgUAtTaNLM2Q0JoAEJJbzKg10vuVRpEEaUY9rDwTnImxyLnThMBYfX8S
+3dnCjzD5zxIvI0WVzPiJNgT8du4NbnH4gtYmtxNMNChgfEh+r/QiSROXhj2kqE64YnZiPi+TM1a
mtdy6FSHRfLopJMmir7iqYNoC5w5BLP2r5VZGw1WwlcbNpodZ3YhFLHk+FHZKSFjmoNtfcWbaK9D
3QD44sSPPhH1dcC52U2OQZylwxJLh/eGgrcIGM/RqcTC7UNXDe1oN8q0wzHwYdjEDcuRtUPlQivN
QadS5jY871+fo7ylZe9tZOJaH6OtUdFTj/C4vr4l05aA99IRpjSjIO5TBzIjglp2nQDRCO+5eBij
v9zvTfo+zVSdpISGDZY2TNADxLSsjKj8jw6W1NZCIdlDsDe43/p1iqAVR2gOtQGMrmxFwrkwCw0b
oIxIzA7Ku+5etsVnc8aQB22Ki6ukvK6DdxMNUjayjxBjSJTeKT5WZiUcB2cTWsBPVSVja8tx4e0c
pRAybXeSv2AZdcsNedoQLGhP3/LiCAcq7ajFISh0nc8dsB2kArNGP6eh2u9k/vUTJ6XVdUP588bV
ePjfLMJ0Ws6fUhTqrL98P34n3NbZCqXvSZSP/E4ys294K+1ANDSVKOzl4pf8r+QM53CN9+ebZhpC
c3UZVfO+dOVxxoiOAIViGtSO7UYLb6u2IT9+OMDkOhbL5jygkbsO+pjKt497o1/H92BdVwnxCTKI
P+ZOeiI49eBtpa3G3y4nt6+uSKSJk7/8Cvpr3ohHBmXVQZ2K5dM4usoEpbpzYqlceCsJxWhacBto
4v1YkJ6Z6MO0zHaKrZEXxhx6ack2H00rdT4a/Jo6AAwNCMuqsUXBf1t5mdKZiGGxtWgbsmh7HkRJ
wG5AxqGZQyuU6q+fQ1Jr5+ZngBM6tL+bZTUtCprFqe8ZXhtY8kDxY9eyl22k9y6zmTbLh7F721Ch
HzZvUUqBher8LeGehiIylwSkUDA3j/bF83tl9hlarEaR7FkW0lLM7Vn86WNbZ/M1847cjXzyfiMc
uiy4QncZOzG8nJrYvnKtCrbHrpNdSPz3ZKhsE5AiD8Ki85lM7XoVsCU5cntxExrpnYzDlhMaEfzd
ZwJNfgFuqXAuO8cAKXw5Nqnas6b5+P+X4/HSkxzwc5GByOeBt05ol7RZ6Ly+FzH1ZZn3ctCuXNcc
VC3yQSpi9NM/xnjtmx4bitXubNOa3D97sVXFcGTRzarVaMTVdyBepk4E/BU/v5y6a44UbyqbfSrR
XLC6QSPk/awm3aN26jyrLvlQteT7+C8FqmBpgybdaHYebZRrimVZTOxd0b+O+Riw33Uuvb1aUk49
odkl49EPWVXdYx8awW28L6spt71CYxJYah+cZJeeoROn7zfPOsRO3PQ83voaLgo0BozKJ0f9j3n+
7kSAkVwa/L9Q6soI7/BUJ1ygw7wOtfnanyPefpXtfV2r56Vn6qPO/2iPU0NUgJLTSkNV2fiF3BQt
EwscVyU9xT3Fv6UNUslWN2SLWjouRBfCY+ohgw/xj7meAzPo7K7h1jDHvZM6AcLtJVvGoFjSBoEP
z2pTTqSgByVdzay/GJ0OFuGcjBcaOwnEBNUDhcSP181ttTb+I9pRWDOs4A57eJC5fS6pjf1xJNoS
M8WYnArw/LsWa623RbFEG3wZ128S8CpmPWBg/GMKSc3Jywa5mJsD4EK942iWaXSge6vCOK9VWLL2
rQpg0+jyhU8giObeWFl81f0kdMPnyKstBW93+YNYJ+dMU5AO0a7pYyPk0O58/u+onQAUnxuDBDLD
0vdfQQBZug3/BQ6qoPZU17E8F2XI+GhlF3enElf6ie2eAu8Ym5BSmhej22hNG7uNuvi5xZ1DRVL5
/Ch7apDEabR2hl16m51yWFKVYxPklyeU5mX3jtmw/D+n7EdWB7r6vE2eExIi1klT4NAzwLerXPER
JyIbykiML4yIsbtXfgctEyMnP5Hfaz+rQUtR02mxghrbk1n+VwwOgTozkIfEhakGkeg69dL1ETG0
j2AODS7KbIew/kFiuDIOD0kxaZ4HJHlbOx3ZfrxQIdVkIazyBuG4bXRIrn5RSPg2SUr6LkxdyGRZ
CnmaQ8r4OjbTnRFswhuoGSY90VF6cp0qGfLgx3QwEDbshfhNyYlc52UhAmuM8aJCZXuuDkMbqKec
eGU3ruUrZcaflwc0fGEoDGlwQL7JbeKg1+pWIkaW8gjpqekJF6NgD4YPUAxpKE5e7RBeIBwe+X5U
m7R9AenmLnV39CfwPwePzIaPAVkoPq0h6wDUS/OcbyOy3rvCduZFs7OqBygByyDDWvgyTwLf9iG7
yNMkmsSqqiLDMCvmvcTDlBt63jo9KJT/AANgneOVNtqKb7ixZqMuF3byzBh7oCogIX4h5/B2lsmc
yKoSxjJnllnUGu/P3ZjlVtAuzsUeK+LSXHipV6wP6E2IMafyKoHXG+xwYk7daON3r5TulrU72VvK
lsBCEXQkIhjcOL4/Dm4ePaZQjeX4xIEyQs0yUO0Uff783vpzn4qIsMhAjD6q3DSHmGjWTSAzvnmZ
4UFMd4kSn3qimOTqH+uEqPfeSDiDUX2fuech+k27yk8vs85tCcMB818A1/14VwDBMHk5kVQpbt+H
j1n+zfzrcUPaShQLetV0NSmPWGxr3AA+ohI2pKTqS26UC6U0u6lk8ILoGXKNMkcH6qiNSaD02kyq
O1bOYKe0SpruuuWlIxw+bG984aOV/3pByXqcBSUlRVfeyFfJcKA049kGBlzq7ADkAGiMnIHYFaY9
8S6Ti9EfJz7A5ajGMoDgtFf5ABe0e8g55slv8yFLYpwtm2Npgo+ztwk9dBwTs1sNkd9ndsIu5Wjl
DLmL8aXNbGexRf063rTlNaS4dFIcglhgr8RfAdDH4qgKNffhJufvgZAkG9cObWXFqPCrg6oEq8um
ByW1ncz24+LTIqLJasD1zZRyWY6bID3riYbAaDYWNzBmTEnacJ88CBKJjt75komhHb+dvrRaawyG
plduW8so/mOXoynvpOuf8Cjj6VTXs2JvAuDGclhtJLtS8NP2pXzpELQ4ZDrsltJGuHmc/AARFrOB
4truXbEkPYyfTV13FB8KBDLr9TNbkta/PENKcy5ssmKjZJy/4ynPDuxw/CUiphU5W8xPvmqkwRrm
MXWg2U+ykHEHnXdv8Iy9tk9NcDrgIOeU+4PkIPDWaZazWlsk2lP9BrH3XkO3niQA6629HwmRLKvz
BKHbcJ/WkF5w8Zk6GvBfhtC44SsmhXh/o8DVHe1LiUojg7tyMBRsZwTTigqt/fwDZW/WfedHLjLs
05rffv11V5uyKPCmt/iXsvdxhpWJAp7K7FA9LP4ppThpo5BQURB32d3S8KA60BD4rr/JKYOs/LBx
4fTNZxbK1bsc+5R+fPb+eXXvJRu09tH27YRuAjF4dbLXk5pfRd+dwqTu7nM/cPe6TMSACpKpLGkb
4oWAYDpcomO4FeT53dzVd8iG6/4S5x3m+PU3iq5ciUNgZbi3rMoNq8J9ROJmpZ7Oj7MRhZD6PgrL
kuG7V851R5ZmGIpFXWcTmNSlZnY3HNNUX2o/c+XP2a+S0hFXJECA0dCoT6XT7CjDca7L5A4njiW9
ykgibamNTSO/IbkLFdwOmmdN2pEXTKJNaHC2i+7gVQ5jSvg3iC52UCOLc5zEq/hR6MwBskgyPxyj
oVsIs92Kyo12mOwqXgJOcPFCpJWDhayyDvlczowJ9fUx+ZN8f6+UzPa6tWlNwazwWk6obx3Z9Ss9
iCQfDczKaK/cM0v1/k0Ncx27XKhrZiTPXCheMry1mEQFoSP5vHse0ZVojMgOoHXI/snUoqLPfbvm
VBlKZcNYqwhsWCgNSXgAQTrTT/Ngi4KZPpA10x4uKYEfDZVeecV5G+nlWeEGB5MxhALpOB+eJJ2p
kn/3R1CVaiPMHdUoZxX4jP/YZdWcjCzqEOfb6Q0dnFK5N8yv7h5rZCw9hfdxOApo+n7OHpVB5yCv
03Dxa9wTxcqmUEQsKrrtD5/doKauIos3fJTyInGcjXHZDBY3qJzaR8tP8cQmDf9APVaCwkiabtpP
nplLdPRncfZSLW7jN4pNcvWRJYN5kADs9KfI7ayV+byAAA8N8VpNgO5hpHU0TAiX+9B+ClEKO8O3
jmTSrzEfjl71CFsEDM6lfJs8hHW5AteAFFOp5vANZIPRpBZhMUIDQX8KPzudIhVT8NXWXe8ntu/Q
oZM77H1zzPY7EnEPYkLHUv1cq1hePViviZxnuuFm7SOTGARiUebDaTg3b0iW6i+5s+Rf/Ga8roJq
LHN2Hhou2FcdXt9xz19tWDKrH7jAFsf3XleaGZ3YupMLuFBy/symTHXYAS1eJkqnQtYy5fHljrbo
mOYuS9izKZhSjbnhTQGTWtxp1f4HReCMgWd1XeYYuAGoVzUdCoIObkfJgws6bS+eWUR8Fxqh/bSw
kyG+96sm7PcdDaEVrPwwg8z1iZofahDt9AmB0y/PUG0ew4MgqRa+JSRfuHhfOZN4VLOKg4vc1ayO
hocjjX9Oqfvtlxftw0MKvggBc9hKv2NXB21dTQ9OvWWkpKuwTALd9VDYjfngDawq8VtzrxRJnmlg
f57Gx9euXwqLloqDqRdZBq8JvJr2FAxWDmPDlvDimTepFjeiv9eWlaCKhexlkF7KciYnKnUo5fz0
LRR7iSqtrvYH9YBBiVpzOMmFdSwQ6fyCBRaWiEMnGwHOeSlBTlF7Oi4BT+mubt6cE0KXMB9sGAo2
Mm/SsPGijBO//lzPdmhpI299vF1wJd2WMI1ozg3KP8nHwpYcbGf8aTca8d3V5Kf6b9rOvuYx5jHF
3pJg+JslcgYT9wokd0XfRFjK35H8VRMo8wUHgGv60Knr1N7iyH02D+Lnd9MvYqhlOt7ZEI1nu7wZ
/lNN01Unr1v2dm5AHiWlx+In0tMdQBlC4lNVysZ/4wThcaipr+TNaaclsj5tz/PH3FfxDWbnDLm0
J/2Z2aG956D5z3OoE1dAt2ECSSgZutk1fDhGkUnEjp3sEWdfKsINqCj7HE/eEBYSbx3wgQOzE1yg
rfmZi9W0/iNTRdYdgynJeN7yemz+HYAYZ3ZbLvrWLBpHfCAerdhJb6up2/wPkftSt8qd5gFo2YPc
yLy7rmCVi9atq+cPcTEdhRe+oCLlNhQllD/BV1zYxQkbIIzOs3XzvNLrxkA0yWxjACocb+z0BHCq
AVbwVKejsKIZYkd2IgEOmuruhLhQFI/uK9/YznuaxxVIK42HNjljlxO0mXrqcbWMWhITQReHIxHt
knwzXNOUYE56T6EBjni6weExgTyQ+Bm/jZIwVmaJHDWMrrvK1GZXIz0ZXsGSXPDM4XkH5KqOoAWM
Afe/bdZO2aBOJjlPg0gF6CoJq3xYioNsg8FOY8PF1id+wv+htZhmL+/ulxdIKtxDO87aw9jJSNsA
FyM/g0pDbDvcbQ5OQfRm4cc1QoJYogLaz5tHtoEQzXvEEQNl9jpZIaYKyZY3oJLyDAKU2guLdGOL
FVp4ifExoo7Cc6b7xa8TXss0d1EAgjvixPYmBd2wN2OgE74dhJyFFOsA5WW2YCw5OYpCZbUmC5vM
pcM7dcoZFCmCqOC7FlcSXnzq0jvcz07uV2cOACTNu7WUvngGOKCTo+xwA/8wsbMEis5IApQJcbK6
lVMc5wV63Ql8CRK3toIGbtBUItriO1xIShgnUX2WTDyywr8TjKnU7BA2wjL6s/BxPHOthtvLMIl2
znSnlwDXuHBAu7eH72Hvdle7chlS9XQz5rt5jBob1SXS9gb1bRSIOY4srlKNF2iVDLqyWruDpRek
PSSZcKf2woW8GzCngQNGf5iq8K798LvoqT0JyjacdhKvcI6V4zD5w/fCIQyQM7B4zowUpSYJPs8R
WRVWBOtUiNCfLH8Onhz6Xjelb/yqSGXfSoU4oMhd3GD2IFbkA7wU/jBao+NdR401fD/IriXE4dLk
EQgjmervlA8BSe5lIIw4eFoqkqvz1R/hHyBuUdcZE9GCHbraUtwGCFJPW9RcEEuxkmAQiKUKAqg5
c0f9ZiDR9Dg8XX0po1P8ErGDIhOA2x3mP7DUiQ3zpDaHyFxGi17YvFcLNPw7Jyc/CQnzKKbIOewC
vUpsyTqGv7BPdRvPyyFMalMfv4xcL63FwDPHbiTQIIezmjG203v6HNDHYlXyHQL1ZVl8zo9QKLqo
6brnDJVhSfLa22wTVSxcwHJkggAqXSRCXBgMweXrrUm7kZepahfdi33XrtIm8sO8kZie1cgMlvsq
GkcJ+jDg1wbc1OswmS+XubxOrnLmc22sLPYSzUKZu9Dp/le7Eq/MgsDKP8QK+PcLjlvrMvrDetuK
Rpv1vhU6/64W0+EDvzG095OnO3fBI2Uf8wZLjA0GwVlzeP5qShejkumGVNiY4JXzzJtF95XrjPaH
qcl3BC795umTsrGs9xWD3F6Qwecdzd8YfljdD9uI0jqDgefwX32BtnnT3IIqeltfzsF+reTc//qz
SOCVSYM977D1tcFQektwBYJT0aD0xr0JQe3ry0I9lyjJUZI4jYHzc4z6Ris1ZTVaBLDThs5z/WnR
Nwe9T3K7EZPSlXv7Awlh+r7mRxtDSYYjgz9Yfy2z4NLudpJn7QK9A17dgDiZ+X72qcm4Zlf7CIOn
rPYvCym2iiq/reR/9o5MezYsY5cJCvVNHLtvsU0t8sWKKi50+ke0r1EtF5bocVfu034P+VUvPmVu
TUXSRJzw8U0j3P5BqxmmKI5jVFJe5fI0Cc7gl08YFzvF9voyNGxqpC+XSkRKBq89JYQf7ylyhQhU
cJaRcItc3uCAXWjrtVIsgNOrsUj4Yae92QWcE1rsONpN0bCPmm4Bepe2ANCaJC+HACGVgnj/zgeI
3SOvaI8AGFuqiaHut++EFY/flQj0CyM1PJtHeBlbbz4F2F3RN4hMIAlEHM8HFYQGAn8A+klxxQmP
gNcN8mbQpflsGpRqdeqljATzcfvCn1UOWdqFHcN8laNntz1cCEyG3KkWlHpvJQWRiYK4Y5Z2rLfJ
U+Drpx4CISUE/KxfSLkxs4metXLutB/xjIStQOHtcy8KedZGm7qAUBYOnsNTp4pv45bmG4EfRMxz
OCxDbtBO1IUyBPZFyPSD6mtxMkEWC1dxeTezkwsvhJnuk9AONyl99WGAAlcTZM59Kh7MMSCKO327
6fqo37EYo8rmP1uu2u1zIjWq7MLluFRNnMwcY/FVwtO18/ht7azNPtScbhmnRff8yeBMg6iGQDm+
CfDC+TX7OmLeMOzY05jh5K1sbtiupicphl+bLEnNk+5EAHLs1AuFwFgDeLhliVd0GrTUblCerZAE
p1ECd51ZC8LoUcE9feGD63KerdG/9xFn8xuFx3wpmWu7mWPWFOXr3IpdH4+3dk2SygeRmTJdco8a
MH5fMMxX0uQSoTLJBku29NX59jb8K8LIKynsqTElKY5PeOher9VuYv6Vxu4Qq13BcGv8thi+ygvq
Wsm50v+3RKbI/4bPRRJeUgpdYMLBXXHwrgDemj3XnT5R3lH2RMqqf8pFwZA2PQatzaAkuJ1BqLlh
b1zQWc4d4mEcFJX6yLDTM197FtjPnLxbN95i+bEcndj7QqKdqhOTOvCTCHqtixrg+lXE+V9fvUAx
mJIRLMllXeY8HERoMsIr7ZBWc8AbnF7837rpTirm3DreT43dvnby9EIh/4cIH/2Wxi6V7QI5CAVO
IOALNXS1LYWvK7k9GmCcVESIIgDIrzgsoIkEjy7leW3Vhr4bw4F6eB/IJwzJJkgkuM9kJ/Qyl6if
EIR6g04BTsIh30Kru+gKHXYwEiKLrNYtYZPu6koMWh1/ZQr5OW0eg0KrmYtLuEh+9oQMSeCklue7
+1Li/87uMch9iK9TLoe/523LszpajBBuuJb0daER/aJ9hIlB9At+sKZQUhule4JV/i7f/wUKMI+X
Av6QcVb7jLU89nVa7n48bNoMBwhh3P+Cj7/X+bzakIUPg7/wvONUSyN8CB/VAKszfxgfeZ9jcmIs
KKcO0CCKbGyXgK0ZkiUDB66m/5C2oqFx8y4bfl9E2+2ZI1JlaO5mUGVJ2T/Us/fgvwg0yMag2b5v
dmhhg75guP3XA67DZJtARDG1D/+N0DLJTQlDv/JrKaiPgerAa8seMFRvwL+RrCHrqCoAGFi11zTi
FkOi47k076P41uZ2GiMjXaxPI2ofVlwoIIhbeiq/P5nVex+9Gcm/6lfWFC5c3Pl2MF0Vk2HjLnPL
w+i21w57ajAXfY3mjwGEOSyHczAzA7PdKfY0ZK2ax9Rp8dYkCZdl/zALliAe31zB/74+PfM6a+kc
8fzTEHsgRaqpLax9NguOR4XwsOgnGC13THdx5YJVLgj2dFEXBFvzoWWpXWU5Jc3Zdbc84YjO7kBC
33D9DfP0a/gKiv0+9H0vTgClldXR03X+mRSufn7wsxgicDcoMrTOz6EyBJjzlhIvtBiMdC2P1Mcx
HdrRckS0MLfUSTT6CdXukfUipDBWwZQGPmCATJgqMJqeD8O2atTG92qtNeopKIHTOqaK9uRBBgKf
ylHDgrES+19xaaNfVEGysEyrEnQNBrNqt8hsTJ0EiC998q1ozz2pBUTvdr4XfMlx5/Wh03uwzfPL
DOmxnPlonYKyguu38yIZnhgugWT8PTNZ/nyUzdzte21LuRSOMflnUltAPp67LZbFJTZP5uhY7+h7
OzmkQ5yDeM0aGD9desQvtZE/UdpFaE5Dh6LbBtxRaLeKGn6jf8BqdjT9UEHST+//2jsvGzaYrsIF
qi1L+uUUO88XUhu9gHf4Sqp3A9yfA0UGJMW6nimCnuf/Oafs7/AgJboBpfKA2sOHnHykxnpm9M68
zlCU4i9lrniVL/rneeqLpFKiV1BgGfkHpr+QQRQJIC0a6TgW/u7burvA/28vGjJzGLUreW0bQs2p
23iRLepXE4dKWTAF9rz1QZhRcj6jDFC8xxhWloY2tNg1KvnMhvnZKZXX7fBAtD8jyAwbwG8CeizH
cnZ/mpNkaHa4TUSo5lxcS+b+tH+TfKZb/ptdG/BCVSKFtp2SEylKdd0J7HO7D0vE1JVornwn9O3R
ppVIOhQSllswEidONwZ19g0bLFglZQmYSzRqRyubyB/3rN7nEqlgojsCcGXRpx9JZ2UTiryRFRUX
n713SdaGeE0o7DJAXiRJeDzi1lNZrvmGlqjAirgKTTCeq+fE2TV42PCHX98DAzAIk1j5jp+kG9C8
A4sSsr49b85vMmz2G7w4nkbs1OoDXMDp2dryrC+ZYnsQZ2TAqLHDshDWLr55I3cgxWgglteLLWZA
DMSq13LtMRQp2zuXlaB+RN8QrQX2ff19UkTkNssTrx47Ax1FBqbi4pQa6/DjVAMzXLFk16fSIhvW
xXOmkfTcf2YVkFm1mAgcdC06PTRq7aplKi4KVsklHpQBFqKz9AuQoiX+l1wAWzrONCRybqgWqn7h
V8OB/016T9PSIQpbZPlFBi+tfovilWg2f79ZePOyHw1eN7tcZqbf/khrsF6U5IUMhvobooqML0Xs
PYKISkyg3ACaPOX+YGbyM5pno2L0OBgKgmVzbBsOdTzMM8s5kiU/KB79gbEjUKcnItFPgranTpvO
LrcTJfZTlcfUfZllPCKY7e9eZwUppbQtgjmloBx6lsYpmgycxhyT7HUZwgGhMnCfu6jGWnZ8GxEy
LhYDFA7/7B08icGpWPnwO9Br2IesRR+jmv1irY0lrljLFA1ONU1wt9fQ44gQ7C8EvBtKVG1LB+Sv
g5C/7a4tFHs5ZrlFgs2X0OKL/kv3k8lxmDVPl0+IjNtiGxIeMqNQvjXiCTg61a1t6/xaGZ9i4jj/
GRieeQ2WwxeSl3aG3JdSETM49WX+4j0eTOi+da2We4VY6MuEyeg5Agwb5orD2Ytynpr2bovXcNU5
xgN3j22/tSpc1wzVGlq9LdCjYLuFJjsizep4t+3PRZGvmygAvM9WmWjXVtVNI0il61CKoJwcGHsc
G4so/fNZR/MjSO52oZQM8pa+hxg1tN0uG0xykTsfi5QZU1uDiBxxPD95NrDTq3EPgKMEzZ+1qKUz
74Gf1pHD5I2E7W47gPvilMg6amoN4Ob0r99yOzNohegUN42DewRLWqSjiS+5br3VOUySMkWqu8kb
MdKNuYIUpaKFfJjXNGXX2VSyzAAFfmbcIbC5qsTHMH4eps386kFBlbHu0wwmXR8J1UfwTZKNWw6Y
8t5oIoE5UCo+iB1ryd8Jj14sgD2cUG2on2LiaQQSfxdvxjiewmaSAPZFtIQ4xx6BadmsCSoBoVcn
Ds0oxnadEXruzIAX/dkfwWYyaMx/JCP1DGYaqTrkJeVE526VF9kZfO/3AD3VhAaqCSs1008X2z9J
cJE6LNTT7fNontpcybA/IMgb0xccrvLO6Kz2g2krEmEQbfpZy0Sskho7Tun4D73y2vQfLKoXzwlA
vBph+S/kwaSFPzwRc3X7TI/62jmeBke/MtNVZsyfKb/HonxgkEcjMowG+6JPOI5oQbEHUHQaGScg
BpzQbGZyvYuJlfCxicll0aEy11KIfqyyb8dn0aUqvZDEhzyEtZJU+b25mFYoZ46ObnRNFQaV6spU
HgCeutuKbZoDoT4tUDe1cEoTnA8Hg+DDbv5HKTQ/26TkiS96TcsY+WkKwjkq78+wg3lqP7m6+DAG
waxwQ0l/kPR+QA9Z0Yq1hDT1dFQuyunm55jcV4hSNtB6jBQKGs3d4iZpwgGFJ8TQnTvoPSBOyFDC
CQtvgVErmZFYJY3RIz3OQGWrdaW1kqzgy3ngzNiojNFbywxD52pIDeD61OXh4o+D/QbWeVmkFI/U
N6NWh5oitbYjaGErukwKtDJFUbH+sTnIQOwRC/BaAjLdflYpucCAlv0Jz09hzR0xjVlWk98a5Nwb
ZSD9TKuqi5/rYwl7Ee0kXvO7IF1n20d3WEvFY4ErePTJseKf/D5fARM71yRCfIEnQmHB72jFz64B
nzvMvHgE6bbuS2Hjtg5GBpukjBdG/FG3juvow/usFIAjIwzwYanQ9hT3ADcyhe9+KLOmsKN3xsUa
M9eWRQSgl2KjSQJzhV5yZFsipBuNjQYJpAKUmI/ulx2yRzgzp87ty9dkxih1MEJasCqpS3ExPlYU
EYvTEY6phvzHFRG3xhVHT7XcJK73QO0ZoVBv6Dsvk+H4NArSdQyeKi7YQh6MMSgoMvkJ8yzr2G3P
OKPGAtPU2aR0j0jhOmDi6sHdfCJ0IpBPlk8CLEm6i3iCFRh0O0GYHEoDsg8OA3j/mhUvXvf892on
ec7yLwhrN1tRFxyRmvMj1zfe7jbDJLqOCPp0BJmxLKoXwM168uT4hrDONgvTCG1kpFRQhZdm+eBU
iIUYaqAyOI6O2D2rU3QsYRJER1KBqf4tEUXzpzz+UmiarwoEiD6EQcXtu6qEteVDPSqcdVIlDqTg
i2XkwSU3sZ387Dq628NFuUeZtrLtQ3A1sR0lj3Zt0QxTC5J56ndWy05nJnaCjYUBkLqao8E3G4wu
gRxn9HNNjB5iaf7pOjfxcJ4843FoMhfbXFmtbsgl7tBAmhV6rp/8uVRqiHdZxwcPUGTbmrnEB1nr
xl2hIWyBU1gOyvlSazRzeEQkEdAT1GAWKnvE0Mw9LQaxxcy7zltyFEYZoZ1ZkkOzBawovpghbxDY
cpjMtJM4BAMDo1LwZ6hZoEb16G/xIpJa1bhBA/JR4eRPQdPFDyST8s/cs2D+2W5EryyPo4UWoJ5D
CjWhdqhBx+JwE4cdz9TSQ/d5pTq6mzwZZqtqaTULuJeXarc0Vla0cEGfocScLYNS7sm6UQdbsCxd
DjaV8E/xI9h9GeHzeKXY995BAeliaozF1U3PMiw3fVg0RXTohqTG8Tf5OROOe029bb2CO4k1pNq4
eGN/GCg2OQK6/dXez5GljAvjPEZDOWu5v86pvmWtRVspjnNrg58Lr/JeXGwwdfoMEai7xKru36X5
wSaXNTIsmvlDaSwJ2qDq1LifG7d3ZOy60AS+QEQG39vPcwttGfgqBfVUr5eC4pG++LehnIFx2sin
h2wlrhc4gjV7/9WR0BvoZqY54o34I9GwZatvPmD0zpJHul7XbtfL4/RdSTc5fB47Gu8cnNOGbEpa
JWZBN0HUWFBzQtR7e9rcaRGngnWWY361hP8S6+GFa1DwK97oSK0A5dgvE6/vVkUeNUPnM6NfT6qg
oY7nF7zF9h2lfmeBs/Oec52LB9Ed2MsaMIo8+Zz630OYDDAES1S6wwpIxu+OcWyyOYYIOCDpWuby
Gl3IHDijwXP5i0bf3rVlPpmmVGmgeNlCGDU5vxJjjdSA0LgVFHk8QysbyccUSEgt92VCcpRQ0XUc
k3vF5RM0N8a1BWyWBJehPl2it9n3zX+zC7F6xxAZHePuC4dkIMg+7RWWMpSZie81GAHIHuHhWso5
3DH8dgPONvfSEuuzkGxq79NbIW6a/xu9mrOnrmDL+P/uw29+okb2GyyoJGEezDVu/F3wqeI/E6eS
vc+9fgB8gtr8Jg9Z3tNBvo5zOjE3OZmZJ/CwMxkggWRcI7c90cUcxQsG/HsKPMlHDb0+NH/hDURT
Gq6qa2w32EbbR2vEz+l8fvVHDpDIlrC2qYwn8Pek8ZIA2H7lyBXdKqrSLT/Nurd1iaxePSvLfeM3
DsdYxHTvePCa2MESkPMLOtdLIsHHVNWgxfsCoZf6O+5qVjnpwLp/OuhRA0nRKO8UnSnpEFw4TG47
pWz4YMCqvX2NvNrR5g2z8SEaYxM1z+o5vbfqFiQK0NJOj9iTl1HIqforYZ2XJNPi6o47EhaETdMG
xdr/NOhF/cuz4lf2C/YYlmUEjpx0Q/7mMB4stoV9w+7zE6D4vuGIlW/QRzkaYqrIUFc1i7ZDDJ7v
fuPGdRdGNACiQ20GCbe0RVM86eQ6IEYxkMMG3zrhzbiP83d0wW+xlSL1ZSkJskGjMHhyYAVorYZ/
dgRs10WTIwIe2cKtsmpHGeCLjBHCeJQ2fnL/AILqff8pHliV5yDEgfzFnQpS9JM0TNJo/b3VVCqf
/yhzSzGtLKHyxN4kEhCS68ouW3mDcZSg4j6hrjrKPYci2OIDhRon3GORbGVRv2xWeMRsds+iG/p9
Je3ac1K6XnaiSBbycMAOQcQ7uS/jVuziOY6Z5wG767QrEjEtm9jODK4zXPptSymaaN3bTKG4aZuw
qc4qaV4mIlKY+Gs/vKByaVt72kO/YFb8lSt3/pQ7+5Z/CHI71nXK2EdNkXA036ha/10j73pRStDM
FEsF0W827Rr9HZa6TXoxlHNrAeBeX6Nfu4ilY/8Rgptvyq46Kjd5QNbG4w2ySWimQ39CT8c4ttga
myOcU0SFQOZ2wg47CA74MBdhnEUpFyaTnts31M43/fpAqnp34L8Vf1q445OhWQkwpqXZ0vZslvYL
taEGqprvlz4pusp6gRpmGE58nnGUsRyZdaSJsRwhTyJswQLVSWtaUjVIXCIxNHUDoSS+rUJWSvVJ
BRYIcgRnIv33Dc5pQb0ywZifTG9EiNZZInDLbnnk0JCSAnRrByrOX6y+8/JfrT998mXBhluvdg3S
WnEGnnVNPzFvDasCAVhO5fTA7SdjiaGSL7Xn3SZQIx9WPFiekHNe/spTg6SAls1vFpxTHn/4N6S7
OSyP1XPlsU2vLBs/zvTgKRw4xzYVcRc70yxV8jsijwd9NOw7MpsUQpZ0NfN0M4GAoYkZ9uVNLb3z
6tILNsXkWvK1FGnSKilRYND82C8ET3E9h48gK0SM6xqmjZ1U6LEHl0+GAQpSsRCuCeLIQgfYpWRE
qgrheTmxDpSfQPxZcadFkPqVbkBU8qIEIW97/IcxsNm94vkRSU6GjSWSi7r6Qm60Ek67IqH+L1EZ
Kj88z5OoXsHZVDwxEvozHLryTxS/5z8dsWCvv1fejg9UvTEXRPjNfbJC9gNjgmHg2vUj//OHE4BJ
uhuuek5wdHYeOgyZQiJ1Y0WW6EMZLXPkjuP44pYQD3pTTOcsDPH8+azOKUfrrw4F/3drQhrKQEJ4
90/URAICFiFj1FzFd4qaXKMiArbcVPsH3D2oAegki4qGuhRqkm8aHULrQO0mX4DHVyhlZw2C8qzK
VdJ3WAK873Lg9/No0lBlppKOhhzyEHoW4nxA5ZunXJazeRRbN/BbzUrsjiiW8kyxZn8huU/SsAj0
IYRvVjk9vjzIGLDXTm64IpOqUOPv5LH5o+r7Xv2lBm7pheKUBSvi0QrOQOwnLOUpJV5eUCyo0U7h
WEPdjjmlydo3MqQc1PyTb+1ZTqdavivi+YoIy+wimOH212RWmEFF0uGk6lw1p+Ky2MwKtDHWXAX6
80kHFv899EoGUhttx7+h/qboPyIvES93BoVJ0xc4EkUUKOhu4UOGxTI0JJmpmLLGz0dEEDAQZ6Wf
LTJB3KekOGCaPgvqaFxSRZvPAUrfxScs2wIHK5j1sKWhoDEKpMV79YHXAxyjBb2vLVuX7rTPas14
2acNxyfRdiGfONunP+dMLTMb4njr0KzOIYHx7efisb0NrKnfV/la+0dlUqDA9tOUicxlPkj30uMH
bpfqVP1inJvqdJe6XxrzhmlP19Azy+RXSY4jW8JCrjKi/BMNhnXa4AW4cXusmjqQB+PAx7qTiyvc
ecRndd8TJay1R10UJGk+Bel4zN1yAdu9xRj/qoyeJEN6ncSbI1CVPwae+wBv6MYgp7hfWARbpSD0
dFvRQxmygLUX2BPyy86valHteHHzpvetXDPsVLosP7HL7FK3ujbV2cm/KkMml/K1Qgk3+h8wOFTe
6YiLYrgV4AmdWn1yUSZ0Xwgq2F+Vyh0A2QuIK7iu4CFVuQnM3l8Vq0nYpXEjOvR19QBKKS+79t1B
VwaUF3TBqKVNRr+bdJSvRC8XAQiEgUFazXA0gDbp0V2Bh1uy0jhRGXaKAypIkdMxv/E0n4KlorVx
fCmgajA4oaiUarzVb7hY7jhidD3NCXRbVnn/Ersc83xeznKqsnkxXcj9oqF8K5PjqBx6f7BAEf7n
xQE1dRtLa02bA4cms9EORXm6z41Grc/rm0zwVgT00MQLLf5nWuOk3vEkjLkvxqbqeS8nh9fRukcs
HtarALiYZkpJZD/yTxbKzwQi4QxgO2EhVR/3yx4jXkqr2xdHODQd2Mq0KYUMgi3VcjSdRpTZAwnZ
Bg71CFwwWh5sTGOdxLsDcJrGty6cPwaihLfaF6jNYN1VxTN3jG7DciOdB5Mx/FCdeTZspN7ZKByz
F86UH5wrO2vweeVNqYQDh3H1GAuxtDSULHkCQlm4SHAxGLF2BnJKcW0+sInaXq0tE6H7qScfnuta
GEPB55m34+Euaq/6CR5G1NmfyJzB9OkSyC7Yzdl8xBTZ/bpixy0n2G59lW/2TBAkbFKbAt4EgBiF
VUvqI1UeUYdR1/M45Ja4H+77qdFNmetSzVo1nmauQJZzQ1oVSvHI6R65DEsorYBhUClbdTm8IOLu
9cP01AnzIJbG1e8MGPxveIptFHO7AaSM585mF0YYGEc2oVvedT8z2L/f2P6OIlxZc8iD2sg0IDQ7
Uw0ySB1rIyQXgAKRC3pM8lJq691iTXcE73IKbsYvqm0dkxnDgT6JpL/29+Wzf6TK7RI2P7PsA/I9
PHKIcBmMyEVXR8ToQu90VHOpvRi7IXbOPC/AZetlXUgfEOgd6UYcqWMmjbAlaBwfQUYpOrBJMx5K
ssMX+0CzY4RwZOP5FWPxJEXcSvrYEH/MrIoWk3NXJQcg3QWX6P+X8LSYIHbUUo728tgsAph0XBoD
LR0NidGa9WSX1Npb4nXhouZp0LfxiTXW/mU5GsAUFwW2CdIZ15xV0XSq6+yZj0pE99merZnCu8j0
sQjpEueoGiLWZzwgPVZlxz4ygI8DPKccbNH9wehItHo/K8WOFR20RXCUZIqC/8jM22sY+RuDLdip
yV7GPAITVVIV1vY0cNE2HAAyOnc6NtdwrNaNWqBwKeDYHIztY1nFGR3nr//ycxhSl7Xm/EA8kuV1
HXG7EOXB0shQKnxddh2NnyjMMV2VclD1TamHDiK70EKSOQZaHXE1ELqyZkfNDKVd7OdUTZn3XUEP
tquijVL8DFxI2G4wMg6jyDp7Ima4/7eJly8JTR5osUc20mMSwHCAioJXVDZPer+dMMK2zQhU6rVu
7ACRFbovUmonfxHNe9dI/ccrbJNRqHVQbX+bWvHtQLo+Z6tMPbOXL5ETx2Ue2c1ACkPIcy8CVjwQ
4hvDx3CGMcATBz46xARq8XaciPRdCmGVfLGprc6oD2shjD05NxkpPoRhB3sb2W2ZleNaB4D5BhxT
2G1U2ua/neHF92nMGsZPa8hYjq0UfhqMauelXyAp6biVKAJ2GqIxhPyPkQs6CIX/RJ/FjxDmpiNE
XwqRQUgEJfzqE/bjaMGcHw5QsopA8RRIYtseBRUDIA+e+YbmPAFnBfAVyooNYQmv3Aq86VGXWT1N
vHbDRs0OzjDlTsNcRfBPDWQZZoWAtk15TgUVes6BhRy9nJ6Ykr+Srq58Y3PEqCBNwqIp0m8cs6YG
3QmAjt/0dd9I7m+i+1qKAGlQyIYN5WeFiiUh/tLLUJu4tq1qNMcW6a2Sw+uOLGSJNzXgL8uZ9nxF
EsAPWMxI9hhWaMgYNU4j1RWH8zhooS0C1/2Q8cclAyK+4iUl7zXvDT9fgM4k6w4OBQP/o0Omk7AC
6uYSrE+9bXVzcCsTjnCkfD4bR7wUvxNH+BrmHC2o6+/6J3M7P7yc7KGfibFZsRfDof9SAl2KeZg5
P99eC4YoO/8YxSqfK8ee8I9EfZ1DcPdLLNKAEA1/in+NzsJFcw5hosowuy7TsaD7arYSmGMw5UVv
vReKgvKG18fAVOvPNgpx253nTB9ZYZ3Iaa6AOfml695Ea41FdADsPBu76fAjjx7jmFzVT4vse8ZN
nNnm3XuKZ8S7l2gq2XODbXoEOXxoalp5KVbGCIr3A8GJEOvaOSbgO+Es5vuUKzflxkfE8xgybWgj
is+QhDnYeGIaxRPlrZV+sZCct0miMg81QXdQwOEjWQ5nJBKuW74dG3FPDdH6zuTMf07UJ0nzGgof
a1+wxa7SnS5+JArukJZKVtUMDhhAdECXOPgQ/KQuNL3hFl0BgSH7p6Jx79w+EqwOHicTn/5T8JTt
I/AifkRBV00HoWTJB4qdyViqbsz4LkjkEnLr7bzn9EgVvUxRZQ5zUtY2hmGlMH4nOTf+NEekQj9a
1WTvxIbEEKKFOYDVnDYOhWBDfrOgToN9lrgV4K7di2xrjRaETkAo7+RjpEjCqZqtTDbJE5UYfFCd
RoMoBLolXuiEznsQ/dY8A98cCpuJbsHvNCjSXD7zq9Fyd4h/F1etAxCKM3apdzRYzZlfRlZtHTye
3aN6onw3dv6aCi8wXTWc0HGnyrmY3hJgVpWO3pdVmGEWHSujJc8c6Kcghfm4mgMoed1TWsgTQDTA
p3p0GneUYpsthfV+bmMmxptQY7QjOZ+l5sfV7d3RLN3WeGqbaLTlwlCtnmyldq5Miito9Nc1ZZL+
NlmVmXk8EI1BLonZ7brIjQrShv+ufQgf7/HAbXxfbMLabPSv2mhXKfitdI+yaz9XNebSjiJpCAaX
AElqmli0V7MTdRlocTYHb/28/ptgFVhybZ+Kd1lA2sNfgFfjBa0RDV5RRYoWJS7KBP5isXdlLlm6
jyQEET/8XGipdxy8b6000Cj2OoHdoD07S3DaWf8TnJbsux2FMNv9Qk0TF2iNO10tbWt1GmKD6aYm
nX7lT1udljN8xfaFL1IZhYmRirEusFjCVxtoch9D6LX4ZS/+MC0zmlIz64IWj/+fOhw9CnNoilLD
zggzt6djxq60oauiWjXWDst4oYMRdra0bBfPBC3otwrF+m05iFOcBdkXx+zReTWd1t5ElwHawQmU
FQX97QohuAUMcT6ydrK1Mr6k3P1hYrX/3jpTHf/RviYXCQMZ9h+8331cZoktnqj9SkQCriDIisuq
aafzYNFJ9Zr9nDJCpaa3AOqgJepP0q2e7XvLSCPZZ2Zt9Rcfk4mNX/XLTB3NT3iIkhT1TsIMNYDM
k5W9oOriBpQCaHLHv92CAgPqovHcY0czgYgqCqt5Z50jOMNd5s8gDTL/Qar4L42apdjshZwBa97x
qz49pw7E/Zgs8yyPzqwbx40pCBxRW+4gSJeFOo2zrbD+qsVDWO6untRVfYH1ujrQ5BwMXR5TipQY
GYCNSqdz8sjKqyL0e7M5U3wjnsQZRhCELEII1Bm8Fhi0KkSkjhKAWTsdzJrBIur8TB4TkohMZi4P
/dZZF0u5KacM/EdLu2GtnhXd+59/+aWuwtF5MNszaNyfXiyvviSBu/r+g1o6aiQiw+xV/KDdEO7J
XXIMXh9/Kw2QbVKI3k9Z4blLPXKQ2y8N/9OKQXxTU6tXFXAwQB+60SlzXmkxxG0JUAQVeqW1sbCO
qVBbM+XizFBZvA8O5dI9cifYO4wEQEgwYw35r2uauA2HL1XdQWJEeq8QUXJ1kcWYNaFqssqR4qS8
pSMYaEl5qgXaOy1mcoq2KL/kxMwfBb7Tx+wZpSlNQgAja2nk/FFyS6dn4dfqPl1ICTUC5y8CB90C
eIMzB4sHjAzNNaQPR5NlHzFzfClim9Om2+9C4Xdk90Mbj0pD0MheW+zn0X8Fcui2ysOGf2RQsH3r
ydGsqQwZdSA//qvtsrVCIvz6f/2WOKLKGE+z6gBmeCEDISenDecaAr1D1a7l078OrBECT853N1sY
BS2aH3AGDchsc5KQCRfO5adC19JDyujdtUOxbmGlEcHQFbbOKKhFa/rHFUkRoGcrEyBbZ1+oDx7j
p8nB0SH4P1GHwb3jYzRBO+qr9Ul4wve8yAIzsHopNMXpESWev1evrf4P5TSP/muB8I07vsbERmmo
sAJrlUVUZXC8Cxu73pT3mWt2TR1nbQppEWEidi8lO/Tk0OAtxJoCLE5sjELuFEnP+eYxVXzJQ2d5
+7ZxB7sqLD/fOpGQajLI9HEtLtu5G4f3UdazAhUNBKkh9m4py/mnUW8nlT1E/CCtNV8CWmDvIMKN
PSiw9SB208t6Oia2hjkceGynr0ppCI4xieFCVgv556SAAvqmlDL8eKUKRgOogfoVh/e41tH22sMi
BL0wa8tiQ6/tKybHuC1obleSqy7DzS9TOd/N41A/RyaQf4eYZj3gG+PAfDGO6JvFSUBfXaylp7oJ
Bj8JDUTOPud52B0ztAamS/Jclce/GjR6JX9BP7yiPYO7zUVeoLBZCmKMHqQmJ/5HL5IKCM+M0ciN
35RHFvmRYC/PYYPL1u9BjX3rl8z5EPqg/MkR5/MrwblwCeSJVB/oka8Q7KgkgcGR66fgaJga5ME7
kUqKKlSbgRMoLdDq/YrHJyZ4t3phWAhTYo8zCAMw18yJ/tg7HZZKEH3+KqvThuajA5PvLjNnBp4h
PLEApiVAd+cDmp1NRcWiZhAZrAb/aeX0gkdL+kqkVin2QREFVmI2Xnh5MqhUk/VbE34xG+TuEwfa
RX/G5BuuuYyRGctcOBHgkZu8vkZlyaQ3GdEeBTrKovZAjEjhkkVb7v1VpsrbjzH5sxelRevRsk4c
wCHhai91BuziYAjkmjO5JaN6YgW+2t/g0/xUKT2npX3mqzVItvoespPTyKAQNpY70RVyAMB2gsg8
AT9OC1tV1KFfMoIpyEi0Uv5Bvd7AITHWNBAaVFRqKWfg2SNtQaH0l6SqLlvyl3h0MBqkuQAp8rxd
4DB+G+MmwIa/Ht1px8s7KTO/wj4mbm9U0O1DHqoANG8PPt3dmZqeEni4ed6+x4lnYOeTci3Yve9G
Qt/uI6Hp+tnIov/NlX/c1BJKL+sMV8oFh+LfNTvPnO2UgsIi/10UVKyExQtH5AkKk0ENDPUHocdp
OQXiOrW/wkyUXZDk1NAZrYubHQxjCc/l+gbj17Etzbtt85RvjrYfXwHmD0xyNclhaiQesa3EbXwZ
UlKthSs6iBZ98PHMgIUx1VFvIlnH/I6660FnAx9VberC5Xyi7vjmQ8wLm52IkDStwJw6YRyB8Dyk
KzHh9TsI1yi/bN7VXfo1oRjqXwBb2HvniAgENNmE4Wt1Yq3JblB2i0eCAP1Vo8VNiu9grVPSZLvR
ydCDexNEPS5zxeID96ytXc9sOM8DzjNuCHa2sLYd+0p7MuswlS072yFYiR8e0FFlUH9m/YSmWs/b
f+Ty1Rzc0FhRuRycIfmq2mZByuA1hOs1JAaZ1UM/mTSKHGFtKgEDzDWx2wfn7P6Mz08flNHP6SlV
npG0lDPAKP0s1EdgtJ5PUerVYOI8KRENPRR0senHHucwiw1a/XPycKQIMaUq3yxIom39wIUV+jnr
s0Hld2FjrMAJhsNUI2egrB4SdibJMCO1BykjJXgGfly51Zk7BKA6SLqnwm+EpaSDUqBriRJ8nyt2
2bifJ5fthhdhnmMwBMtN5JVPJHVTCQ/A4IF+RrB5mybylt4WBOHEk4Nc/xcoQvU486GgOk7NT4OP
BP/qknYftepTuUmWPQ7YzCFS6pI68G3esaUOdUc66x4fCbNJheeNVOo5crx6EAT44B3n9XUSZpI+
6JknVH/KVd6TpCUDKItJLryTRCb58bQsRkvswUyj2tQWV7pzwAKOgTPKJj+BnnZc/c/K8qWv4suq
kWMAQfOoEQNUExZRmAyA2g2E8/eOSSQT+MIZfz8ZbigmJayGU3EKRuJRyuFnpz/uHURAcAsh+ITF
xgwAiZmdX3dZIa8ZpAVVQAFsHNz8Q6fO2zt788gGCqGRVt1eClu1/gltHuKtuyOP5vgHk33RqfwQ
53EqxDIb/WCsS4hjtvIiLC54wn03Tc/aaL+8hNHOdqDFUr1kA3Ozfo64hZlb2Bv0xBzwdrEM13wi
g9cHk7mHaNAeV0LwRnPNVYkdKkOVRQSsgKbP84Om0ojtyEg8kagDmxcQSAZKHriI18rX5HrIVFOj
NQMy1Aab6MJg7AUxPxu0HMq9LDq7Io+m9sE9hnhnpe4pfgKCNAvpO+o6kmapf4SQwUMfa9aRqF+d
z5DcVLSn9A4NkQOBH/vIXUAROywRP7YEkFxytT3df0v28ezUrimZPryKxZ3TJ5t21Y7vKq7iB1Ju
Nl3wJU4jZ0+s1m/RJVMhCx/d/mU8sHWaI4DvtNUpxqxOF0ViWFQR7O6L0r5evKA87YxqmOE8c0sB
HNo9PFddfWH+3Espi9gUOX4ZqYHiARaa6uheUJIxp/n9/FKAMHO+bisH0q23q1r+2il1dVvX8bfR
SbP7DcN4KWbZSWT1igNQbrVGk6KUZ0w2eF63bcjXgkLxDSpm0G+G6PVFru3dtD4I7/9tqVSfwJKh
iBFv7WJPu2jMXI5tyCq/Tse0YfCCbRD+KtkIG/gn5NYrJjEBRK6kRgUktPC8RuMauNjZn4xRxb4m
nLc6h0DwrYNABcgTdNdhMKOEWZF+vRPPi+TYKg71bCPlOn10A44IpT9DCuAZQXSKUFMI29r9g7vD
J8g9c8Vsza7tH4jKKJAdvyOjqySRJwdfCabNpNH9lcd3uo8eefaZxRxizoZqhGzZECe62lIx4riF
UmK8PHErUmPxXyPENT0cMOLXyRTKo+NzUQTjOEAmVotafvjpR97SsV4cAE03zBHDV85NA7SkpuKB
SHrdAe08Jf4rdzCi9Vn2baOBXUMLnwttW5PEN2WhmpxUBbuA+Ax2Ek2J+JAtijU7thQTmwzbndG1
5MhI62PQx85MknrHDsQlBKZnx4TcE2AJkzKK7OZ5T3slAtklnOwFnLgRRMn4nWuCxScIb+YHbWQ1
lEPiN5jsRiucnFObCxhHyinSwxWtUSaRmzVUc8+vYWc2CmYfBcYXaWwWyKvYHKDdoR5QEMP3E5f9
bOBRNmzR19TGJOtdBL2sB1s/Tv81tGfqEjEIqejOfa9tvBcg+EPR53JUxZP1wDXfkfW0guc2Wqx/
IoV4OIWSHXC2icSLMUnK2OclaHAv9TIWdRTNHnCnzc2vkdUmmyXUnkGQcyHMzCDtIacypaDIeeQh
NzsQsAiogsI/nxUPAklp2x4YefnZIogxElTcYGk1B7G6wRCKMADrhE8ObQq1OcHaU/98w8enCbta
2mezP3VocJpnEPX+d1UN3Zwk3znBhAGJ+uj6JEcfq9r2XhwSzrgf729deLyGcFXB11wnTz2KKhAD
OedmbEI657BNdia3tan4kKjYk7qGyoiWWvcrLTi8FwZ3O3PJ90Z0GGhaVCLDGM4F0OSkyUxCOVgi
6kMYQbi2SKnf9hnIUn+5eUDHG4hA0hW/Hs14Nox1YF+wRHlnVtgg6xjRx+x7AORbrkPUoTiyw1Qr
8eF54ZlH5/heSkDhqD3js72TOmKIFThzfiQpMRXRGaf+Y/fuzbSnZyoLmfpqccRQgWVK8WmAKSpR
D3o5KbfcgmBGc3aaG7cyPcx+ZX/Zw2vQS+hS7Q+3juQtiXwlz2i/AsuSpLC0DAyOQd6szAsIkgvP
CFDOJR4oUAUd/vP4wxHaZkUNyP0IRJYVJ9XFnzWDEj7fdttBePGjg+TlEzxBptM4215/ulZJ/s8W
8UN/wwI7TGj6z2/tijQMgEbP/b0Xk/3u9I/Ct20NqHZ6E+yWzfZchH9oaLmMlkgBM+S8uE/TrUbY
0E17A4gtfNrn629ueZM9YBykDV3NSyG2b6L6PNbmCSdt+r3693uOl1voKxmi8O+R8iuoIcocpLFD
wMlFzIJLziZTmDI0RVvzHz4I4rzU7VwIQkkI9pOIJG0RAaZzXJgsxUSWa/k1CpTYWudX4Yf+CAx/
xlL5Ikp3JDWb5P6ViccIc56U/msm+mVPUpQ4J0Pz7TFXoKXtbWkWcInvnRQynloOd8oN4Rsdoruz
5/CRtNq0LaS9TBQiVi0UFW7u4SD60tV+LVw39qZ9dTdvBcjCJbk8wUBLFhEp6tzkTkfWM2DYquRW
rxOPh7x62ILCJBUsEPdHywmxzX4UXn/SA0kL9GBClnFAyZsAiZk9km+yKHm4p0HZAbDu4RG2KPqN
dtMrHERWmq6tsUHgKn58AX8GkYc0300Dzq6s5vNwMgrx8Qixbjrge/+KGZ0tym+cF3W7Z/y7av0a
IaNQHlmNguKDCvLhCrTirKkBmanU3qRZ1Y6wMtAOrvR+YAWSSAkWDLtDbrRUGOlHnwpHiIm7UKVL
lCG9VBtSrdNOn+eAd6pVhGGR7JDun8KUA8/YuPNaK4IE/bvUJNdHmNPcX+nrWsqWEdP/mXf/YKVi
uBYJwFeBzei91YWS79XSU8e6c4WzQGfGCg785eDR04MVA1kuLgYry4PaTUx0PXirugtcjVIlH5X5
QyUkuecXnGKBoo7VJSKfARkWxKPXAd9X6QCoqpmf8Bi5UK71Onb9HXG1+7SXNrc+CoNjH+a7Qox4
lWLx1N9lmrwvuZntnxhuKTeRDT1B4YThc+HPpQ8d74SjEvtWfXdSiGWFhwsAF4RCIf7UKEGtn6wp
qLiszwNU6yOZ4dNBPZs5rlx5mJZ4w9o8SL45FzivG3jWEhr+tIean4hRwYzS1d/OmFU1ywHXVqoN
NyJED7vgwhJczqgUKrXq17CeE7wSXLC6Xv/mcHlxlhrpu3LL8vtA00l6YLb/AMNgz0Zks/FBMSyV
8THptAWyinkmnqajn7uMUfA1jSadVNxGwMOqa2TVwN/0Ahn4UAXf9s/KWRAZQI3HrGRaD4oE1MgI
jmkQFuMFV6quAtiW3IcA3UeHzDrXA8QTWzUZGAnEkaCcjWDO7gx7LCYXG1paCV0PN02m2mCsu0es
A8oE/1avEPUDTHyguIJv5puzJmOsKy3z8cb14VvWBg7meaA3rIfu5/fE97j6Na1Q1p5g7bgQhbcw
7VszXaT6Wu7d9Jq5MOLsLE5sY3Nsp1/RFpySUsyyVXR0nQV9JLeBu9wUZeKEOst1eG4J32WxPWHL
krIw663vbYKyjiT+mDX1wh+/5taFpFU5yYwJdW2gi3bV6eCfOdcHWZP0y+HY2a3KcHAF5iP/1LuD
q+19qm4pwxriXjhrJ0f64ZYtwWdd3JKp6ca60t/ql8NCtaMfK/sPvOdeCOm519QbGH0hwCLJewvO
iBCPefuFRj6Z6Mb4Gw1UjHiLoSA5Mjz17AfqgeJJCZ/dWgsktc9mdag4d8PNZ9PrwKuStB/hESDA
Tu5sJPdmyF1JkgZH1m94zYqYScI+mwQ5LmylU8bS2o3sDKEDTI4KdvfMPWKnjz6TQb1/Ld+86Irv
F4Rj+r4+LVdj0aP9lEKAeiLhBhDLJgXA00pSACMiULDuamIvsICwJltMoDW/U4IzwdWb0OrSOqbF
f2YPPAJiB2+HW+m/hqqiL21gvdK3nC7Jojk45Af6UUcdAPUt+Q75txoXae7tXRu3W4t6+weiSBnS
ww/rA3R0TXVLGA4B6tMU1h4C1R+2gmO2pIuKzmxZWj28JIOKshiOnB2Oez4hrOGu51n+10zE45I5
P+CG7krenimfNMbZihvvM+0lMqu26kvFcA/M6aDerFXz+PR3fJk++PvQKD7zfRWDHKU8uan1m3AU
Ulub+Z0SRye+YVa3HkUqQPf9+J4f7+mrVBI+XD3oythQx+YL4PFXwv3ueYgTT4aCpCb0vNEWzoGd
1ExjhjrgWyHtlMiN9ns8s/DPMrETYtv97KXmy4V9GWp6z7gy6h6zMJAX985fna3NfKWdfROgkF7H
M1ynpUn2w/H8e0afK9QXFgBtQhoHTRX4PePb+hJfRpWifW/C14am+tLwEfdM54GsubJ/ccTS68o1
3BTtQGrYT0yeeM/iuy+oYu67pUCkTweV3Y+FBZ/OYDB7mHeFpwyLZW1yQFmlefTfA7TPUYG7PED1
kd6Q6H5qG5kTyJPP/9rCCYUEdBQthEKR0ffIyP3QgDhF9KeX2QXZiNgTXURrY+CMUu6nthKqgvKr
BkHoooP/oLPfOcVatqPLBOVA8E434yLkMKbnc0zvAupOqRoKub8xqBY+t4lGIWKqoQtTye1GaEGL
DnCw6M09HNWhg+YF9UdzIqCHvqPgLJj34BmX0mE3fCM8ea57P2D4kc6XfsrjQU2byRccvoomwA4y
AaV+Zrq7Z8Tj7BhGG/KfP1KaUppLuXLc8tGdjHcN8OHPHuq1sJ0lFsK93RF8r8reJBS7sO+yLUpM
v1hX2godqzK+zH4G/pQYEERszYihbWRSMLwHNg9Lu2uJ9XRg0MDfdKbFOj1pP/yve4GbGuFtrVlb
7uWJ0mSdc0nEMHRmdcj0ZDqkXoqlZnK+64FHMB+rzldxy9IWM7ZQ1G63doQaxXCjHgBApMXcsKlo
JH0okQ6Dx2CV+2r0VtydPpUek6+YUI+h4SblEJ7t60TufCEKCqr+rtXm2x1ynpYCZYIawCkCfOOV
jUYbRMb5UpWSz/SX4I/dngTNQLEPYlIhZasxgcoRPilKoME7vq28SrxBfx2QqSmBDdssyikb9f8Z
1hVMEq0YiP1DrwtVV8yE8mm1uGrEJHsChMkDcsDce3d7yupF9pKWKOI7Ut2ImfvRN8wZEk2LIZch
1P1VJF8WOrL9IO5bEZgjilVtXCteZshG0kQTBPD0X8BRTePyB8bEqmVaBFQOuxalSEfI35A5MT0x
wjzbw5SL5/gd0jVn/Asv/sHyvyMQvfnWwYT44jc8b001EKXPIccAqjdtqPux5EaxjPQrf8LAmBsq
j67A9p2fWK5IjWvKL2YEq7DiQ0/IOFQoQoG6JTQyWkIKiYMFDpvQHgR4bB+ZvbjnF9uCFekHavi/
JHI2UK6F5UlXWC65288joT53hL1G0WhRnUqmXOvLo90MnzRv2w3GbteUn+bPt9sFRrqSFEZXWBA7
3U8QJB73s0vc8CzW0kNVtTikXZf0+nqC2M/iRZFfl1766grswJFr+fRKBNwrWjsz57SIkYTHSuf2
+2zjizPaQAIERjydhQzSEERC9KqZjYRo16A4LTdA2JHy7JM29KSPBZfgw+ELyJD2xcuNskqJ7qtz
f1SUepd0kahlttgQzsei1Df+MtLYp3R3iiL1NRfj3VjlhEGo0HgyvNBeNiLFtlOfY9V2no3ySCuz
wOIhmQsD6yCpgcLCJoHdXDhZzkCyV07Okt1n2jjc4tgx7gNKC3zI/nms6DfFw09o/K0kjIBm0llP
Rlv+lo18hwfbNtXZjgYNzPrWhr1r113evxtN4l7rtBblraZ1TutY/3SwQSfHjaUfu4swumLs1wLq
LAjATtKXJKWom4T0x3PXKPzYhNLYH/BxC36fLBUXJS4So7YQGflzQu/U7uVcvn0oSJdsOH3TC+BA
xFTFkrs7aq8hpfuDJvJHOdNPMHudHWjNuOu2PeDSeCY1ZeS7YDFJw6xt4wGvcwnMzKtHN9rzlQ3g
BahszsILYbKQPJz27taRADRAc7HfVu5hJp3mMPEED3SEdvTQUiJajOYUiU6VlETXqliSLzFLtrx8
1n26Bqs4aZgcRu3zTBWHQXtjfo9bFqkNJARbTW+ZF9GKqr580A6Fhdxffm2FB6BSBwoD4coUPffF
AFS/6lKJ9zr3z2gWbq/EWZbZPeylP3it1eQaU6Tw8u2mpWalq0owyv4vRFwyBJe9efFqD2tggnUS
xeAMaq++8NCp/xeyKhC3/tMUJhGYbYTr7M6lZkTv1aU4upi6bGg9vc3g8JGZ6MYZdoAvVJ40l+7R
fRIFfum1z11IzOjTuU7fPUJfuIrQ2DYapn471l4Lnr1mZrqXN6uVFYYYbcsKDRZuIkKHRmKStMOB
+dnN09MHi4ZbHe8ZX/TKPWUIqy7sdiu12d6ODc3PdGnKFieMFiuGorYjhW6GLyYM6O/5B4/pq6rJ
ccsygL73QjOGW29ac2vL1nQytn8tJAIygJUuCEhN+DJW8AbeLp49q/smDodPM0lZGVXTH0VrF2UO
ychYFOywW6Ysk2rK052F85NMLLtv5O7g1qzP2vZSkB8rIj4Ke0LIO+svsuoJ7CCyIwPFj88aEfxD
qRVr4b/491b8qJ/hOyanbs9+ELV6w4AMuu+IaLE3pgy19EoVLbD+LCjyhNZPon+9nlRqyF5kFpsC
RJIpRHsNk60JvUMv413pzIcFfNrlgr97/R1ZqldA5SdefiHBMcx1snJKBVRULcK2YpCFJVeajSaw
hq8pq5iI085+ZEXJzoEiNCD7Pmq9R9NnhDvjri5EUZn9So0FCRnq+XwagRVTGOieAq9zZgGQtLPs
9OGCNj4pdnFI/44gLqPf7SaUx9D9UHl+XYhtssM43Q6Fu/PSD42CT9jMmlmL5Uq89rps3ldSulWJ
/dSn8SWSWFxZljwjplNAAxi8dTmuuQcpZADgUCWNFllLMOY79W34KldQckX/lZSUHgynn58trYn4
qzzd7qZtSDVk26ev3gROrdbCIwHwSgkFRSqf1xDnKMwIZE2WfHGCnGWgrXx/mEAu3Bit6y9rJqDC
KFXwpSuYZBd6f8/pAewNVR3+bznctXMejuXFOZ4NhBO76NZyWuBs/r2M5JP6kv4WUeyyMWbqgb+i
SIUbE/ms8NfLGYfBe68PBQtSTmzIXP1FaxZc4C0kZJVNu2OtwJHomzaxUUcJRk79eluD5mPtCXaQ
mGwyZOz0/wT7/CCkNEhAjXPJQJ/Ay4N3l6fQnWDwEfDFBkDbAD/UtO8mTPERxM0tibex8Zra6Zkp
WkjiBwzJE0hw8u04FjDH+2KPeBpVA0n02zxxnNZdFtbnkrahmWisXGARjFSmuE6US7xe0CE/Ae2j
ctFSIb3UV33VYcKe35zQQGk9eMhs9elZzM4ZDVqs//sjqXxzBQkAtRUZva5Hwa0RR+kEy2VeTbvk
KNcY3P+69wLBB/Do/OvaN9rjb3ATmzXllMleByLGCSyI0f7JqD415lvOiYC4KfrbnZAlCffXUEcR
I1/mX1H6O1gJehWZf+3J6Cw0k5uqgVvRGlAmSrYWgJxtNI+9nXs0JzKnlDz8oBo0k1mV8sfWf2wB
Un6tbg5PpFFt32YY+CkjzJ5GYQt0ATIZngKlf2+j86/dukQp3SGEuxOw2osFHKY0uRG7QZV0Prbm
Z0i/mfelDcFOa3f5tJbbQOorLOGt225zW9y5XrrwMzTrpyuLDg7Xh/d0UkS8QtpiUr+LXaUnR34i
sAXqQwQL9Lsp1aALPzN4FAB2BSSKYzkmTKy3CZP/yhiQIn3iBUFdAum8XZbMiSZdZDh75WOTp2yY
9WNtflq7fG6+xz8U5ki0SqAtEPTsaQiNoFzGagNruY8GUtWa6FIb8Zi9XiDHD3IxNV9ahpajtgpa
1B4a7UbXPTwuSZiqAXZwoGeL/B/JjMrDzTaHRcZ62aLShNLYm7IRs/CKTwQydADc+VzE641ySTcr
nVfHFnvBMIIWmYSGB/dcHdsBfXNzt7E0C3KtdWUCV+9uHrn6hX+aIBh5Xa/YOtrK18ZwC+7rpESt
HHJPkmPtoNuSg4giXU8AQ3j2gqnki+6dU0gR97joo1p96wASM9tYg7D8VDI3zv3AmBDYAh9GMQlK
y9Q/J4CxtJFjFRaPWpAw347LLQYCIvNCRHyJT0GfBML3i2poJFkktvQZSWg1c5XtE0XBfkFjf+zW
rXEB3lQ/XnJRZfyQRcAVmwzz4HjMxQ7hC74Ox4KcMkEGZqVCcp0YyNLfrzZuu7DdJFLS64gC9iej
ZmvG+EMwtaW2P8X4l/FniG8EX/ks49LlkbJU6q4KDBMzmokW3u7oJQT78I5yrr/bFUuvyxVbarEc
ilJVJ3M5l1Es2Xtv8bAb1XwW+Tbt83cmqre8ZcxFBa8BbErotL4/8PPH9hJiIWlpd2wJL0fNRjrt
dF6fKZjfpCl2xT0xUQnpJ6dBSGtj2Wxh/VvrhdcHoa/v8kt6+zA+zUb5IICofHLc6xg3M/kYFpAd
03lQ2V51yZ5GZC9i4WczRq7UbGewa2BFJnMVYCsAoWy6XcNjiu+pvuJHlIxzx2ecLCcBxAWJglng
smYtsIo+26rFwTSo0kO80lQN+YSUidBWp5PMMiJhk4FYBJNL5FCIdNHow6mZVZZRRr0I9VBTwhds
rhbP5pY6hyyGslpUnedy4tPbziM3JDG2I1Jq+LsBaHcXlsbAWn7Aw4+SHBS946C5GJYdOACBEiwg
qrt7O3huAbjJM2GozjJ2Sv96RT+3cL4o0lxRrbHwEyoLUZA5Z7RIrNl/SrNN7DRv39PejKh6T9LJ
sFm737cBMZy0d/f55kmEdx6fEQLa+te5H9NXELEIDQlpf7HFwGhdw1LJ+fWj0UKKQXE93FyFOhnL
VvK71KBw/Ft1mBzEIy12A6666e695ClsChKgwRNZB6m0kcaIhVa4feNcPERSJaTO5YiNBy+Yv9el
h1PX72ZEjT2Ozao8ctFipHIoaoHbRuS7khwLE5DRilsfNDhxEnVsaWZNDKBDo/ID3xAFQdfJ6mHc
VwtF1nB1K/TIXeOEKhvN4+krNWaD/LwCMHHVA8AbOfJrk1E+UceXhDoMxhc0pSi0nIZIJ74wr6Qu
Na+H084bxQE6Gva4rTKwjHJMgOgJMqoBtbdycG59kYDsPfouoVPsn2L6E/jn1/Ba+h+gmKcXU7LO
eBNVjFyKgNA6UPv5jApzzzX1x57m7w/Yy6LzwSedS7LGYCDxR6jK8wehZvHMkanPLMW4IgrjIs1T
G74AF/lopOaAG3MZefc+tTGDhqxI7t0pS5ODPeJNCk/HstbBGuYZdbpMpIciPd9IkRtQjsYeAjkK
Z+d184RGJhf6CCJpN5M54kR+UAqliJWLKGfj/u9xcFHa1YSdZ79dqlt2J52u8DHCfVPTdsLalQ2d
6hoAIaj0jgsQdzAHe6xCmJGdDswc/53xlbFDiKNnDlfXSRFFGWs7oRUTwB71YgvgPzEsMR39Q4mu
rnebVJ0SpSOXD/MoVJzvDXN1l6sMOIfoNLdIZwRhtln74hp/bk0YIoLwszmLyD06BQ0IXpc7JApi
C+aPKRThO6wyLKTMguijsGT5kNJGyN2OddN36waDsfreCVmvOYOvxa4oLZlLwcf9wBfr868Uk2v2
S89P28OkMC7CDtrbJcat4Za1+46ZgsJWWPZmXekTuQG3skw/zRz19e6mYD12Vfz96Q3TUWSsPTiS
/JK4bxXzEDtrEB3CTZx2Z1MoR7pqJ1C4a3GJ9+AZLKcaYcsItsHBA4bUDn4X5UWKaTBRmq3xFmue
DNk9r2LzXVnfvbAjyNvxNlQ9vRJVlCXhe9kymj+MxYtoBVJhNigz/DpbgTcKQaHuWXhxit8kg85M
hcl/LQwu8Wl2TA7NJRCl+XIRk+gjMI9cubQzrqM8VqgbA6XQvQyA1fIglEL64XD+sa6v7mmJj5M1
2XwC4cGnPH5BSqhpDqCG2jVz0kdSfAd7405yZEGSdmX650+g8PFItWLry8cQx+igvGq9je3xt0be
eE0NNLlE8yaQrIwKrJRFFdaQ9D6H9lZar3AZ/IlHKrb8ZKdZe+3iX4iep6zZfiZGbhAovIGTa01d
+hEGYalItqSh0EKo3loitQdGeIY7LtVRywrEDLcvT+mTQoEJuwd43Uf7yx54N3hmH30QpkUH5Ihd
Tor7WjTWvYkAck25/AiswETP4j7oLt7358vJgBKzs2FXdbvIr3++UFIh6VzP3xBKeArH3uPmLvrF
ykJmNtxQPYpgClsJn9J0F6TczkxxEHIw35n09wSaGuD6UzUmFfvjShIW5a3+/UrZh0xhWSqN0+Fv
FvPd/JWmMqCFksDxqwYkoIlrpREjHf/Sgm2U9WLTbDa9sTqCEKDb7UWzG+J66mE7++Ny5mklacny
EB/bEKHr403f9lAIfxO3x38fbmgNFVgjhJwzQTCYENr/UyCAi1kUHh6MIhoudALWwBizdLWU9hta
sTaU4JLvGEjTqeCCNNDEbEZ9KE0o04AtVMvYjRFpGtwaWuvZb8XKOM0OPkgj5pHKKNi9A4jLHfsw
btHnFgT665GLE7yIBljWz3XSKTXRbQC4WwO10jjpyyFOFGfqUwuYEIoIxdWBguMPQbA6D9xKDj3E
1iooLNFlCCukfFDX86RQ2jCoOVZ+VwfL1aidjSMyFs6gFAH86edHY9WE44wR2cOM27bIHMXqdtnO
zrNheYlRZkCSwUK/IfZUoj4N6wHfz7wyyr3k9X4eWTLEbRse2NRc6uK5GXsPnrrxS79NbI6+ZuEr
1HmcQ0iCNb8EwlTVoCxcO5/r1IgQiWtCU2mkSyP4bQrLMjJ5Gtu6EYRRzoOyQbWQEl1wDJ9XTe9Q
dnRah9VxTXWMdgQ895fJhpF4KtJ9eQ0HZuXPyqYj/3PJRHmsFWPUIk4/I9pSnTRdxr8gllHhv53B
je4NxCLRBBT2kZd1T57QCxCJjRjRHgwNumlkBvj+p8qvxOS9/WEhBxEVrFVzms15N1vsfUGc83k5
V87gblR6/cfEDqSBCSB2WtdjWbULRsd/g4QQ2m3QLCDEUEJIj83f7/nh66ULfFOemutzgHXBBkOb
brswPNV2YVUGtOipvz3YJmxdeEDUTi/jFlBrTtwLU/LOTNddwkTMlsxoKwS6dosrqxlsJEnWMR+D
IejyFwdFSBIsJh+AeTkor5z9oU7OL6AtnbRI/WbJXLqrVvI5ZwIU1Zsgm18ZYIy91GenIkggdhgB
mv8d8n+VIH6QoJvNdMOCMv7daHC9PHYAIJmopJqWofLqrJnrFn80x3Kg9HQJVMG6mOyJCb7fmHMe
wM3u+OtrSzYQCKuhig3sdqgspjJo9dlPJMSpDIjqPqF7z2GQXNCdvLvR1omuLD0945Z/Mr2Bp083
h/sIVN4sSUiYdnE90BVkV3nQ9BHEVwxBcwsNuCTm4X9XANc3pUsN91zTNHdh3UtYWxPJj193/m52
8I6PFg/uxUe2EvWStdkqJltOYtM2KMZkq5As/ZjSRCZwxhzl6goc4MTokj/kbFzZ4i0Zi2ohVO4B
CgxG02tAy3uG67D2CXWAtc7InYyeEx+iIwuaZUVy8Mf3SsedQ5GZ7ab00a8PV+JezHmdpaMjYUPu
BAGUt4hUiA2nvKzKwQTMVAf0X+I9aPQzh3V6C6eUZcMs+OlYrQiF3XVaRaReoMs+qkHFzGlKmm/E
XnQnBJcAMSYCi8V8PAfg9T4JvrJt3IFUk38vu6sd0MAisP30oO970u64De30skBJJjPfW9Y2ic4e
jOQZxJR0ZUo8qyY1WUziqbNeuiDQrD9EN5bWOPtEJvQw+G6wUU8TrwSQqR/OI2pEAiRk+rRnBgJa
ngm3zIJBwRXX9Obz+CWf9g8fiKyGpUgTHgNUy9nT8QBjU3ZRsFHTIYSr+56cP7dReWtKzm3J1RFI
OS2HTYFcPC6RbG+j6pRIXZosYHiG/AmrKTayIozePWNXJgVc4GslNmvStigswDXVk1A29yNSRHju
JrqvsEwE7kTyay5we7a/NmpaJFNeOALP8Hkn//1WqBeLIxAslkJzRI2hq9Ti8ZzEjm+Ir5Y+7PYC
Nmt10Oa4nNjhccKBIYuTjnVmoU9BhHDYcrrzN1GSvLm6+F9dnTmjYr3ZF5bH4EhLZIFPajxI/v8U
DWIMrbXpD/7fiuyw2Y718HWLYZEwVsI1s/2THpUWOmxz9aEVHsClTSRDfWNf2YIRJHQxEq84UyoT
GPoBlneVfNwaOUgYTrG9CAz5Xbd1MQJp4fOD9vELLyLUC7yhbD3MWG7yh02pzt+iCxF3deRALbW5
/CsBBp/O/tQj/A4U7cZqvwDy+DL7hTHPRKo9/QFuUScoCrPhBvV9C6b5Mopa+EMsTVoL9g8wj8Sq
0cbVE4OOrzuRhm0nemnbpCEJUgaJ2rKt5EZqeH80uCNkS8cfV858Fxj0aPdilRh9tMKQ/eSgRu9W
3Y8/SyUpp1wsjGhfRzjJGiXi0GojtEttdTX/FsucUWZuWU+KojSaxJ+rldCdlQtBSJqDONq7uGnT
8hO5Vehkd19hYHA9TXM+XXlGkQgJzKHsCAA/m8HoJ17Px2bxViFrafs2YoKKv1vKcHjnL2/jlTu7
QJ8+I3qeKA2U+bIZAtZ8+BRo1q0spIeVpYIVA2yRSbNKWYA5SG7ePLLs/xKpuKTcmeAc2pUPq6Nc
KSiksA1/roOXI2GSbeS1Ti9qqZRs0gUjJOLlyLsfUl+lxi/JqQOTU+1ckvMe8o4TOqfeu54QLYM4
2G5YVn7C0/JirKchQOy1ssfHyOsO6dMGKY6UggQjIlTEi0Y6SeTW3uRcPLvaKA8uKPUQfYslPY+b
d+LMoyQNJB4saBxBD5sPlMNMfj0WgDxQ+CsUD1qFlLjqBtqC6y3vMjFB0O3LkphW22l+irXgL7wt
WGxs6RyzdKa7MmquVZjtOuhRPe7paOmuA4+oHZCu7PUe+99vBJPhojPsqQI4+dvqxe1/00LWUksU
tYriyMcr2C4+ypeCNKuq2MDu7gf4xmop5P1GGcpLmjo2sxdsln+geqoczpsSwzE+ANl1UmzhksjE
ceIqfoPM7sasPSG21FHKoRXqrlKSl08baTWSoFEf/A/9Il8tbHxvlZj7fPKbzTUcy8Ke9BTpjyfG
6k/axgIy3JLj6OyIjSbYtCLDNL6itJbtRyDANmT2ZhCRvvJ/429RsjNfUX3xzKVOViz38/rlud5r
F9XkbZz4oqZnmmARkWEiMyCJiKP2pHNF9rR/sMW+yKQ8zVHASb3HWOA+RMPLE2o6pqWG92T5OugV
hqTV2ueIDcOwai2OUXae8APke2lCMrUgTwc3bjbSVUGC/HmiGRmPFtCjwN5V/WnCpOuqztKGpxiB
Dhs9BAq4GY4lQuHr6/dG6XdWykKDHgmtcoPsEK6mTjANjWNjbAN3HDe0LQezFhtw4wI5jLjtxH6Q
wgzzqF6wBjwi+0TeZABC7C5/XN1GfdTGP2S66jdQbvqt6K59SHMa/IiiilWQqNRuaQkSygHmExNb
06fENSF6zdEORQ4K5Q+/4lP51C5gUsVt4ul8PBroeMppvfQLJNKCKRXRkfpd7WCqxKYX3mQPq6MQ
DmQ+QMncXoqYstgG25Csq9Cjk5jOZqrWQDc/XhBEYZzlEpngua/F4OxtdY+ZSLQWJE9xlMy5lPAj
cBkyEIgkKWaAh4s29xOGNuF3AH+Pz0AVY+d+aWN/K3nCGIl4sPfgjxq4/Dvxmfi3gcsruF6K4rwl
0lMqNGbrbH0FCn8Vt252bE6L7x1c5s/sp3jZA5pJ0eZ2ivL4UAF2Q8aqJe7BKOPc++6VNL38ETIz
dRvCyIP798LtgwKT4sJMYUcEfvAQBLje6GCrFx4RzQtsnd1Di6/QJpLsp7gCxo/PVQTi+aY2d+pc
gFN6yDkZ4ASklTLM53T8jtcjJSt63k2Zak0m73EREuYDXZPKD63tZaEbInjqOAT+RbEcGClFfC5h
n6KjBKcSwlf6uHtzwNl9FSVp2sdgpka6NGBECq4seIRlDQh1HPHn/YXnfL46fnidfggCGsSUBVPf
q2Zfiqc71qrMs5omk4mlGULWOEgFybyEcRGP6NnmVsN795XUf1oY05jn8nImQ1N2aOMQO7Qc0TcA
ilu/Pn6S/+iMVUUp8mTVsgfqqTGbsFdvzcugvEnIkGbIxmtjNFvXFxDRIgiogtKO9sWTiAb/OTy3
KX7QmtbOPfSnzMgEmcj8ifVr6VT/PUbmWpCylsy1l2VvRVWHwY3OaP0HQlFOs93mrRhb8BeG+rUJ
0mT1zKIXkGkiG+0GqNsvHI6gWfcdwVsQZdeMspdEIXifv6UC9OuHx5MCqFBjQJYWV1yVacIa3DwU
KzNJk7+a9oiAGYQlBxcmZe4DLjA+Zbhsn+o54Xu0qHE5hIkUrvqxEKXEAO7t+DC419goV9rHhPPq
pOG3WrG8Ml+D+d5N+8+2lgL4ItefkTGsrjQLQJG5UjuQPYRidaxMie5QM8RdMwM1X51D8K+ewgx0
h83Q+r9GGFlIcIi76m2b1VuZ/Go7Zgmkd1lnBpC/u5eyhlQeUPJCLZDELLa0C9+Lu9MsMlXCtIYq
4sYvfEpb1MiNNOFW5fpN7EJJgiYSBkRedUUomHrZTbS/GvHkPR7YD9fNSin424zQnD6FJgNfk9d8
MjmrX+AJdT1rbCiuWaSQkyZMfRbvMcG6t3t5VKRXxnhtrJBTKe8wk1CfzF6HsoM6IBactltTX5RV
dcbfLaxHgNeL+hqNWEhCCrTO0Ievo+cXUf6svdX1D2yVnXKI5voTfpv7IWek0yMWIUdHJgzFNpzh
FIi2t3l6Wbm+7AVGgB1Fl/Kn37NoI+5t2IZWtdDJG0T9R/F9J2lMLBiTHaWMNkecajOdHCCgW1cY
NptOrIPhVfJLOxB5VE43ES15IL8o/rjzofHx/r29+xH7ABMhH/TUd60c9c06LLJOd/PTwqw0x8jG
WttZ611vsXpKg/j6hmWKH60xRk5B+xy64PTd5CAvVhNsBaco0d6JxfmvT/CJki6iLiIbP4+ifsU1
ywflri0hCiOg8uoJGgvL26l7Lkg3mS+PyX6jfvvA0UXNng6rQ8f/y2ooTzSE3RDinE3OjUmFxp0D
u/wkrKNzmuJdnMw+yn6I1K8+RxfhoKcwKs+1tKeFwZUrboEAKc69Pem/alhy4WkG6jNqVEj2kA65
c8ioymnwNNhkcqC70FIHtS3bP1scalCIKvzXRv1juEVKB7B66f24nW8HAChXBeZ3bXxBD6PPOFTS
J6lw1lLT2/LkdylwacjDt16+0CbUJs65VHRT/9vOoKkXzN5p4BTvDT3FGl3Vptq++vWqsIlDnKN1
4ovZuGjXUl2lS8L6AaQEckGEWiKgC/wnTc9KyxEHAYlbnjfk2RWw0jSImfIHZrDDyjsc8VKGdjTf
lCuxt4GC79w8PTwCgHa2se95wij0FJU6cOdDAJoJ51cCbasPl7SfNBSBT54TS+9p+g62I9Khcbtr
Morv32MyXTATJaFxcwuI7nYv4pnqZWK/hHe90QsQXzQv7oGJvHNpqVnfYI/oAQQ0MGoFw0u/x1Ro
K6LSq+AfnlSa267djsYw3EKnIhihglv/pAKNtKhJYnyAL6KLBZ0zK1pxqXJD+MnyIbU8/yTWaeHF
szdCr08QWIKBFvQyXW8C5+ur5Ykvu0efqGBwpVTTXhGBaQsWlSZqtZZY0xLMmEq3ct433mZPfn9F
cRQmJIZoiHopb+3+BpUu9W8xhmAXaCYnstb3yBLRnTNJ7GmhBs76pY2xl/472f+6a/1R/Q/vCq6x
tvc+RpOYwMHQNDMv5CvbrD2YH1SQZSKWdZfmALTJg7qU+KrnjSAXQvp+/fjuHUFB4ws4DXaikNoG
OJxYIfiXn/RqGWUMWU7zP5tUoNnjCfj7U8A6B7bzh3eUD27kKzItLM5enVSUzB2SlxI0jmGCsNlL
NZ2Qcdw+RZ/ZMN39FMo+1oKgyNJbL3brHxpe+n/MKl7e1mFgkXJze0vFtPMDzMBlK+EkyDN/gYPr
khBnh+Hn1MrY31IcCnU2S2klj/jNRKHjy3QxUOC9piAJpZBu9zN1ZcBme0LLTqfZ+kZGq4MkEPHF
Y/2tdFGe8JNRMRiWoIJX5X5jizn9lSvMzxiNu7h2gAnm2r95rVOwNB9xX4W9TV9zC3gMFMLhXtsX
vHXXRIqE9GEbzlwKBAkI/XkktbkPO2Ee4EgZOvmUrViO4hOuC2/rAGv62AJtsoQ/FG/SapTvZkHX
LVufjNWLjfs1AEYKP5sgpHxJY+o7XdCZojzjn1yeM+usuWyRvozRxpxhAmmiEPWi04T/3RLcvvXA
GSuSElvpc1ufPvL+zbVjBW9l2L92y6Hj3PvwBEwLgBmaAnc24MkrtmCe8/4AvigA3mpC2IsIP1BM
/9AvD7+uztFSG1QvAvWjEtodEzno8o4/cwSsdqjQOpWufmo26B5IluQdZveAVaK9Om4mwGE8SRVH
vkisCpdWqm7sM1Rj3GxuElN6JZOU/A/uGXZFzUjoT7ChNF1KfdDLWRhmjr6mBOVoHMCVA8AGv9nM
ot68CP4XlHxiBjYhqmKMyQC9egxmGNV74zUyj5JG4TgOaf+xxYPniwSoeKy9R7SFA1R3tJWk6gPV
6DryajWDzoadNEDNFE03uE4DsYkoKHM3cnTYJEs/+BXl8kkxh4pHPVoggCNf7GF3S0s/JCg5+o72
gDaIm+XTV0KPRT8QEOjTi8KN36WMu0+0wPn/dwBO0/8vN6XNOHuu2YtTP23itPfx1KBo1Qi95ub6
CuNN60NRbrZbcy/fbhO4+RFZzTJAH3UA+HREkf3uaIKyEfhaqVFj5e1BRt3QcpHaioHaIPLxGjdW
NHWR73066HqYS/SHXtZA2y0JivgPLIQqw2XWRmEm1CH6cIvw+qx4UF1nfnQPm+swDwhmOFnudUlf
PYTdcTVzvW/AD1agOlrGq4Gew02BTlhs9Swe+rjbqmHG8ESnmi/46+MjgylnmPj5SmoxjtdsOSZr
zlIu23eN04cqkoWU2r2E/ovRmanxOQFcC+O1RKOS3uCP0xzT71HZhsA4ZbbRzBKE/D2Od9yalAzB
8ffHDJZAH4WqszNRodnw6aT1A54Rs+g0UYVx4tQW2SqV3VU1HcwKG6pxHivzB0W8N7fzYGxUNf/e
uuC+9HKZEVT/z4hD2ZlF1aY6QekPQCGcUxXHYw8CnC/i36jnjGy4rPz2UVwwkjQI08NwAxYQbIJ9
UfvJX05jrpS+58jHHY/UcckYeKH9Wq3v+yLFaleQ01Xva4Krht/Tqr8pzkKuoFVqJ6JkGZo805IX
R8P9JrXKSwbjx7XJXH5tA6GZmEhh6Bw4uZ3BbgQMDkZ3ApB2ROyrv8WA2jjMaiZ2baMrkmu1mdaJ
eHMm0gooPBCRAvlWVj60EpcwfsKU08SACEnjSmaTP46EKB9OIQ0MfLyyAneMpvHEOJD63pcLKIzj
04AQhI3rfGPnahGzpR541qvwxGOm2QonoH0t31GDiiF10KQRavN7EH5fmb0U0DNYWTs8bbKusQj4
eP1TaF+ByPQUVtWr7dKB/fwOs5PDQErwkGGapPrbRNKdb8hXviMa9Bw4yARiDijQWMIFT4RWfaWH
bGh/TXZtwZbq5JQO0iU9yzIYXWkOBLyOI+qMnlsNdiy1Z2BT2yckPYLYBbyxxV2tFwqWbthHE151
n3CjxQPScfrPX9kMSGw2tW/Wd0W3I0PhuAPZxHzp46WiKAhQ07wnmrMWtR8RCPdItxpT+sCLehCA
rKE8/UUUkQvqrJpRoae+lul85+1hmitykQEvEF696mNX78UnLFV9Fdlgdo8yHC2fR3shMaXz5B3g
cJdjd3klMxTG2CMENwbxwvaNFJDYn7x+0SFkF8L+hBjKWhRJzrXciRuPWgGqSSrZnbkKQl08JCzB
sY90qpuyl4U6cJDQrFcdHGht7ZaT0WPCOE0T3a7wuJLZg+DgWKcF/uYE3QCq5kb3P8RAiumhZvLK
qCV+8/OcQMALESO5eSUqW467gXlPvBMHiIjhYc+93/0WVwq+Jx1KonhvSsb3cP/S4OSSMf9tfp8K
9ae1up1bkFMbaGG3ls7wLo/6DQPS/jdIJd93+hlQcqgnQRhxWqCOccO6AXwrTU+/4Ppq387rqwmB
G7ral7+0jEF9d0mmvhNGPnYeTLtEY2al+X3AKv/c6PoA5zKDBNOYdaAW3CAVUMi6WCbW7MAtmxm5
vF/nba8iuHPT6/SuVzaY51t6FtzCR8F4ImRkeIOtM3yyfLfjMF6OKypd+Ob2oCD7emApXF6FMRnN
le+u3sIE75MlJ4mitWzTF1zcKhdpcHpWAMDX0qEF0b8CVFLuBT0bXg24AaZRd635/IXqY8KRSwpc
OWi7feOQ5FLLcEH1qIdwp+GZl52+qvBfJs5gRUjnZZ6Ml7xVE518x8H91cahCfHp02A60kDPWVln
hx2av3vIfBIsmbgHJqyLYz1333vJ5i/578ADpt64deykeSiNl0MimoIXny6BbnDLMIdyzyV7UBiy
awcBZPTwdO/BpNhvsuki2nYrl/i8LA0cqSDt9suPraWFJbd6yaTs7i/+0qR5Xn0+/JkfQAjY42/6
TAbSiBsOOjWi5FC5b3EHi5iIpB7mnGciLaOE4czgz8R76gEO9rZAZDMkachL4TfiaXZ5NBnjZGi4
jdwOjgAOxxTK9+6uOdvE9DyPl63G0nSi94cm+LHDWg/qPnrmVDBcANWKk/siLpeUP2h+eKvPpMeh
buOmWLn38auzhVBD1MTlZGJBDTr6yqkOV0QEjLQaGB4SJcxoddt2XCWRe85thXCjEMm0IjODocO9
UHYI6rKvIJS9TV76ZX3+frbQO7jSuHYxJG2I4O8retVZ4bYr7645YwW+k3hotfjezfcFT84ayrXa
wNl4V3Ca2xzWoA+qgmbOBu63eWGYZHQI1C3ETFYQM2ShL1hkjMruFUJn+GTD7KLs8P7CAVTZIA4m
XNXl7GFIzAMeX1M9kU6sPWrl8oI0jbxH+YAUu2IvhZFnsU7z5mguRa4XmSSAybyay7jBUXRYt318
FzDTQExnmZjJD+a2Rh0wrsAyT/9IAsuXT7cFboAOBzKzQXH8HHVf9xXkjqywPoPcAylMCcaOxW8B
VRcgZ5zwpjtZAl98w+UD23RgYwVkdgoKosYM++PE4oH46tj/vg7KtP9h9eCB8Z2UxdcxMfkncKb5
qohZtC/uyJDmCgO0vhufbZiMyHHg46FA5Te5XUjeDsW50FN0IE6gAZUtMLrBuMp78vN/Gt3TNe46
sV/XHoBQshHBSNPGKX8+3ObJemUN7hPrsLQkWHMm8ImLfEMA8p8e+daA8SyaWV27q4M1EI408RK9
myXOf8I8P7sjhb+UqTKqdztKyPSXFHGFC6EdvE9VzaAvUAr+IiDQrWYeXN9VACjx1MbobwSgdr62
ySV1VYqGUrWWGpfdDPHqn5cxh3bKDOCEhl/ZYdNsBFSpphW5SXgpw6WZzkU1m1f92unA0Y9RXhTF
/ZBC+V922gFSkkGM6ncgaZIIE+mh3xLxJvTCPhgkbZB8dufh1HapyNCkUNY1eZ43sapVOiL3nOm9
zJiBqGXojpNvR4gDiuV3k7oFuublb2zqux/AcMikWg5CXiTNvUY6ZC9A2XLN07o2GVQaqJkLhdzP
naRio70wvczOdHl0819rKtfT0XL8YptT+pqmIYFpHtoQhC2EKgAcZOb2H1iRDJ3NuQv1it4jFcyy
BrrJmhOSoIA2llJrJQD2fb9X5Iwat8f9DW3oVd5w4ZgArDRVW5JpNRrk8fSvVuUVIRI8ZfHCm9M3
a80STDSDwdEscNd2le3C95ssZKo4GwNP8OMgu23A+cjJtxz8NRL+KpDRJ9W89H3TzZ6WFfCqmoRT
VziokeQeq7QzDGqOK9FnUgKRxpwGJbzg3R2oyWVKrz/vCG56O/jAVyz9fU5nLFkfkcurqP9LdmBs
7iEerXi6LQ14vGCUmzQzjmNI165YPQhMAaHAEI4igSOaoUM8AwhLBZkJajjwWe9HzyaelaTyW/cN
PJAewpnUzonGsaXxalNVJmG/3chqk5nfSFTUJIno2ENfuD02UYafNU80ISqJEUer3BkBBbpJADCS
1JGTqwRUBd7GYLtUNSw6tjTSJHtnV77x+2gbA2OuaqdCWzLHQf49zjFiogd2Kuv77DKp/AQTZ1Nn
tbxRYf9ZclIbue/ulCfEooG2WyBaJs/Yf36hIyfLkoUV1Z0wjI19U9Opynq+KkVgA7WfEkbVM+9w
AcrIfH8yI6YRzwrW2d4mheGG/0R4rNzNckmNd6wo6WxgkQYue81JGW9GgmSSvFcBMegNgFxWhz4z
yoIO4r5jKzrWnyILfpQ8tNgL433PAPxZEvkYy7hQWpMK6vVpeRGGCC+ORiUdYJZ945XFcaTPRyuu
WJd7k8c4FkoEWe+vXArqvV/eFQ0sHaY4DdR/dcsgk/YU2YkPzwFZLTI/P0xMwYtCCYaSHJY5R/h/
CFW+rS/ngFKNYfyl5zA0bkP/jxcQwMFgcjpw7DDOZgOcX8r12J2BjUoOGjtoVjXoqGuvFbRayQW0
ICMGr47VRQ+6LR8Ka6IG7vHODiawLtW8f7XW/wJJ1fT3IPUNUb1wuaT6DjAO/cXBg0galor2Um82
KwHBk75rIVFBgE1ULlDzdMdzidvGYPp/4gdPKw1tJMnlZ7UNx226z/dJOYojj2Tx//G0VPgRxBqp
eRrhUn5kRDoz580d/kkLxd+9Wfvwb+8QlOxOFc1SauTORO7S2wvYlcRxH7QWWIwqYs1X4t6SzdrM
qRKYozLImqqbYf7d/0T0gfYloWJP8QzLht60C21qXuOdVZA5w9uSS5Aq62dfnB++IcbBmOqqsYaw
e8RByi3yFXJ2ytFL9iSSeQ7VCXDklpf0Dt71Hpks1hxVBIy58OtbwWunJYap4xx4EHiMWllOHCYg
rWOQv1VBBsxBuzNCIo++dsbzUXkMzWAQ3JCgoDvJ3UVd29qopCrlgagkm9iF3oOe8Ml92w+C2LzJ
PTxSfs0/has1wd69V9Bl86SzsNd6DWX6eI2EbppXEEAIE8tQcGh4m7QlYo8wgjt3DgHj6J++dSoi
B+wWTpXWoGxHRdSc5F7BQB2pFhZ7/9wz+EyJdvr+DhgbGNmZ21H+FDGQHwHb59/LfUfVUdX5Re1Y
KHr2tpsq3+2zdMnjP2s2aW2nGeRM6zALsWF0qDEyYRjGGelKqQUpYIt/otniTrDx8p0KKg1kg6xt
+2bTJIPjvzcc0cc+KZZOzQSqSfQ7Cg2PGZ5kKc2HudIN7Wh92FzDlGyJiq50IJuRwVACNnLd/Wxk
PImFP3WB+uS6SRWEL4h57yPnpdE8Rav76/ky28CaxVRi6wJpwWa/bTdgNUf6Vv2BtoCYkIA7IrvC
DVVYRhAJw7Tv1sNIrI6R5/2xV65M9+tpYLIfApSDeST9l6qNhQ3rTuGbAgLYuauaz2Z0yjSPOeqN
4k6tAakD8+8VjCyL+XH9t3EUHTngztWDHKLuAmaJYfRoJAeWN/l4XRQHvkMfpl2Um/i1/eyx/hPZ
3Sionwn9rRcgaLJXeWCuVAXHaWl0mUBp2MaXkPbxpHlOekJP+A/zp+tE9WanYoYkB5F/Vz+YAgeA
lFaERtuqWuS87HOKZhFK1yJYCEXA5gElrdq6265bam20FxCnGNsNe8IittQqdr0w0R9a6aYuTrGH
lCrc428nSvVH2k2135UFaFG0++5MVg/XeW4V8v6cBvLMxNNioQvJGA4r+BzAtDVW106eAxrHR/BY
/Wn+oQXMnrhGOJrvhmhHGI1udJ356qKteyNAIIVh9KMo4GV6LUsQzYexi0xWv29rSvJWDRIybGJM
dKgIcTYWZYDKFyX4emQm58nY7QtolSXEv4Fn0Po687g/1O6HyYHqHBrz7y7dPbNhMXrOji4B3yxr
Rw2FhkretY++W+iWQ99+gd7hwSAqH4shU0ay/f8/l0cQlAvP11neaS4tnp3Kb2q5dtnmIuaSYDEj
N/9Jn847qazlkYlp65oRlJ15qrY74T5PULRvveMco4cJYetPmE5fiAmM0BDshUYtFnl6HRMvm065
mvjbcmtYwh59InMFyGSU5sWsHSrRiGDkqKFMpHdzGZTcRsYenRm7YEmzcMP+eB4L3aTIO4BUIhfv
B761+YsKTGM//KjATOMbmsgm1pmUF+kCvYcXweyBXWvLY2IHuQk7oE6zvRzYDS9LKUzTQJAF1ieW
wmAjnvQm2WrtQsEkTqqAZyc3Ls0dqkpGaMnRJgjUqKkApigXFfzCzjj6+JVNqNHeH9tmgiH4SitQ
kiYl3qTRN06yENHaZstOoWDrKOYQC2gPdMmNfgdD6KaKBpblhL8qqGFzj4sYi402izIkRHaI7aWP
Qb1ZylDBn20IqZ0gB1o/Wq6IE8+lLHEa55WJiR2JJV1bbecB5prZn6JWUKIIMFr+SSFJAsJCLJAp
XkNDnTIF01oskEQSh/lpv7NZV6LMb9IVFuPWrBx/QItWsjcekVjO8EG+r7lwf6kjz6OvHaFsrp3q
s07cecBPrqtzkOEJp/+Q7AOfYPWIublRHWLTYAYlxcSo+5srBlzMLw+C36XZNzupMsKb8j5tdb7d
vIPr1u+am+E6lXpg/6AZrvDebJFmabTglyqxGfWQRVQOEdcD8kdTCmzYrC/mnbP/5aa830dexsPy
QwMehhY1uho9Gt205OUHwugxTikX6Gl1A3GEjUP4bn+3WEJbxMqpEtYF0UBg6UgANluIexNmAhG9
MoP0FblwoyW/VyAaDkh4jSF1zmpsRvNiZ4gJmi/RcjSiDI35qw21CCoSXqPdI/MCL36LySSidJjj
hV42u1H/8D3N0AzpLcbzJscKgvs8oOUvTkRCZJDEw+9nscokhiNCYHTFynEcyaquDKIAVhB/y5tc
XXBK8sly3mPeY4ep37FaGi0Kfd8DAyePQWpj0D6t/JmqJv/XnXZuxXI7icCPaacVahEEQ/CDDPnl
WY25Q/yx6zUe3X3Z3XSwbEYU9D3Tx8jyYcsl0HNo9c/dZgN2QRQ+C0VG9gsoAiWDyLh6K1zrz6lI
7Hs6yKaqzt2een2tzU+1+VMgv8KAkQ5a2BibrfhFLZM8iwvAh8I2Y2hhezuT8WLuSAQdgTGBEr65
9VeyM76kN2Qe8SSU45yGM9BFo1G7QIdCnOHqmNID/w4wTuBXKrAo4De/AhI/okMp65eB25f6ez8Q
a38gvDp3ubWeW3zl3oqTL9zD1xI+nwas/AW7KcgGiQhrT31MqzNPNvEC6IalQoIOJhXUlQh5Szsb
PILgsI6/sfm+wq3cxsJH2eBr5ErpHbSdsZ+3G2nkGV+7Jbj8y64Fz0ZBYw9jhSa0xtZPGw2zLDjT
flSAQpclm6Jf5vl+vMO6IF8f4XgT/gBrnWTOdpRa/uEadckW7uOa/9IXe7NlwHsdLohOK3FAG7sL
VDkl8mOPC1KfbEmJvOw3AD9/JuAYXbGtTQBZXppKFbiUEo0U0oRcS0fwEzF4YqKWt536UK1qqX6B
31M25W7ps66tlcFcpJLAjlxtBk4tCMJ4Ev0Wr5+nn56Gi7JSdwVv03+UXWBrQXy3hJCumCbHpA95
W5csw4ULzaQSjWTkHGhhRZppsfgATYhrWNVNH247CetoIB/rR+jU0FrZR0OtACnZZcyZI3mGai0J
4BGtnLEu6LCQ6M0vLEa4MuD8W2juPMvTi7UCo4GKoQOcIqzQ1lMlDYbSkIPvtmaMCLoczqGhiVcY
cgOp/AZEcJFW0DYoM8g4lFt3dkjVbameomDB0wUBiXy1kYoou6Jko2ywUfe/3BgDPM1irSyulHN8
ORg88DAMPvQCE5au+u7or/dIqY/wenxrndg6ZXGb+cERR5KECuuNAUS3ZVFS55jGFer8YS9Nbjph
xDYSbrJvh3SCwb+kozFmX8+odl8Lj60GuFO0Iohu/zssM+ja83Dxf9aCK4OrlGzYbIMs67tEbzDV
oHw5F9lDFk8bGvYgfpdT2PPQ8kO2YVEbB4r4UcOnYPCwWDtjz7A4Y+GjHTVtBJ/Jv8Nd6yYnHSw5
61g82bBjl2dPhFQwoxE8N9DhM/OTbPPByW9PvuZ8LXPXU/DQ5191mb/znPlawbguxHED3dFjxUfO
AUAZctuENMNgxl7ceZEpsGVdCA4gpb2gBlqe/XjU2cF7AzICg5qUtOlTJAnubiv92bvvdIwfMgoq
ebE3/MGCTSc10zyMD0KCK8U1J8Fmg2zEP2NWwQ5CytVkV1jAdwD/BSWDuds/RHHuGcQVJxZAXoxP
f5c66eAAs2iVWjG9Rnj1+lFfU200HGSKdJbAm0A1EBzM3UUatkBeBxk1VVLFRB2Oe3ya79lRqheL
23sfSc1URa8FtOSwtOQuDxllFv4Xp+rQMNmOukxpPnQvVyFbj3qOhRoo1sBP+y+XhxyWMLKFCoO5
AZDwI0f7CC5JMLcL4HZw9zhqTcfc44fSqlrqNHWO0rigQH+ytviKYcq7G1ZPLazRSn5/I+qF7BzB
vIWnh3wsbUAQD2/jtn9q2KNyymLA/3zz2O7l+8JENnFpmMizoERVPRKf5pLA5Kmd6Et/zSWT1ULy
86QvQ7q6jmLbjnd42sA8hsEIqBcTa0FFdrvu8US0jPYNgP8ySXFJsOUm42smiv/KMN1VH4PQSQIV
mCaed0TjtW63PEN7lwX8LNWHgg7yL5e8znOAN67NVxCbn77dMqPIEsePT0nRp2Yi5N3jBeaxLlPR
B0au0HLdCNafsPbx8TTQtYZR/7jSgPWp/wsv6JOaVb0x8+fXM2s4cp5Ep7VD2YVdNewWLOjslSdB
NQiG4JLtzUGB3PWStToxyWiIS6XdbsmT+N5zS+msGDRjomLtOB06VP904BFPing3zzbPVeIFLszP
mAxA6Q8M5RYYCTWIJNuBWjFOt6/EhI/ke7DII0t3xGgV6qa6DRVU4W2U2YhMt45fU9B1diix3QWC
o7BayR+rpUPFM+T0501mGvRhTfo9mX/Zw8dSuSGPhTApzcs4t7k2g4pCGQagt66U9RhPQg1rD3g3
zz5C2K5bwjjoZiYuhf1uqMaXyb2fPj7p/S0pToghR+lnHMGo6yUyAqzbX6tJTbBOvBTOB/fpI+6z
iDw4h29RNgnZuByPtuba6R7LKUja0OW+lGGF5GCRWdOfxdpPMdC859KVvYtxMzgwhS8kf/1RqMux
wJNvax2qEQ2oOLDT/s4jdwxBG6tdBPoSSr1mcDuNBG8DrmdOEm+Cu00VRNt74Nj4Rst8VKy3h2t0
nRvIRf76zuonQjX043HBYhHNY95wRilQSYzp6smdp0WPaZYNoTvohG1zCCBpg3aK0OVbuorV97ag
0FXo6OQ7CRDmq9gtFRJwY2u+RT8PWejS3sCSb444jWO9jw6DswuICYrBD6IF1kz7+k58DyqBUJGK
ayOa49Chz5yuYmOjb/PtRwGNuo7wPSody1tm5/jp3wySqpF2tCbARRC4h6gLijgISkeHmbU8uCdc
C+3NGbgBmTA1vqyMg4HXP5u1CL6+TkJ87Sgw4sK2VXJbzMEhMiQVVg/EUSmZkk78B0S+gGMCq8WT
J64iEfhgCL4VakqQb/Ru9J6XGDvgM9q6EZFpJC46SJX5IgfFx7S3n2ouCMSU5IAeAl3jqCJ/U4cB
nIG3LXmqt0avsyVWbRSz2HN5xmzDvj91kfR3q+ebzuKdEzzN51FZBEIK7vUtEpUvk5NLgrHiITC7
8gPqyYVZtPs1gK+6seWWiT1Jws5QdNSm+brHVI/yQ64jfrCxKXDUd9EKbfkBverRhQcSGCM4hCBq
7E1hQomK++bv3LRjaBQukYRs+HB0j7NbpKodlPrjHxroLkbZhExVQVpPNrEKoNKSlHbYp9BYwqD+
QOXemgza9eDTWWd/FDKuVEdZlRwUYSvOc2TWYoFZUQiJwriWUO+QCzjLgbiphgdJgJRjZbh5/f20
IUZQlSfULmkLH2q8HoZUtb28zjSj1wpul7gbk2uI9jFBaV0fbbGcYMTZ3A9UQFywpWL7K7zKPQww
iTQz+PVEBi4q+j+yQkh4uJ/QbGLdbhDuOYXd7tRw1hOW0v9aTDTxgWO6a+Y4TTMR59wdm9G/wq7T
6otu+xeluhlrAi4/x6Dxsijg7rtyy0viH65ZT5bj/n8JthAjpbS/ZMZaz0AV55e0R3Yd90zZZ4CL
ty42zI/fsVfku+vOtgIrXz1z23DCQ8ahZKEZBjFYFoXTb7IV/fSwuE3VrVVqml5Syeavl7A1ymrP
RcTj/jqyBAwltZpdgIjcUoT+9VQBBz1yqbzi5FJaiFZjJ+hZR7o6x++1GL7ji89hq4gzF6wOtIEI
+8vbUgLElg8xk7QFk9AjqPMeyXgn0jxYlMbCtq2676Q0fcuYWSO2WQ9GotJFA897Z/8XQ/fNRKue
HL1jY0T8PDP/WnkFuJGVi3HaVLmZWwpeTT0tPm0afzU+N+XZxr3nNqhV+f5H/R6gcgUPYCAsxX0J
VYDJQA1uXgEMmlsMmjxfd0sc2VOGcwNhlvQJvz5U2NN+m0/6kBPdAGfJ+LFCm78WVFkZI/0jO9De
IRgXv3wnBzcniF+nEsafdSn31JLf4Htvt/auJgJgqJhXToBjHs6SD2qVpy32beKffoYP25rz4ZZe
4MachjqBGJSNm0WqrKxjUjCfcu8NT9o2Bui1l8Cn9kL8r2T4IU+TaSwH8bjKCGjOiXZ07KczTWiz
jE1hVTarN0XZKo9Li612oR9ZEhu/0xoaQt1EZ4cJmheW8Sb3GsHgTjLEzv2gpmteCQcYFfNhmXv/
/0tOW52L0aZK321C298gzfQx33q1v+7LZgpWpmKMGnWLsA3p3+bgIghiz54e7fkLYJV+ZCJtt9en
5+8WdeXnMbwrpNn/j6l43CwdtOmz3NOTicVhDlfirwpqVV/aP/sPCbtwrscPvd2ZWaTB10H3RvtR
QrKKQ/2HF5V3Lfns07RvhErvLiStOWKnySQ9kcCqHbudXfNKjRR9hY6FveG4RPcJDS6zhaDtB/fU
3jGyyHJRTcyB3wo9be36FsoGOmDO9zLJU3e7tWq4xFKCKCIGduR2ARwf923cPutIFzi+7HMTJ4wC
RW48Q0gIxIAOBFvV1GNfWPK5gA6JYTjF5hkotN+SOYt6Al7RdjHVnvccWCgwgejbmM6w5dOGegWz
ht54MP3oWLjJZaLu0ksx8x9n/ngUHf6rUA05EdkVJrJcYzU0VhIPJeDyuN/TjmEwIC4uAfseB1DW
jYcw3lJD2UqORutP3yMDJZcT63yWXl1KS9CWJ1te/GpZWEx1naIoApt+AozaiPaJ0L/mUGH6FcX2
UBK7QrfWvPRVegP0gTsmGg1+Hlke2UmMkAwKXSb0+3otXcp+fEOhBJ5OClK5q9gYpN2o85+hxtRf
jKQNFAz2pQ/pXR1+g3zlMBSysXTpmZsCsMPbJh6HhzQC6SCfsy9Xd1KoZBh34ld6iiOGlqpXoN5R
41Ile/b/jiU5YXJbIhuVUe4OM0DGeFf8uEbnok31CFT8GJGu+N9oHsEs6P19TCgqB+Lk8cDGOaO0
0OPeUGtgZ2fvTGPuhUM7KrFBq5ztk+U6aKF+eE5vwp9A+C5UREMAZyrO3Hae4Gk52rrq/3RRGwmS
sMzlSAc0jGSXFFammcsG/c7CwZK+M8uQeb1MSHoiKvLqr9cSHLHMFz5QVT5qDc20mdqIHXRY4DvV
PUSDhGTN8XybB4ZjO68AOecit0I9lgdOU0fVhZLZJ2OyryVijKv59+APPKufzGf+pQ5RhNJCNp8h
Ou23v1/Z6BPr5JVZCwENZ37L1bt5/Jgyw7MLXdyoPQBvee8IvXyyp92aktoxzyWWjmy0TDf/kCVV
CgqKj4maOeBSDuaheGxrj3McUNNncIVeUkDtNts9VxakiP4o5OMDY7WQOwf5hqr8gb2uY+FmxBkf
W+YT20KiS6NyVKF0L+0dHbeZnY27joeGlhxRn2jD567qiT/Y3uU4B+AVkuVxgEVILRdxE8rsItS5
3Gor4fL/JrS96rrwVjqbaT91YzOjPPxdPPGdM7DmPe9jx1g+IQbj63J8drarMrp9GRITlrTUluwv
PGzbSGZNXx6pm7vLZda1xmpNZkLyhx82nCtwYXv87ASOBLGep4yJM4CnpaTG9bKk+SZW/kbNDmHR
KCoyBlPNrPYx0H/4yiqSpXM+1J4DiB5pGWFaiMZ8yq/E0+yFuWpqeYqZnwqAUrXIxbdMgT38pnky
gRpbHhkk5TpR3Dl7vVAG2hN7aG5vurw7UndxsIE5E2NuJG6BwtdV0KFU0kDoNNF2u+JCT4LS2VSP
25vq/mfSu7T7d/BXa1BiRY9pH+X7SBqJ9msVgijp/GnFhwKKyqPII5Kg1cXzrIPGaaiojUVSyc2g
ELkxbhfJldkspo0Kai+3Kt73m1rG/IXLsBQNBpvQjtUCySfaOr0jpVuw15Q4kIw/UW/ka4PalOAr
A515gSIpMCoqjjP4CCQZyIctVpRycKe4jzBc3DmMQB2wBrASSC7cMjqgxRBinyPbYNQEFd/8JKrf
iuaExbUVHuYgVuFZuPIEiP7yeX53yjtTAU5mTKGwiZGwhTnH5tWwjyQHNfD14HqyJ1vXNjUJVCBz
Jwhfzge1eGafNVGm8H6fEmWT8d9CQ6jPRx4Py3Vi0y+k4quW5RXU/aG2qDGedeIQOL9teEidZ4FG
VwMj5CufTjHhihYFuK/+HL3r90Tz+XAv+QZMs2c/O+FYdgp25fMklp6SV74wCoVbvUOTYLaPGXLT
mRSMF0PLWfpDD6lSKeoBjQMTmb/J2xelA7FKqEmN+1avGnSrNKnxZvuF7PyOTnLUrMko0Iuyx+yS
v80ZAR4bnVdkMKGmShC+FVkOKLvT0l/8DmGEZ4l0/gz6y58+WlDzqayhg/9TfJWFIQ/EPNDaL5J9
RGJ+CTrMknBAHnmNdlqxQvuxkN3uSTWaOeZJBABmQZA1rbbUauEIUmf/qDznLha7pFn3Qkrab5UU
mtpUvj3DnWhFT/rErrtifvNI8gygUFEsqswZ5s0p93cI63whuw2nRlkH+zsJ7QS1eBTLlzEt382w
d9eE3d6MueTcVvbaz2AAcLl2GJvKoaJ3mgf01JoYXTaRQY0AK+J2Ee2MeEjtSjPhkZSKGfdYiquG
BysfEtM//oVAnEAzhSzSg6tHse19wb1uciIK7doX1wgBZnPWeo5kliBEU+5/DEmhWLzbE93XlHem
+9hG4/kb6VUSP3QjxyipwDBdZ+yPxyeOHGLfhqGaP9n/V4da8k/SYIaMrhO6/ih6ayF0ZvwzlO8a
+DWTfwGYivbOk+nicUxmJYVL38HfFxFlOnPoDC1Zx0aWeGd43UzWf/XBEyfgoy5LMIbdh7kL8eEi
6i9Ppr+7w/8lAofwrYqkn4Feuu6r5lbblMJ2scpaYSuFciEE2idB5hS2wAXuB90oF3adsLkS+Ap1
Vdi+WsJ7XS0Jz33ThhCjafZUz2bG19T080KyVk62K9PpnCZsIAtwNGIr1+3/nTRHAKs/a9t9ngoJ
swMzQlNQr791Mj5B92EF6ROdwe4sWBpmIRi4b/WnNNBFAtvXZrXgBMYS/FrJxqd2OwYuqxSmYo9S
Toi/u04Oq+1tHbHOhexyZNMe2wT6zNLlLanssGg4u1ayv/cmsl+qKbv8yoqsFzBJmi4wPNoghYQx
oc3vyT/9/ppa+T3BF0r4XNeEcPKn5Ui8k19lVGymdlw/ICnld3cPWQ0fJo4WsuWf85fyHuC5tzP2
H7MsShnXwixYKxbtH3nQ6Zm9f3zxPOV5Khezrtf+lcpX8PAcRNrjq/Kuud1gemWuvJ/Gwnw0SR8R
s2h7XG6y9VZGAFqaZ8CoTWp4ZahtWTZsXdG396naji86/pyR5AlVhmCn5yfj1RQNi7XC17XVw7ik
ZRFWe3xelcuhvJHG6WSuELmM9ddQA2GqcphhtCwQ3nNSps85qGVVlFLQenVNQwCbozmMg3Uwu/aE
m7QmhN4ttyx7Dn/dkiVILH73i+8ylJt7m4RHv9bRiwzvOrnIG9nObglsGqBLCmW2C31rp3h/s8or
7u3Jyb4gD7iZlKWrw2UbGjKdai3lOCWgkm9zBpbgAps8FtmWIefW2evySq3oUu1bcUgjVaiF4ony
u2i3ObkXhQhpp5SBCHDSjURfWM2Prupkaf7Cxfq7GKyX84Z4TbWasYsQCwTvHAK/V30KXyNQgJ3z
hoBYojeLlj5O4wQFY8TPxf3e5Aqgm1FVHsn4WlQuf4Js1iSJgcWc2FIl7gbvxthFAX81mwnMLDHZ
qrwhn2NFMcIo2F4SzzfkZn5JNb9bc8Zje0DtyJqoifxou+IV0rZ8+zvFJyNA8LAKSxT5u/mDAJhb
CR2vL4oWEkCRN7pJzrAYpR4lkqMS3ERtkTIg2iiHjSsXc/sVR3/58a35G9ZRwJvIDC47g8H6I+6B
phokwrn+tYNE6nKIyAFvZoTZwjysdhzIA3BDwAYPfzfPLNLPjiqV8TGDLAdZC1q6bpLmbsz+w+S7
BJ66XaQuK98vZWA14CqlYqaV/V6w9ivwxLNsIh0YEOPv7wQh24OFjH8qCnXsVpRfi9ypSb4WKqzZ
yo2HRPu2iEapX1NktsOtTaIPkT3B48wJFC0juN0CROv8krbbUmTVYwRQt26ubGtt8c31afmX1u2w
EzCKedzqgNI/OQUpg455e94LMWiDw3eTuLjn2TaRqsh/zncOJR8EhWUkx6FYrQQaCwk+PHCoXcNy
BhhE99aLZtE1wXQzyNajDszvptj4u6AJ/8c+QkmGxLmjhryrvPf+8NLitsyRrXcSxM/ZGwHw3hwK
OdwNiw28LyTzxhkdfDQrQgLW99QWe+Mht/BUxImmWMEgAqgs87t7cdbPCGHL1rjm5rNGT6A1I9Uy
DPWetNrcs7w39687tpE/Tp8TbnKG8rLQ9Jx4B/Md3SoWHmlbUxckBODPHi1FwuCXlCQVzTzZr0My
K/GlPLeaIIZtNV1ktnspg20aP+Ulo9QbBEfkKswFp0xIDhU7omXEraDCPQgTC7aDvfHYmfQBr+au
hmL2w/8lvMpe1xniQkdLuEZq2HWHjYADmWCZeB3O76UWx7CJVEn+I/sx9P8gr5HD9Xbawf1MWMkc
ckpEFFClrZUmI0MHOrMgB/MypBjsCrQwQmJnmBUEdkhM5UrgeE+1EqEcaQsa/l+9RKQYXh/dNHNa
n9jDR0VG5lGqodYUGLpPJd9RTvLz/ct2LXWJ+dbKZQPIuRPLPGe1NHbHsXtfKDbPH0nD21wMDUoR
WU0xmZ1hsfYanSIuKIGoYuEjz54JTjwSLgdTgmY81tq+vKpQw0n/GadRTwUCaGFerU6bregMqg3L
SnUsT9BM9D0ecFoVdsoJuurZ9qgwrfGkRKCpdiDSGnl2mvDF5CYL8NVHk/vKCEnqbDHL32SHUT4Y
u4UViMhzzD4FZjpiatfhp6sHpv+uPv3vl+LvJeeVXk8p6ts1X83mZSUBZnuQJDbBF2caXRyjv+aL
unmjcv5bfGI/Z8hqtxf1IiWbAZJUf+QUGUaVjRAD31E3dZhzaM0Smx0FJyKo3SeqQJ2b9MFEYZ45
/lwKX23GSIrKQfatIvBStwgESZOLFGCkCujVpPgKAkQxvai0BGad54mMouADJ6CLIPsFPD6ASK04
HrLFA0Yqpo/PsDjz7u/zvVjpDVTqx+tMOVoPJy/H371OhhD84GPDH6lz6MJdA57ckanUwQOCYri9
AJJ39Yv5/uyyTQt7Pi0np+QNbenFFfVt7FYSJxtYBw9LkJnz/btuwPyVCYbBAqds+MgposlfUOeD
z1PxBu7zbj1nzuNIm+JoEU/ufvT7q/f6OG/SdtwmcRdWFQOsbYbM1zA2QKMbJfkjzrxXscYtoxop
h8Fp1bfSIER0dxVXOQzlL25JsKlOziN+v4pHfgGfgaUKFpnux1e6Zsbq/mS6TI4J6NlN22jhpw5I
DSoK50W9U+rTj6XXWOnBQjGkMbsGkipM8d0vYH0RRwg1IiG/m8KKigiCliM+TF3Z6aPh1XU4LvcN
zyRuzAT0JI99Nzs0hNT0f/ScA4S6AkIGReyetBDeAGA2CjZjwV1cjScvYYD/LlBYYsjTUNWh39O0
/GoLXESGoMaVfY9BcOpROdZwlv8MZg7sZ7f+M7NQk8LqQnJn0uoP9G2uENsMdZU9K7aByy2fNA2U
6BfEwh5TM/lGV/kd8duUr61SNSk2DPPTnp9wPugEamag+QLCx0ujYR+D13e2E0tu1iZuwLpJbsjo
lL2Q2vZicPW00xcnpamRR8jBeGBnZCYT7jFZc/UEAQN6QvweUi68wRZlofdzLeuL8ZRlfQZ/KURJ
rA99y1M3rW23AiAoJPHvuzKk3/QY7gOcyUPoEYfT2c+Amqw24h2ZMO9xGzWpSsr2N+Knt6E9mBj/
nDZIGpla3LXxVoIr6roA4JWP9nRcxYYXWzR2J1L/8YVjLpF8/Mvn8JGRYqaRRHhyK7xInTFhhvcN
oWd3AaV3kG+h7sj7R92B3ATg55ZFFgOTWXo4HP8aou5N/Hoo0a/WXRFiRYQSSLx0ewhdp4C/yziA
mKDKSTucEceX4wSh4/bimo2i8kcVzaZVgmABjkjexUui7nMcJJWEfEo1lXMXBO/64DcimGJN/gk1
uSPNpjfNw96ShWDO9RLwRC+FKU5jY5N5EXG8AaWl2Q8KrHRb22zzUXgnmNyyck/7BwG4gwixkJAW
6IeAcrpDHA1YpbxzqV8IhZ1Cj5z3z1BGaxfBqYYgXgzzw0VlH3aHh0ysQ8SLR04XCAzaHFA55AXe
ko32FShOWCtFmkTP3txjbaXm3CABZ+vgXSEx++8HP5Pkui1ZffUL0vpgHoDHS0XiRO3najVGRULP
tlS7ce5tm4cwHwal6LHcTj3XgwjNZZt4MEQo4XitSCjSuOdS0v65JnP/HHHTRfKrCsOcqG2ur8+A
Mor58Co9J5iDhIydX3g3aSVWq2LlbAMURcQYl7Lj1avNHsOwF9N6DF0JRYiwIjM2SDnaEdygI8PK
Nfc3NH9oHBdlll4IKOdI3ktG8xeqqxW2ZP4byBZi1Qg/ln1bLmZwDse9JhunJhWEPIAlbRyH44Au
XU3EZlAd2uD21tfruyuo41szSq22owXkbmCpJhI8gFcYvRbfxwJuZ6upTmszkyKdN80rggxV1Rly
Gr5ME6OPCboqmnJAKu7YlUeB4eY9Ui4tFY2aLDADyouY6+U0U6RriYheAFoHuFILCgIYsUav1kSX
iwwkeLxq9EjEMQu3VgWL+nJ5He55ud9H1iv5vMDAboYNcpMCNMh7Rf9kXf82ZfuXdY4qHOIBcUVF
1DTvqa/IUvXgAFMwlD4x//MNiIUZrlq1BA/7+kVyeKFobe4TacaZwe8Kb60aYa7tcKxQktghGNhk
gNvORMhCZO9KL7+O6YByiPNDMImKCzle3cB/PVvu76xH+FnpQITsbSV6T80d5NriM/aKYMy291u0
zyVFzOPiKD/v1F9jIFrvnJ9wAUsvj0nLwlNuJW5C/9C5HCu+RZoZYnvYcZxJJ14J2dXPjj0MIjdw
artxQOum6XpggFxwyjtMkG2wwUuZNo06YZJ8fMThlKZT7odakwyk9KpMmuslu3pj9sys/s49qIgH
AVScVzT5Oxf023b1g4ddxeKGlBxHtutftAGITWBjCru6+8CJjhSi+spK/iw7fsJzCtNrJ38jMXqC
DrSp+QP8/RvUr8HwcwrRAuNxO4KzLsVqwFkLIOch2oALZ2wJX9+PSyfLRK7VJPBuJXEB/PHKYtxn
9cZov7fxSPdet2ew5eXNI7ZrnqRFyrBbeye3apfJBoYg/wlzqkbeZN0FHskHJL5eTo1qYeNr5kF8
Mkf97bFngY41wcLOnjhHr16zCe3MPHEO3jnfuEnW+FWLOXxMl1t3WBuG3+HhbYC5B7eTIGdic70Z
kmzFcAdDvN/pQwZjQMB+hM4e6N2WYBbhMZ4Fp8xoNTkluhIGJf3erbTLnRksUIuA8hRhheSjNIRr
jeh5i6hcsTKzuN08fdQMLHhKrKHAnKxpRvPTalvBUxDack1TKeptSOTiVu6Twhk3Kgrap/3/qRPv
D782iD666dp5WgOKKIdi3N+YrA0Mo/iZPcV88i9tlLxLR3t6YkoUpMVFEgwa5aI/SzU050laeM2P
m7PxPUBN5uZwkxdBB7o+UOqxOu3nJWEnaXn6hSaR1+f/+CZCXPZYRoyMUtlsveF6eknP7+P1amy5
SAV5Q0utK+bZg3r+UoVc9k0qKuUJWuD7lyOroSE96PserEXfLkTgnRpEKlej9xXXqQPubiT81Zqq
dsMnvkDMkNHUaP2UOHmvkhcBDDn3PhdTh+F7uCgxVyKEFOVv2ZuGz0XWT5xBmJunXvvYRin1jIGC
YZO5qZ+FaugtjGiAMkmCgexK/N9WF0aOJVfMopnz0jYh4JcdN+1h+xitSFJijuZkOdv6rBwGE5Hs
GKQWA6Osx9Z6/hRCogVR+217xnq7iaeYBTTwe8RwAo8MWOcTp7aRPCx3FSYoc30CUiLm3Abzle6A
Wd17UyjSlB1VpA8iVX1kiggdJIwsxp1M3hnmoeQJ5t99cI9DdTR9bCXLY2zekdS7LceVvQG29OYP
UkEMYKw9bFkjDMc/fDYFiwupABeh6wGY2qa2s+u9FUf1u+15egT6IDb3HAZuVeKoy/GbWzSgney2
DlRkdUzXKfEWgAnhlFtvTtnRM8tSli39x28IovxRa1nwYvFsT6aKmG/Vey7WOZ/gqowMLYki2khu
THdzJr7XEqxMaTkae9NlREubbG4vlfgZf+/gVMe/nk+Eo0fMndl1n+Lei4W+N6VhRHkIvx9+tGpl
OUWv8lPUGz+mzvPbhsJT5D/Fxqe4Hbj+4J9li+ChvpMbSV3V1ZyLoghNYcbTwPlGTioBeiQTgUo/
uXtRirw5EpLCz4f6tKwauEcicwCuQ/ASj6URdupjOlvVJr9rFS+5jV6hZuFIX1pbwSXq4GM5RQvj
D444N3Gyom/DmfTQc3ron7Mta3E9eqtPLFF4XnfAG5ww4WAmSEkd+KNVaNfItvENkDwR8BtY+JdQ
YxcADnmG2BCyGThSxwpQyKx7OXad1C2tpsldb5XN7nZQXzaoMuwxXUEfZIx0euVCnp0pf8TKMpTk
zslsqai0JIMTJgdUlwZ+o3y9/P3q8W3sUNkVC9RGsWX6VsQG7xzfwFdsYVZoor32/0ORO9fldSTc
U/f1ZFHF5bh/yGfrPi6n9nU/Nc0wtn4DpYq+QdS8rLFOB/sc/DYIZV7jcEZ2YoKaW4L+hGlD7783
R1+RBbi7NO/0rFkEkuJ4rIBck6m6rUNdtAxjAaEWjcRylvKzbPUrq24qWG/tb+kmQHE+oF/J396y
+hEeyiaWy55UbLk7ZwbS9d+KitVSFowmmjl+ehXX8rgFAQSOjTE4IePZ3/bVVjvGjQsXwXh+qT0/
wtFb16hk52L774bGRkI6LukjLYV4LbIY3gvwFnSb6+GdNXWLbOtJY7UIqOxZDr0y2Pu1W19fmISg
Jf+CPZZJrb2lB1VyZ+ORhwUD4OP//hAUXAW6W3b55G+ILy6jz7BALz2muIWBHtrQoJgiC1o7cN1S
b99G0SzF3u0p2IVEQJ4Tz4IWiG2YkB2l+NKM7eLkrDBpLsz/A1PoWLOyY4zT/+xc/j4eHazPzX+s
0ZScYaYvMBn8zcJVPPYOZ5HCh9X0sGa7hxMUNIN+MSuK71rlWJi9D9chqg2cCw2svlTwnRvBM+e0
HOlpETwNvUxwevu1aSCMeLqewKCtUSmIkA2jlmbxLOATzmGYqcs/uD6bpbt8Mdn7pw1ajT+7wc4z
JnkNrbV0kqRrNeU2iOZaVNpwl8h4UxurdF49XOVKs4+40DbcIEwDo/3Ut8idMpfZr5EHGxIIPdi2
G45EPOJ8iTdyzYDKPynudDyAI6AzfUKg0fE7NPncP9U8VI4sek0wX+f8AqB+0PB84U65YnIJwTAH
5ga8u+iOdVfyCQw7z0qe2cgfmkIWpM9PBlJ6i7mYkVLpyDilhjNMEOymSb/4hYzBfwnKT6HcGW00
XF3eLxf3BnbsAK4OnxojtJGV6iHHe0ho//JEV0Umnj1fxD6j9EPksNOrRGQRiOkXK/VNeN5Aanme
W4gu+/okRp/9Vt1tc5OLI3aykoCzVePLPbvdKd8pNy/WJaOyBea78GRS+KpWY+DYRF+wN7wC5VA2
h0+rqvnvrTWDbk5v9Z+tPq5j0+iVt0ja0tINXn7KHtOyPYMDBpX0nO0I5oaTTTP/06WWXq4BZiLb
erF9VzDKL5vENK6iv8cCKEe8g9SMP3Jxf9jzBSBypfdZ6fOYo4auebDmZ5kN5kQ/7KyIWEgNVt5U
thxrFJkkt134IHdsyv5CY/Behp1dosfsFdj3qq3RfDwoDFvt1wBLxw2N/VddkVMXPDcWbL0CcXfw
y3SWlWxZky0QTS4zI1Z51ICSVWaE3mN6eK7SsgUNkdvtPwuofD2ZU+qYkuNmb7x9cSAOZpnD3N77
EB/GpWw3i4yxgAJrFiTxrW3O5oVc2/xJas+SBekOHy31KSIKmIWRCvXacVzeTUW5i7DZVTfNkb8e
eQc0jTQWZo9KPilOrUzNBYzXPWIFyCtS3NW/w3JlQlhCO1nYJTEq5ZOJmlhla/Yd+JmjvChuuYYQ
jMtOVPnSdlY0+xEoYyeNuuCBS3XTw0Hfr+jHjNWgjNxQGgdhSAu0q++R0AHF9F1zgWGYEbFzC0R2
kWipk8d3r22yhC7VHdWajil00XB8v4335bw0/ALeWB9kL6hPFRxHfeqnIkucRWZkxWoEiUPeNBp+
eTX7WtCE7hmJ0u0oT4DtrurNOZBavp/OH0zPRopsfZnWl3NgFdXQq7E/7pSTH9CUFWnDhPM+0V2M
oc3bUQw1PuXp+PNV4GlJRe/s/2Az///acPvC6KwP+LrbVL6o/USNCnNWd2scsPbTaLpCbMHa+Zx4
ToGHGVONTorPKlfVyMIxluk1+Y1mzzg46UNoKlDQ3fsaH5j2fNn23pidvPDz1njAVmOmrIziqE8n
KaEBS97m5gXbMQByCbNEHbswYGjTpDZ46jUtWe78VqQ9uZnY19DUNtop9u4P2t26MOhUSWwlAc14
rTZxiWwis3HxGaToMC870ObdWkUsZZXKqWl+y+xGjPNYAQVNau/5ufBIsZobvZAaNfPRqwxK2eBJ
Duf+gHu3G6BGbfmYFGV/ngWM6o7OZhkl0hHgZVB4aXHkHpy/wQh4lp91rh9sxoBMeBev1/0r7Z0p
DdPTTVViG76gLluWKHZy5uglxng1dRbk3w+ui0h64OAdKE/zKRlTaDJY/Nmt24BHKHPuWNtWsY00
cokyr+Dn1LuX/UyiugCk7XT/YXNejiAqNSkAOWGWWlh8AN5v4ZvDzhPusA8BWU1HxbAe+EhZRvxr
uiGrjolC5Bp/l3H1ByOEAqmiS8mrR7YfJ4tB6lwOpiqHD/0PPHVpJ8wJlsOwD9l4HfH7+/lveIa6
FdBvTxE2GLznqYF8RlapL5vVRVeJtetOAT6c5ByZ9/iyib4LIZl4dEC65C7nMqwZFkCFXcnKH+JG
MY+o6/M3YZIwzM/k5myVsSlt4UGruSC/Hj//38yM6l11K7ahatzvL9URtabj0Jub59SBLTeHRwTu
Mnh+JB4/xi5jDSgzdz8haiN5uAf/fYjGgRgkxC7tGxTTSFU/k9/1A8Bd0NHL+iqHXAkDPaNb/r4l
1Py5hfy0IKnl+2x0RND3ZXQVtJs3OTSg0LqQIVDNRSAvfBft50MYXXX2KJbMoqT5SCFXO2Dlh9ZJ
fBZV4KHcvgWkoDARvoep5+ZCwHPlPd8wE7qmLiUlHFacoCGqGfDcf0Nz16htgreBTBTPUO1ghF4f
WuAjjBmbp2ZgpBUHdhu8Dtb2b0cgO0fwaeSUTdOeMSBCXldQ32IJzljP1Iy98txlKjrxsg5p9mO3
5tGH+sCOxAAaxEtm/oZDPg5Be+1ZtRH9WKdOxPHZPy9mFgaQl4cwbVKQw6b3F+LMbyIvGnRP55pz
OBO9bBd5bPvvDaq8DmQmGzRduxi4yp/9lgZPS44imFUoxeI70AiRFu+ZgRTJASUrgUT7zq9vJRQ8
IJ45dofliIZBOTpoPeQVjK3RaoO6aS5s29yrb/JgiUsCqPrFFSojxCUZtoMaeq6J94tXCK06GoKa
bQC0ubRG7+cXesFvfeh1L+5RpRtQNCCqz/SI10nKDqkLG5G8q6E564VoXeyJ+I1boByDq5BT80UD
W9y4s/9ZQS7p5mq774NxlwP9HgiZTO2skYd0pXIEqyFa/4y0W/FxLjqTx0fsMJV9if8eEdNf/GNw
ZKF62WGfNeWJ89uQT0okPQtCGyHqkIzrmbxA2XrmIuwV9kbftpJ/RV8WORLt5bDm0hznEIgSj/0a
+DGiVJAMkokOQ/65HwFB2bkakfj4glc3LeyBzjB30ZeArAKNlDSDWJ+Y/sUkGFX0PZoeTgT57apa
ZP2boZUdWA12RzpJZM7V/4tgQDaAhzzTT0P7BYMwL2yR08hz6Fz7KT2ZE7MsZFqRpQXHpUiH0VH+
Kljp+vH1vGsK4rqO7OEb8OKMY/L1t/goqk5v+bRRYYAT7DCX+Is3BA3chAtfwj9BGpRF9AGJ1/cE
AOBifwrKWVU7AboWr8y4XqEG6Fb1zpWGknw0py+dh5P8T0heDbBILe9wtRHkGami8p3GeLJL2SIS
l4j/SxQR3b8KZc9ni7siVj0SP4XQxppzgR28O8ztgOoE/0bq+uuNdBUVKTfkStNX8tG/iB3J8ZiZ
loyAJGq8R/oCcUL0I2KpgSkxKhmNU19Xgfeni/p3ohTD5n240c06RwDaDKNHLvFWcxKupnyEsCGB
9aezo50VHd8maaf9Yj4WyoZgCnJowOizg50AbR3rAxTVaQECzvhQHAYfL2VTwnH2rn75XCl2VxmH
f0nAwH3DinXzUrxCmSRmIDB++PK47geXVU2OIDXoKtL3AbXka8QEZTJsZaJRQTu3b6Y7k7DJmDvU
sSu3WIzovRdAN5TZ/FyAs8Lwl79RYGI5ofX9fbXpmeDCeAPEAsdZWeaHLx3S6AYnNbnuA8Qz2Tbt
2BVUFL/bxoJuSDEYB0AYi+SJofhvpKVL68NLvPW+tsskkFxdUpE3tR3zEQL9BL5Pv6Jdf5c1XX7N
i0R2CdvSBWMSDM/sYXZceiTUY8bGsfD7CMzDXyI7qpXm2zCGAYyF+RB9hcMlIZB42mJldlvuQLyD
770xS+ra5CkRjjQ0S+4t0UvRxTKmO2ijsCrlitoZR4DwWcMBk2v08/ODWfdkveMZKiIZ7bxMUNxG
QNor1eYFwgga7HhcMFCh3rPzIfBecUR7Jm/9u5plkb5b+8Io+uc8EaXpph8ahtORoYgqFHu9wHCs
gsFUTsWYLQ08UcfYZlZ18tbmXk5ogGL7FK0xhU3zhy/L1KmjgIYvOwOhw787ScD4fVyfVrJIWFAF
ZW3/lyUwBxX9BR5fy9sYEur2D3ebj1Q3dubhGKIm5gH6DoZogFjHfapNB69SGen/6QdEdSNTLpYs
HoMRAew/UWjgUzNo9ST+Hnl1hRkP9ifiFMZJPgaZ6BmSLZUaHpboq9pyvMlfqwgqR7TXSFnZgeS7
OAwDLwFOH89Lp7E8Vd0tPvp8DlA50M1129rTqjHKzFitjD+1f/ZBb9KpcE7AEG7xvrsyWvao8eVw
REzb5rmef1xVP26YhTNvjlkURko2Ub1wlLiOsqXkbiamS/U+yL/XK86ssL0Q3BQARnXyu8ZJgfNS
Zk4r7zLyxgZgT3HU6MOEcG+2+75+wlr9hDwUJonTUGvsygwXcbTyppHwiXB3Y1FdjYxmfbQmDIpu
wHCzAVHWzxb5XLI6rOWPwCiwg5/VgYm511Bhz/8BSr5NjCavQPSFTmg1eSGb/jree8JhaPu4ppo7
4bjJxvLFCL27YNKTAP4vyUX3xHEgC2z1gifr7O+KgRFtUJAF9VrSfQc5BVlJA7Ywnp3wtQOPICzx
WnZqYXw6/xb9y52PIV0lhZSf3Ws6UBTSlgfv2kxMjR+H2AO47dqvG/4VZSLF21NrFAKpGnylfyT4
4LX3JCNZOGn1zQgIYrXRXMqNzvobLoaJnTWWi0scgIo2BdTeCJm7tkTfCR5PCHLP9be4jfOz3Dia
NjLrfokYgEmvqw3rNDkM4BmIraqa37KsMuz6uTaQ2uAxRKO7vTNt+8ifwktOr7mdrd92nn4yQgld
B6ymvZnVhafnfeOGlJjNY8FrpkkkfDg7l3mUrUXzaKhQEnCLMr2W2xHwFp5H6CG3VYjWmfpahx/R
2FM0TKIQdAIVOkls+Zs3Pz9PKMb0EPuPSK6OVsnxQhv7fwpWoTcntOwrk5IMRrkGbE6sbyPrKmOp
YLt9b8H0c78J3Yc+h4HxGVHdMg1HHprIM7PHLUFLPP4eIvGc40qU/wpDx0r+2tWutJpr8PtxPIT5
9ANbJxLCVy3FbyyiUfmDYmB6W6Infv7w4XqvnHl+nmC/HNPLOvPHNG+obUzsZtScNR+JkKFv5TmR
Ypn24UhcjrBADZqCKbNjhCvyB49Px2BHdtNIcG4+KoIk+96OhlltiLKRNFKnSFUrPd6n/M2CoeM7
YmlezExneQswmn5b+DvUe3f9ZkCepmXfkZhao79Kd7LiJZG0nEt6ENwkhp4ayDVfYO/IVw4aluBJ
kxxKb6s1HeZoupcGYg/3LOko/2kVNcFE3mXKECg17y5/CfFBkT14+81esWFPs/b3QMbZGw+0u8Pt
BVbNEFhdn7ySJtvJiALs7TrjMxVLmxsKPH2CbV7r03nIcUtEqgHQwzGZOd7O33FDTNfrLn0KMsO7
e9+N86E3ZcYq3eJk6i+CxU8Ar6l3M9lrSM3oUTerOuZietQ0sA5McI8RFowsrOrwngbzN3JEjVfD
ufkkb+DCKMcHWoFsCkAScyUrZidqMApsJ5cryLtlvyrI4GAU3dZgJjswQcbZ2G0lDowaamulfwx7
ZwbfGIip0rJi+F0IzLd6eZpvvpl4aCl0xqqDZevuihWaWyHtPLeXMW48JrujtM0jO0LnW4gXlcUX
krRzI879zE47UbcJhZ/G6dOyFbyHXx2mg26Ybzj17N+MMBRa4hXFM9NBnO/WmQxCNdKnIcHTkmAk
GyRJqNtGjglTkkXxib/+O6NjOK1M3FMPpdMpA7TZCExNtAGXLgS07RPPAsc9BKbL+mIDYIWjEP5Q
iwS3GYHPoPyN7zTPVwGX0mHV+le4VoTU35P7sVz+kA9ZcrXpjG86uMJuc7DQap0iumGcaxKYeAC9
2QY4oEunZ/iwJfDiKnXV2IB5+O8jQ4ZKCi2FaJSkPgNOvvS+pZdnRZapmxc+iYRUZMWzngk0IceY
clW84fuyfq20AnlBbH8LpPIoyEr1ZubhlyBhF2JDCJI0QUDPa+P6SV3vvzFRmCMCVfkXPhTbpViJ
1Qa4Xce+zmGcSvfxcs7QrmVUt1R+X9RAP74B7/uHhVfv3GZXqkMdhD3MWUIvPPNTmnwWQOTeLn0t
0fXZLEIed8Xme1uKYOR47izP1Hg3MotcJ2KivX/6S6EYRWPuKcZSL50iYUEet6TWKB4+wrl7v/vx
rU88gQD9lRdGx6dsJAih61WolK+xvuGIy61oR/DJYqSFTh078mTzEMN6W5n2nkdfFs5gRvq08bWm
8dWdplV2qT5PR3JdD5y3Cqh1/kjxBHQA6PYQKVoJ/6nwkHjIZe8mINQ+jUsdK5BCO+P0bkL7KoFe
gF9eaJ3OkMBLIArrX6r5yzyecgUChen7yVGdVU5wRP0KwX6AWx7M55xFmN9lwZ7Cyz8ije+dYF3s
RVxPTYXzW/gp8zw2bNS0oWnt37di6H/fVAQV9R0d9fp8YlysV6Ep1OmcvsMGlq0WMpWmW3Vovg7q
JMiZhQ+c/M31Op2m0oOBTcYRkwUX+Y6/+6k6u6imDGB6wJP597MXyNEybECfdcU4HHKguxy8THQV
WWicyErO6PSf2CQEXDjVC4ZQlo2WrkyTvF4wAorofBG4HeiwY959wLGW8gGHJTkup7lxazTCHaYl
53ch/mtLDNBOH9+7wVWYlNr78s1oTT7SAB8B8OGsgwmUcBb6bnVU1EKVn3HkDZOSsILwkBsNfhQ1
dkiZCREyw18WHfoUO7KW0stoBWX9S/rcp5BzI444zQkMfRAvw8js9YJv1NCUCcPInhocFYAnb4rA
qCm246rIqj9jliEK6ThTzjkfXS56FOqnhMCaiWAjjgHqJVZ8HIXdYAsvN7wtJyG3UQ3TcXfrZZV9
/C4zSbGRpyJzLlcwbE+gxbv2DRchjkFh20j5PDrGkJ4ADEEXt/14r0Riw+gKVrKS6VC+jHAisTqK
6TaYU4iYOwzUXxoJ34aifqclTPaczej9D6ZYRy3dMrq4LRisLq2Zp59kFWXxOW2tjdlGtB0aczqP
13DQ1VtERqMK+5/deLRNEWGGVhux6Xlxe7gBSFDbgXqIk+EzBh1UIKhCzEshQgJYE7zVje3wRaqh
aRoQYPbssEVZETNwj+J7xxA8wH2vkcTHTAMCZKnjjnXjZp4kaVxbH5o7PueoM68TXR/lH+5viIrg
yptmIbz7LJHFtbQfy2E7hYk5+blvQ78hdwJ3ba1bUWo6RsVfUz8uyOgUbednjfICRZrXc3vVWR0G
GVtZ+2nsc7z5y79irJOD3CJCPZlvqyw6VS/BdHHHpoY6Up7OJpw6Ok1ynKbm21KALg2KYs89NNL4
7813r/1sgmlp5pL00uvLaznkvli1QeHn1SHpBu501LW3R04mCevc+5VLIV8/5BDOJ37rAs9y8ROF
Djzyuom8Fi0O0RR8+tYSI0CWFVHrixQ8VTSdHtDVyBzVVJ0NRuQ0IfRwqhsA7w3pTAwCUwN8FjIY
qxtc4//BGG9nD2S9VwYSyTy5RyQXWUgqnVKiQXZT8Hy4VMPV97ntaYMdX9P6qSj/YWaFmh3pbDL7
Ynil7DZYIdwMZ/8Iaq5fo2Vx/EOoKp80loz0eeVwDdUaSvgbOCWD2VMB5Q58eAyzHUdwpQX86gme
D7L9kSM4ZK1H+B5/Ugj6rBNrDh4QmTiQtUfhIKSvl6cHvLMRX4p3ZdPUTm4xk/2epy+BXrVOOSyc
gryeS+wFQgWv6/6/W4PUcpTJSMcxAVb3oVKoMwpZHEKTJCJ1yBsNyKO5ADo9udpvUQv8Hd7cUMVe
XIrG//yMYUodrAUlBFA8pAIAjsCiMWoizVteIffxn+ytLIw3iP/WXSPbXyKm9HgsidiSSulDfCuf
7bWkybIfoSzeWxm5DlHZzZivVjyllzrTtMzN1Hwz6lu+xaqtqZyYsgL8tzKalSFjoM+OdvgIsPdi
JCbU2WJ4mo4zXXSeRd+T5wScNjxyQqowCTdaf/XE+mZ6/AX1DUaM7GWxKBkM3sU/F43XCXSgtmfr
hvKjj7AQXhmqcV8pcgATx46W40nNQOJXB0D6GWfeJKv2bIheVbts7yvOpm8+Vo/vdtFpn0khl7QH
++jKgW7O1+xF37RQE7a4AeYjTKGGZWSToVJSA1XtJtHvUAyD996GauCo4Nu8EN2mkl/0Ulw7h4kH
vQNUuAY0/IDZwsZhjc1Q9UXcwOSmT6e+GQwZetr+3JWKvd2LFGPR88kxSkfQTSBVTHeHgsK3POcU
W/XAPcskIt/0HNKXt7K2BfS1h3jd09AwPVwRDLI8XpFdQnzCxQwXK3u4HAOrjEnWsQ5MVHWc+Mfy
/QUIVUCOCUeE80bbs5BSZEwWOmejlP+sbQhiyvPwWeWrOqgBAHZS2XbXOnvPRIirGTJHymSglcIL
IV2P3nqifgX3Elkc3HgutKftX6A8jztPDKRk+uJCy4GZM7cvJMhvmZLERIvP7osxD3IWC57Jjqxc
ky+OFy1lHEJP70CpYLpeKmLQLg41PoYZ2xvfo5Bc1S6f6ZPcjTv+fQZysWRr8aEC9t83yZ/JZE28
GHs7xkUGgx1YeKz/lPoQOg/E+MzKZ00uY1pVs8ZNY+y78gam7Prt4G+qjFycyhi7XFq2/lrwv2pe
Ah20PtPbGEmTuqQ3vsp62XaFJ5RouPcZ8WlSSfh8eywiSyPSZ8lA42O+eqQrzQeAL9dfX8QTmCv4
JjfXlJ760txgq12TFa7B9jVeVmayNtCeuTDL/DuGvhkE4EjRCnUMWnwibbO+mBMVUPsKbcfykAY4
Jvw2AZwUeHy0e8yK5tuhD0IvlAHmRhE4aHkgIi3srySHlWsWgOzMRicIhbEE1Fkpqwhq1J+z6FEv
pRvP+1VQwweyqc/84eBZmyhwjfZAAZxEtYAxb1HPMnYPQeEsDZkm9QXRMoRN4VIVrovDCcITj7Mz
9usbFk3wGrau6cwaEdjgiinp1/hPgUS81QeLBVuU4xu+2sVMt7VfrATMHSxt7bH9u0RRocP5zd6M
kp1IXB1IC3LE3rdc1jb+I60AIPkfqDAz91ONRfiMjoPTAjxt5JwFpPUfXwYLYdBXODQN08WVYmDf
W16KbavJ8ded+2J4wgH8XpHEn+ccrJMrVS9oAXkUEAL11XMsbTfluQJgVc+I8e1+qm0LQ0cE1ipm
X6aMWCQlzrvWF5ccaUz3ovjpfWE0AEBdU7ncXzExN33bCZT9DGJ/1Qt1LZi/rlijWRduOa+T5sMH
xl4KtGyxIu9bMBGjWHV8jJX0x93lL3/4AioY0mx9EZ7vRixtxIli6JHPG9rjnZiuJj+cVmZmHb82
edlRq9YKH8OZip1Jsnd1grcXDSSlUTI3434QuCdTIirop6XOeuzgY8W0U+TxGADx4VkQOXNl01L0
B4tzxKtNFI+Mr46vY89FuM54mta1pm2TCpJ/Wp2NpTVkbsdaPWEPiH3jgir8TaJ+l+fWUF1ytwWG
0QQ0OJLNDdXJGGR7I7grpsks/euVyzUpqEhi1U7VAKYfUH/2qVCVmJfr/eS2pzOot92Jlrl+Tfjo
Hj9gORtmogLL0ovtu+UE9U1lFKV6VSY88jgI0nZ510LGc4ofvkBat9C9YiWHmYz30e/OcJU2+siD
iEdiYu6lbZu8eR99kJmOzDaGFpGDMej5qNJ1rWkNJiuo+7Vyxa4LZL47RIFOcgC5XoU6WZdX3VW7
2zh6u9redN/FlxYIYyfcRkF1O+cGEAkXNSltkUYs0poHlGYfnblIYLMjgjDkn4RjbUzXhPdvFJ84
qgho6n4gOUUJXkE0jWTKWnJzTTWwjPaU8AOhN/4Vo5uDHsSS5+7Y91np5mjcK2/Pms71nwY/F1cm
ZCWA24frgD1cgsYEGjFwIF7OFPj56vKDd1e/AOxk91PTAz9NBxhFiKdDDX1Y983lgl4Nw6C1Ig5n
T/TQMOv4CUZ6mURHs3GV9QBvFSjfgIpV7Qdz0GcfzhZHiMLteXSruyesJZ5byHn5OuErYEIniUbP
3Hd3KFAfgHRVm770uzlvvhqM3i82H/VMr287GypcyzjLGfzxY81DWD4tPQ73IvPRFPNaqd6mXYin
xMHPzNbLqBz51/ZiClZun+3rGnVmTJDZqnjh8qhgPBgPasKRC9QucqJmkDqYBEJh83fq51Zwvx5o
W3iW4uyJB5NHvNibMME8qkImoNCuJRh7sA9wKWx0EYpmWGkIjkhr+5Phoc167/kbXkWt0D1cXTA6
HuJ9gDzYa+uHH5EpHByLlDaZ5qm/ixRxO7Sv8LnDAtzOOMSBu9SSqlsH+jWU97pRp9PR+Ybxmtf9
Uytg10qtcSUyhMhKfWbntfTrncUYlDB1/wm0Fu1h/Xp/u+7MInPeEt0tB6MDhvzScdNm71e7LGzh
dC+H7p+IwqJiFVKjdyplz7RBdNkCvP0LMDZUjSKwPFGbPUfyUIzqA9uw7KvCCk5bnl8WOHFhy6eG
4NCAoD0O5sXiN0qPK0nO7Q+beokOCmU0rwhyvTF6oi0PQCCOLU/i9IQOgfl3/HtCVXPZ4A96WSmG
k6py6oMyRNpY85/fZw6L+2qNsO0cmKSRz8onEP0r6/kEyyh2WcsZ1m+Qx9Df/+cACV4I9TH157AV
ynoCWQh4xoW09wK7ED2P+G5q8p2MQaeB+jpRYx0/0DLhrjJl/lrPDn4sSe2zIjp68W2gaGGbOvSH
aHW7Yh/jvO55wg+8/Lw1DCskNsxpRYChzBwdB7rLUptQI8qZs8hpnKhyyHMJrbijx3zRdrT4OQ45
tvxc3ZGtlUGinBYxGaYMHAo8WrvT8wfAA/m8XBbb6k3sgzdPwri97rH6dUbY5vxC9g1lieINWjIw
eEYU5fZgTKSb6FvuFVIViMfYJ3ns/M1s/5j2xFPCV2pOwhkGv3UHNYpNdU/j/XrKi0KmUNpCaILI
Zsi0g59oeP6qoPhacrHqtVba1Bcxod7DJ4ZEfCODWzuhhfz/Ah4ksSZdjCmxkIEBSPLrbQISS5mM
H8PipgMEIsPNQjf5vB3VkqvrXcuGRIM9AcIEqfcJGc3v7QKgIc5f2ErMreHfxx7S62YjIoaKRjzR
vO8EF2FyFS2m5UNkb37T6xFFNls9mc2OnTFlycWIfs3lmCEzV6/xRLrML5r1zvj6FRK8S4XLfvUZ
RcQKIyR3VQpoqhAPjzDbcBrJFmFfjbCkaRSyzwN0O2FxLyJrqrARSsXFgl0HbRJOUKY0BoFGNavB
OiMZB1J0IqSxhTdixDi9NeotdfHDgyzkdiYrdWZiZzr+lVF6xTQdCH+YCqGgQzzV4jmL6GiCVFyz
nm8+jNwHQKYD4OSFJXbUYOMBMQ40NJqfYQhjcBDUr0xV4ywoUKrUslONOsGkt38mA7mefiue2unb
yKT5A0caDPzl3LQsk0MMluiEhYzO+GBo8cJYffgorrmaJoZu2x+k8O8gDwu7ME+EHYZyJAFvAv2F
daiCXQwiartxlHTfCzaBg4ogHhhLgm3sZgfCgN+yvXgojc33NbBsW9kYJO8l7InIQWYy3yhVWlYn
0hVYuB1p0z3mJROl4a5KC5tsNobuE1RPgkYuCpjF6cEAB+6Ss/LMGYhPaB2NRbRO7RC7KI4nBEy5
cknZsdCMpGYxZBZ55TBxU2jvgaIhHojyWsid6RYPdX09L9gu7STdFzRXL5n+H0XvD65+mZ7Ncp+d
CPGgs651V+Zr6c0X0phlj2boMG8/eb2ThWlNkOjiAeTJdbB+FIERN+NvRb1OChp5JkUCrpqdA1TW
cKjhucvZWCLI++yCRBjTp8doIAW2y0jyN/JNE4naHBf4UvhOf3l+r9YQc5iSXzs3aig0DGkxxIZV
qM9ncMfmKaRrYK7SZuj87cBLyMKInNGo9jifGsNQDLtK2cw3AUpu1h70fgE0gNBc2F7zKOwYoBfK
gwsqYk/KQPKxK30ikGzsV5sTDB1SUvtToqP1o7yu7karp8zIja58l1qO3xIdNzhGTm5W8sZ2q49I
k8Ho9ONn77+Z7V5tb5QEOmgwDgVd4/TALfiAW6qRDctfS9zTDxP2CrxXnpt9wE6+Mn3PrgDfQ4zM
9Cu687f+aaBR2rcSjZmsLqn4FZDB4pDayxVJ85rErLRq1wFMM26hs7hL2dSTGfSDlyAjB73WWUv2
E46UWJM2BMWTRJtfJ6PWwlbXSy6rhEeuuMi5FmnLEuNLhNPm1wr9fhYNVSRz+VNQN+s+omDN5z9v
BD7woo0Vxf2j+FkqmhNFrhjIUJ1vCrNw9sdg+9WkpXd3LGumfWuuTztw7bNQ6Q4kzIF/oVes33P/
z1S+JPNwtaz77jiqHceKVLs1Vxk4M/GMwB6fGj7ROBaQDI/BosYxLigSFqrgDtI94BRiqQVigMdw
UN3hgzsWzWivMe4+bbCFl7UYLlAVuNSwRUs/FNxzttYeKsrrz06QwTM74EzQK31Ir1BK149h+/UE
BBBgnUdsFDYDMHOgwHUxrCq6JJmK28t6Y0dd0SvIM8sWjEduA9txQ9CkGgBz4yVeRhnkFxw/Lp6s
FC44CosYBHMqT51MH4soMuhJbC+2jxe/lGKq/rKAJzpH/5qO2vEp7iooHDBDs4XvJSXW4JFhrcft
frpHRYuyKNuWul4uBRsomHpVHmt5J31OwTlLndld9F9i+Oul+GCdj9RvWBAWW4blKGEBLbkZWtQR
wPq+URUA2cObGWDMiggVkDD53KYLU0PJNYel0Oy7PSNoK3/BKNeys8nBdU0Wx/55/njQu5zgsju9
YLPlCxWYsyAfWtaKQXz2ERRl48INqQ9dEFAtkU3QTZhe6YVGUPETwKptqXj739vwg/8GzsvGnau6
F18LLapDmbpvAquuxFDH5VI1YqAgBTRq0xq5ToDrrYx4DVo956RbEO9qIuCRWoX86krhKv1Edtne
ACW9Re9vsjdTKR7Kz0HasruXIQPvZKQmbRVwWSlBFWVGN83yTI/Y79bcSZSPaOXCS0F+7YDgMMjM
3L+2ULWYqTSUDkhiHoEnLttkx7xuwU/DX63kZYpC26Ba2jEMO91Q2ctheRVMyCTSiqBHiVZkYDl2
NY4lNc7Ojt4vXlzI6WZDtWCSbBDeqduDL91V6Ao+xOOcJLX92L23nJ6imjVnlNcSKPlwTAlwqvHd
7F68UIC5JVJ04Z9Wo/oy49siiG0KaApzvnj9uotTbcgOaQrtfZNbGzTnig9HWVGztM1ftxx3YOPT
46/R3fYQdxV245siyVx+DLDfa2yywVOR/8wJWJ2FnAR4flZYlKi3o0IN+M/BDXUlZkO8kT/z0xnp
o4EmExHEe3O3HmXVAbRtwKjzsNa75sUylA7a9DB3J5LXqcs+MZ14EHf9Cq6sgVwDcBKW0hZDd8dF
nydb0U9mqHDBUQ9S7wEzc9DgCRROQvEv80A0iHoQeVwFQnQIXF7Qkxxc7FHjBnnkb6vCn01I0iwn
d11Dy9gUznbe/zjGUXSDsW643v5WrAeCiiFwC6lOMBl64Y2a2gpzq1tnLcuaNto8tL8Pz9byMH7d
gj9knJd/sk4+p8iIcCQPYfKADZUchRinmsR0gO1ZdET2LN+cSui08Srgul56REzejO/qJmz+Li2P
UB+aJjhXzy33ya9Mg7t+/ixGWUrLRhttLEAbJ6lVI23prsWJRaMwbIC8Xzi9CcFr0psqdiaVERGO
V2lttJELR1YJv9PwtnkETmWGs39lUNj7RRuepRfbK5DSYM7w8lwe4P0BOeGHVKQcuXgwCcCuS0jb
zB3pj/DMKZOFxHa/DbilE1w2k2c0duIrXG1ziSY3Abb+gaoKxioKB4uc91TjMpdbpGIjbunlGUFt
0PbCnnAC58IXy+tBtbQZ8Ftt7k0rL4ZUmSwKWgDD74KeeFLL+a3dYO4/daU90vlLYbNTxnwySbBZ
NaPwa9MHiawZcLt7gRMYXLG999vRkOf9+czwKn3e3SZtQAC80qBJeEwMZVIg2ccIu4H3xm6rBVaS
CYBHMLkYEoT0B3qLbn1k0rWvaP10/rJLittAgyJXvEBZSFrYm4egFxXk9QFf/l+SFSgOPAOtI4sj
5MxPCfexyLhmEiyMDNwtw1iREXQn7Vngyes2KL+FGvzZcEJmOUq4+jPvUAQwID0cHHZzQscRr9AE
u96ZLvoG1ny5RdwVdDG4zeYmEfIatixgzKpunOy1N2vMhKmMeDux4PZ/Iund7T6yOK6g+lfIDaDw
vnomX0j0lQECdAtVPjpZQom36Z7rUCQidB5iZQv5lDRCbxk7qq+K5ggyI9oAlQ+UrK67OOPaZicw
D4vaCStnKOHjNvt1PmN4P0sGUDIo3k6n465JbHoVyOCgLJVkFAb1t6SSwKXxbh1tPZ9SGNdDlXV+
y+07ZWiZqKVq32ldtnK1bBnbb2Ags7u6aoBsM0U9e+SIGkMI9dvd9S0b2x0BwJFmV0c9G0/7jZW/
kyWocI8mleXnQlbrc1HbGgRb6AIS7d39Zd8dPyBu8hwd13NHJDIWk0+RVOqvEuAqGQSVJh9rpbKv
0wzAh++SxeOFn8XgeeNK9iF5bqjhAVpu9FXo9HU23alXMB6gd1K3WdxcGHOb0KBpcTxGbJHe2rtd
4/Q4spSOgBr4aaV45s7CDfgnmZDOKWmk3keGtddIOnttP46PyFeO77NMbTylCfSW7JvTj2fbe27Q
53+Tgb2jGINBM4AA5Cvhv1RtSarvb+cqa1iO2cnrQkuU1wK85UjSrBsF0IlDuEsrGAC6cWLucb99
MKnPJws0h1zM7gfAFCIVy/in5FBWJfkZ+Rh4o9mW7Hhy25162+3D429QEkjwj0xwxDXkCsM0+E7q
CMdfAj5Aw4N+BFes/2l0JoJ01Gz6XgIXYJ3J5eXZ1FDJ3+gl/sMz1brNIsGDKtUQnCnMML0XwGQn
kM5CLtWFI1ISnjFaK/AccdirCmD1sqewMAfHFiOAnfXZaVkdoykIS3cIxpWNIqHBkttb8qDSf33l
fCIAnQSxl22HrG8Ju15BFSKjBYcaSDBEFTHQgjykkMiVd6up5aqnuyI+9iHGVRoOIQ7wDCZUMSNd
fGHrfFefNK79sKMgYfGaGcBkFAv/xJZmba+YOFdFeBmkumZgVrPrqWcv/JRDnHgFnoZt2mcde4bO
zRy3sUUbBD6tjxj9WtX0nM0g/aCd4P3x3NDD3Ryt47gf1Zxc+UGK0GYgaeOdQtjiNAKCIbbrYk8K
iY/y4AlZOBG233l6O6TTVsCPobwepThC1NsgGRNKi0lJmWg0iTkHXxFlRJU0zv8+rl03x40WHmD4
3gIXBdqREluFgvL4RZRYRuYVAn0aV9BsFjc75aDdD5dff7C9vGDekWrgTSIo2Uu+MlT2Uc+IzuXh
qZp82viWf+l0xTQst+V0z6rMIhF8A+4BL0s8Dij9vWJ4jdZNB7K3Le70oEjhT0gcAvCmz3ekZ5pv
P7J8SQDwR5+96aQ9vfxgOpWrl5k9dq+c3yG0JxcQvjw1jYcvN2Q/2xqyRG5W/KSYJERiueSN/qlS
kbbLvpdvEa+GiQ+xxPVDdQxtsdEthsa6YQfxWsAiS3XLKDq/mXQIr+l46fm0vr9Xt49HfduZ+OEn
vtP9V+jHMrKOuikWaivCpNUp2t/MNrWyTAuwU2OcUjDf6Mu8301kNmTu+2jgHQDMrEnOHbHbc78r
rWhcKR7zIWGpPuV4fMsDd+C7FYUKl6tr1BV7z5QctVKirzu7mNbMQiqZAjApt8RmaIlQfuvgLOI7
zp0SZCnV/jYXpop08eEZsh4dsQJk2czufU1OB71i7o/JQBe8V0rh/WxzO6GYv+lU01pGcju3MQ6y
UJbUWJXjTy6dhLCZJgZgALjMo77DtRm1Z7FpkYxXFXlSRlMecLiVvMMZ1lqTd2c9scIoX6UcHgLW
cWqp8KMn6gmKExiJKDQPklObFaM+UDlc6CiEdOp+kDdEJUD0I5T3isCPL6/eIC+KT4rIy2nw1YSv
EgAPFcGGkWvn4C1qeThpC2fubkcSpYxQBM8VuO4qfUzNmLcc9PrYzs8D3Uk6J0EOULYWauvVmdhq
lzVim9C+WA05ljljex6vBmDeZa5aVY3kTpijZCctnh3K4F3tQMBebiU4xeomMvcZ8PT/FgI+0BO3
lp4+8Ih5BckqIiQtGm+zZpTamlJkRtHIuxFq0E9m3pcJpovilY7/ashIo2BreGe1yYK2p1pIVRre
bkupXsU6rynjqXTCdpLmcIpEiAU6Mur3Y/x1ShWWlPcg/ySeueXzrgDyA4Q1Kdn+X324JV/FuHgZ
PLsD6Mvog6WiResHWCkim4POTsm3aZSJu7F2Y8elcBnAEyziuyUL0RzemgmrbolVghKKsWm1a7F9
t8Ln1GlZGrvWAPMckxwzGB0qG3YyYH/a4LMVWslLue9CtpusOcclYJshNKTM8ZMRlWiLOMk4zcrj
P6HNRb/AUO0zBWBNRA7Czlkxi6U68XGG+W5HUywoQrBCVtG2VbTXeAkOs0f6VFJL12ivR59vyF8a
2fVHiyw9Sm+iJEljGy62r/Wms4T7ucbkzrqWmhxqcM6rQc56373j+l/TkSQsc8XtBVUvhhqatQev
EokwDd4uDis/eBgs5K8wtKY55q3wlnZ4gNLa+U+BvwLP+c3Fbcaop13CSf+G1CsCHpx0cdG4JAr3
UPwhX09/PG8LPS4HCd5BnZUWBLRvtI2HDEyG0DJ8KiyaEbPhWXBDXizQBySbBYwXNiw3ldExfVqE
QsfCYDT9KXL+4lbthsNpyplGieY+vOqEkpGsPAUVW7mnvN/Gg62yGKiloUTn1a3df9i9o4n2rem5
6/8xLZska+TVX9EtQ4R+x8c1Q7TUIKfi9mmQ9tyD9QtsmKx8CnfXNjNE85beQcS6nQ7fnkdhueLh
aiJdnb3tPwIf6Zp5bwTfzjURNoo7T6TaPSX+WIB2kDKWoXzOqtCBtkqAix0auzdcX5jVoNzuC1af
Z5O+CMs6GbFIH1sgcqVkv5C47y4TbjVQD71R+X+0cuzV6V+ZsWi2dTduzGbE5PRw3kNxvtp53656
KX9mLstbwX6oiB4uq1ylfow7GZgMQ9CCbbs2AINKW//cILT5ERlEBVsSEiI5DzjBoi75QxyiA0ni
X37kbI5fQw5CDg5VVVT090VM+OS7J5u7KDS3IE1DdTz6DX9HCNBLbwzZNNXKt/hc3L4HtlCG4PjV
pmmo4JhhnlZOmLekEb/UhVC8jt0pY6Sy+RA+WehxeE6guZdHiM6OH3+SjpvwA6ziqFfN4S6sYzUZ
NHq6gJRB3n2kwXAZvtCAOwBtLQ2IRX3AxfTntnTsuRrnhTQmDyRdEJ1jyIWrClQ7DJ2NQ9EpRDVY
RLaAojc2xXWE8Zf8XUnrW3/G0RE1YyIlEuwJ+PHhGsR8b6jAQanzjgT75aKk/g+dGFYgtVHlcPs4
ND1tLrC+Qay1cd32xrfhy4WkJcocuwalUx3PFvKzTVkWdlA8n37MG31vjJvssrbAM8yX+sWoZSeb
ZSAIwVjGk/0IaoXsvo14aavBXcUIgv+n850OF4hLsgmQI4cUKIadf1L7Ij6blwQO46lKWhU5iIrZ
MPvAl0IDy5ehKNlDaBVStrTdqXuniOJiGdM86hXI64IVae34jewZ3owZqSApbY9XpKgGQPr5PtE7
r8lhGR0G1ZnUfkOoH71lXqJNWDcw0RsMfXzirc+DwHUlRzCk+Qpc8bx4/PFtxqS8/ht2r1q94mb3
CA8w5MGfk3KgsPiaeDHpna0G2TqyS4TWSCGktbuBoVhfcIq4reD4PIdx0qRBuQ6sS1OFIDuVaoJa
r//p6cMeiNDDKRKoVMYw8cbVq1Enav+al5O/9Fz2VJEgxqjLEXpCSB8Ch7hVNA+NFUOTi9V0/JKZ
yg8XJzTrzONwvrCgfMQdLuwqyxFFZfns36JQx1thehi2+Cdb3XdgEMAYes7CqYVxzqTvqN2H2nu3
uOrUq5THptEOtrjwmjE3hrHiPwmAXlHD+f9VPOw9p+zy+FhkU6ErE4bEOoTOSNj/u0p+Nm+MLfVD
4aSnILW6qmXeQbGL02zR5xDTNQZct3JvSUpuybNaLyJg6AETuSxCSdAbseDPB7b3+8tpIWSwQOut
lIm+9u4+FXHK0DjmVZOS7CnO3ipaeoealSkU5lzVbRsxCwdC452hb8+OOspseLglWjS93qjOpa5s
bpOm2fQ1fasjPhqWCteBiywWYB3U+ASb4cQbTk2yRIb+wsGdtfP+T4cYuLhtOpPfKmhgbxx8oRa2
Z/dD6z8UWv+bXcnRvoUBYlgRLv3gNIzGQ5mTb/1tGrUe6Ias9jbmWhfGUJedH1110omazjGDoKrJ
dg4yuDirznwxbhDcOldqcTWSZYCoAZPcc5RnlPnSeFqatuL74RTEPoyVG4/yfQHoVCygiSpOF4R4
7fSNvpEa4wODu7oklPQa95Y4LZlAeGNFw9dXFJCRiNd9VXMVm/W7vmS3haG12r82S0uFtrXLl6ZG
/zq21M2CbXE7Uch+mfy4LnwxBmZn8yj+zlylVGOcHIlo+EIXKtwokcIcWmMYi9dGVhbzf2UFxyb1
fm+4wH8/b1D6a5BpEwFDkqp88vKqwbyGlokWtQquSLF4n0SvzMhSNzn6SIJ9T8xMRMYLneHN+rI1
48qISrzJkEmWmXPKiOyvupj8CWrRCE3xZ4jRebW1D1o7YkRAaIcH1ZIBYX6bt9jvvAYTlrGu7Od5
JHkQYgapDsysVEDpa6wzGNa6otAjGWyIHZD5Hajb3tjliNKjRXNB+nXs/k2VOdJzKmbf62Z91cXo
lWOqYwcwqH99FL9+mNc/YX62yLI0O2b+P2oOB55Zt3IIH4sXuLkJB9RKO52nm2NOkPi9CKIfgRqM
RpxykYhVXzdrCokWtHKOfIC5LhHybwMUBt1Sqr6J6AaJgHsk/7fFull+1i76TVjiJ+bH80iyaOKn
w5ElNe2Is+Df966RXEIHx3Xe/SCuMxAmoEvA21IbaurSpQab5+hmvePptB0gYlXuIXnAIXg1Utks
NMwLvo/0qHCZg8HIv2gZ70ba8Dggp5+bAWLY1iqsF4CfHnK42Mngjf78aiPv9qWBBCWVwRKjk0fq
FLaqLCfTin3EMaE8amXEIgx5eLGXDNKY7PxeI6YIXWBeQVZAOUX7YRfvTYZUv9/RL7sxga7wCaYT
dWkMsTjYWoRQASNv2FZ8V7Mzvz3RZ8q6jMokMTkEz4uq2ujUMVHdlDZALnxUcQPVAl0fWx6xDhQf
f2RgNalt/vQbliQzZMrrtygZ3FPuuQxoqKCg0sfhvW3Fd3tLYHl2/nz1gukKjIKqEstZA8NsA/Xd
eQX/IE0ezLQ/x0Szclq4ubhvJ3R0Vauo/iowp4ACNcmoRr0kHJKQ7LnzcylkT93cxojSKHLR4NOV
vKYAT8rHAZ/W54TJjF21MDoP94/d49vAMRJWQ27CkpYBMrwymni5IW86zHf+unm9Kb56yjMwLMAj
csxEHBV8fy39rn8Kx9a2mx8YZiRMVNxJXXry+gVn3oPZJhmWX18QTQQwwwttczOIZf8wzFVRxhN9
FFeBu7aVGO15U7i9D/nzxC8eWrpxCAVkc0WiIV+h8iaS8Ai4lFmVTPgW4GBVbYj90eAhjmxX38/T
9S/24F69oW6WRFFVElVsALxtxnSWqaV6pxeJwEo376SqJnAENi2+VMh9gJVzcCvpDkZOo9WZhd+K
1nmt7VwvMuOrcrMzGyr1aOg1eQRm3sWHkPQfOG7+PChOAb2yGQBT2SK/x5qKrxZysMlXMXs5obW5
4YodtVCiEg+AqhuKk2wHBMQtUCWJa4KswLXssREQX2WPyKRLC8M632/fCA8oHx0qhlySEfWT14ao
LKkzhafgTd7ld6mj/lUYDPzvMITQamixds4m0KJdU0UIfmhSEGv9emv4fjwVP6qBEHwTuFA2jU0g
IksKr9O9WhhFnk6BtO8wXBmI63UxeUDdaGVfLGowzeruN0NavYcjJas0TRy5PFPrQq/InLvVsz6/
0BwemgfYthhm2wuAcbpt23PkqwzB2MMskN8Au7QlvdVedtW1agsDpkLIj28VGs1zRgVfC8njM4FI
Bjea9sLhaz2eyruw1P5bacqYSoI7cR1/UyIdw+2+RYmDiu7bwLg8q10qeE3hJiZDYWziuKTehq3f
RceTQuF6g5Wb4NiyoRQ7Mb9tik3Pb36l9qHGTdEGHfaVD7KFfbM5Zr/2IwxOD8os+dr2RG+DHqkM
kE7HoG6+zskdDgek3qPlqLey8ebykrD2TPLZL+6zOIyv3qmGOCcTvGqa8GT/EpMXEPXUXC7/9NcI
b04UdFd4dHOxVpqo/Dqe5tnLa+Odm4fREh+OoL2GDbnIpWDpv0x1ed+44Ph7moNVsFk5GNSrr+pV
FzrqmnD3WhtBn7X2/hlc5L7FfpMjg/VSuCT5TXR2DhtaQGhW7UtnwWsNHnr4+FL3qfg3qtpiOIlL
6bjVPig3nNPtogRhHPWuHG+zZ9RwIgIs7Ld0x41mLyTqAEQ+F77cjYjbSZsljICCjUIly90mLM70
04OWGOrbDwOMLc9QSGGn1QtrXvUsRaobN/73CBk/y/zxhijvnNaryfzF34VlhBXj7PpFfXsrbtqe
IjfR/RhogBnZao7PsFGO6kbdPE1YFhbQvny9grwZIahN8z+ZG8B2AaED+oNwYhTiYklARcxsaniC
D/OKOgc8ATYBrZJzi3bKbGNWzOJcoHY7Tt6qJZ9Y6yg76l0t3fUjlMp6sBEXWmOwvaMp3wiGOZn3
3J6p/ZechDczrWYIcViUyNw22JjxjqxnJaLo+acpFknumpum2Y7mNRjeFT5FTF39s2xfq7Yidjab
i6Kc+SFUVDUnfSHuXKpVXIcKAXjPADFrb0VU0ozuNngfMN3/7hrgbFP9TavMNnnbnl0o+uYn8qPi
YgS4bzuNxpL23jcOrza3d83/s7HnS6NfW7SACPSwUMSRGe59/AQdV/aC1eVjCbM8ucUhl/q2+OkK
Ue1g5Msi95u58e5MfRaA7G0ZxMWcMIjHDXKe89eOluhHeJs4R7vNpub6mZ5hYhhmXoAE1e8J8C0+
CrwGrTWo8rU6NebegR+X6NF8s4TGJhCi/3I6WozlUVwWGHDRvyyJ3oPD+FZsRUa11FxUXnGPePiU
ojzsrRu77BkQi2YjpO8jrijRw0mrKouFweSYZgFXVMoUiB02F+cyQ6NtKPtLVQlRHXe3iLzp0pcD
SnDm2ZiVZkIu8u1rQRCSd2IYnFMsVTPwCESC5v+TRQIvmZJuCpkyL/O0s361GY6xxYpzOJ/5hbkz
mOiHpzlFuOZtajSWYTV2maatLLIFhIHydgJ+KVxMProobAYNWk6mr4qAZbWZQgoAuOL+F4HMllFV
jQ6scJ6be3glgvWUYFxCL/GwqxftwA88vJgNlYKHGKTqJLldKMwl7bDrJLKlaut1dT7dXojwcvvb
APTBRd+a6xvDwO3C6AyOnhVgzFupgvPKLZoh+uFRVI9xG4Cl7A1DcR8KJX5q+k/ZWF65jOQbmY4O
nOAX1llrohM7rNPRQ3Z4SjdfK3Cl5XuCk2g8C5fMG7JsnhKkRbJOiLUXWgKLnRn/Mh4rDhy9bSfy
UpqoUE4mOl6A3bQADX7soyErPqTUnke9VDmpzWapPR1ILOzIcLktmXqP0kqZ9kPiVRgBYFdNSN30
ontwkLyDRcH3/he7y+iZKszqzOXWiBeKaMmmuEbdl0gnz8YY0UTr6/2uoG0h2+RYa7Nizb5aMfRN
uRE/2iG7kRlAGyJ7hxLUbV4mx05A789bDiJLP7HrQVsxgT+e8k8BXhtT44wclFgrK4n7/FQNjBtp
s+k3z+Z03tRQkUMBjQO+aDORyRB5rwXJS41s9MkowIIrnY4QrqBQFhHK439zlQXVpleFlWdD311S
ISxXngxIJpp7MFv4qZucq2S196KJPVEjALa/2em3+xPpjamJXEWqiwGx/J0LdknCoR20xQppCkIU
0qE0ccP+k79xREj8gOw8Tch9qO006BT60R6CSzTR7v4XuGj0munkUmT3Py61VsfW6Fmme8OeWD/K
8NPItPCGccJ02AQoaeayeYozfV+NaT9l+hyFROabRBuYz/SWYI0TaLMfPeBiE7jI6tXOHQvdJs2Y
TgaWantfAFe9CyFASXK8M2z7c8PzoC+9FL2FL+U3al08rkqQitapfsUeje8/+gaBxbaBytHY8j+X
I/4EbKKN2YnQ8Ddzr8dWijCwjDlAlQuH6ApcrcAd6g5a33Rbbaex73pZc1W5SqaAb9xvgYk/vDsv
S7vOZRQOQewj7Vdaw7tdNGQCo1pcAm60RwKOcfO2jj27sspG6jGKj8pLa1mWrnEwKLvvVQPTSwtH
JCXUCSqTAKoDw5a0+8LzEhWm1aZ5Pf/7EAnwlPZO/WvO2sx/z76WfHKU8h5tukZ7WWXmiTRuwazV
Om0pLVfUMGZMA0MJVrHkgRSIpU72Au+DTF6ZHvC2mKtju4ezGOKpieKBvtIDbvPj6fwkcpBJaWWR
W30/ygDTTPkEEfm+n0jT7usj4BP3hC9M+2XmmzIbNjZ12Aa/EwMWHNGFaPX/ieBMPXyPaxw2WYLG
uwKuXzQn07IQNSAPWL5e8BJ2JeMvQfwEcx7HZf44f8ku7Z128ij3ohCuQJioXfmeGu4soh3+NwP2
p2HMFRaqcyGIti9WUNrJr853KylM4HDLUe8q+8ysG6lEKDHOi9HEFyjf7rXxoGEiI1Myee+kQAOU
tNYhxZ9JOQiGhHnlFB+FznDVlwcDefPKAypfkeqiUQLzqiMW1wk4hvwna2wQSzA+AUywhkHMvF6p
M5m13vNUDeP3ZScU3DznDUYBYvFNfioip4j9EuHSq6He4ye+3BaT7NumrMHpvtQA54jc4rWZ2Nfw
sp70cRwuBHc7qCeNgnX7n+dgDbGyif0qHPAhRhnvsp6PszvGzrsQy8/54scTb4/yQg61ZPS2m2V8
1zMay0VzqiALJARO2jYlfUwv7nk7zpk6HK8n90SmxyPFGQ7Pu7XucPbjRB7SMU6C6OdeCNjBzBaU
7swXiaTJ6jkfXAVk4bjSthE19NA59nrTSXvXXHgy5UUvNfrDKQ/djy+iprhIctXVURXxkxkFGcxt
VEy7MVyA9cU9UzwcHbO3Xdt4Cfod0ieVih2nN2p30Fmy6PNVozJvih5yqga+Ymf3cacYWB8gOkwf
adh3CVl2K1DXwYipA/bzVO4cn8hk8vGeZqQHH9j8JYUdVr+0pyahoCBvnUEr9U42NJccsIiB+Bs5
CGzwLySrBNM2zOAQnlt8ylagDOL8xhY5n1kLVo4iem5YZy1v0VMzlwDvISmiOPtaAumyKprZUQqO
YGki1nPaZIiqfQO1HG1bK1SYxpuKIVrzs5bjnM1U+kBLFmpkluD8Ry+vXJuOm7rbc5qIuFgZT4Wb
UYjSf8p09fWwutDkH8U5j8IRFn008MqpIaCsGFkJSUPia+0gL+beWDYrd92RvGcH6ht+u+H+NZCi
jFsM3LOto1lqUDfwxSnarxtmNuhwzZxX+oy7J4MQiJnJLZZxLr77AHixe9FMi0NkWIWRNEcdD0gM
ZiE+vOOzvfDKfLweYa8gb2D3M9iE8aOvJ3ut3pl7aXVabE5TGF82t44zwZl6u8+jYZ44V5OtJk4a
furs1MA1HdiTHwoUB4zn9VHZGNEtzS0YffT3tDxBGWVsJpkM2DGQJ7dXgtjMSa2LHy98+m47oaMN
ivdlgdhnEGPEr9mS2GfmkHt1rpv+RA1gfYbLIeKCa4j+iCe84UP2FTu4vr09e4/amGueNR/9U8RI
yClwCjHmi//cXlRIQ2Q/1EHsI4NzTfXvuFBEu+sL0es4LAN4JN1RheG67Nl6Z49SUgaTwoYRunJT
ZAP5oAKofrZSu2zkT/c8Hud7h7K8dIdf1zm6F/fD1e+SblgPO/xGdCv0CzfWSSmPDB1ybqPKBCW7
yAtulXuy4OM3hLQyG3dzD1V8Zg7CPhztyeL7MmM2xi0lnfaspKD35jqpsRZQqk1drI6QFGwwkhfL
hCDLboTK8LX22YWLXw067AhuJ865lhAksGmEdTRlhzxFpvx85nbw1N4udZlpIFIjYO/IN+PglFNa
sdelx/t4hupGbP6fE7jtSs3G/CRhzIhXUQe/n1rxpUc2UqHdhv2YBWr9wy4botW4pmN+HiqSRw9d
/ktPUL9l1nqh4DPX8jgsWe4rpOJRgNhSO17mPMS7mYYLOAOcYniPfujGc09bCmm0atAMWbXtEfIB
ALaCXb+4Py7g2myoQgTmObWk7JaxDJQX3aW2C6gXJ00G1pZl57ErRJr2qzVC0mwp7W5JqTOcSF8l
4xGpqKiwdhbQlRJ5JTUMXgtIIftWlteIstWsSvD3w2YJFZKGATYbe+3+mM//icm8n/yw5vHzdCm2
uayMEYbShFGw9u+mJ8IvvGckI4add3M+VXK0Cs90MraFvxerym3Ensl37vTH5mOwbY7Lz/e4lRt6
2QKJAJ/fOa/UqDGIkBrl2hyMSUVRUGq/6blCenbgHtDwqZvgxKqrO1v02LMFveAsiH7Xzqv3Rj9q
xpYHvzRbOgG2zld4laoiLqRGZsXm3o4aGmNaOKaH7AIJi18lPQL6t0WtdxRbjLz1vwaMOKR78ehR
6nsy+dwlF8eDysOcVtAZ87YHdXati2oUliyWY/QEA96pb6k5TOCLhxRVz4eKzm9BD4bUmWhoUhNq
bSpnJW1NQR3QU4fxIx+AOXGMslz1UQsYp7tHDubvNlPlof8TNfjJjZvmXYAJfVr+4O569HAbq7Mw
98fsX0xMoktmk+gI8VHOymfGIg+h0apL0fxvWakfwbIXJbmN8btWcys8drTKeVvvnNRqXfB0zntJ
jp+1WQIvZLfS0/978E4gqIBFNldc1Fqlot5wOEmf0seyLCk+1gRj0P1KOy0ac4aAAq3IBS6x7Bwc
/3+N/zeqLae6ZdsXV6TL/XlRf7t/0Bo+GmhnUN6q1oqaKBrSHwG4bWBFV8lDPLWDhK8VWnPl7lvx
uM3iMHiHsDG2y6vgLL8AXm3TEeSvqqnjKimgQDSKJLXuhUem8wPjRcX31CzF7+9kErP22wQycDZh
Pk59KsPUGF5LJualeYnJ3kgcHdl8PthsuZ0rZNRuF4+N5O1NOhNM+ShKiwFPyZEgF/I+QpaC5TEp
E5dJOJVS6PG80ler0t2FDxTtk6toCftRQHVdmPGqGCo2uCqaJ4aKuG8OZR1+yx6/zgMDn0IAHzZU
16m7WM9A9mBxvPqR58jukmydQwxLXBSod/SkZY9K0p99bPpvdCG36oITm3SCSrTTF0CA/WEpH7FY
nFEEKL+i7kzoJszHrDyj2/5ZF1AXzRR/LkyX3X+nCwJvzHD3IomcJ03fndri37rA0NLpt46E8FbO
ERAt/2vK9THTqxlAyXAFSVqIAF+xRYfwUkwNWjrQGs3higCQm0KFYFFYFo7ag4rIhCeFoxouDq4M
GDjzIa9Ee2siLgIjKKq7Ad1YhHSKboMj6U0zidPjq9FFD2AzfZ8dCl5GeXx4qWci43bXHsc4R7qo
tVo7D7AYoXuo41NLTQpgtYfHNyrcwdXHX0dUjm7OUn0GL0otEVEGPh4wmJNfWDTvi9XvoejF7ajC
SjuzBwRpJghxGQDrV6NMINZma+8greyagXZ41TDwI9n1Er0+AWWPUBuZXnHkHnhXg9fntYJaJLUP
MR6OmMflGNnSkRTYlxvjJuJ8Dx4zGPbUNffgl8c6Zs5r1ZJe2goH5ds5DYdnk1HqUYWXrickG4I7
UaRUaOhiFpyIbmYMNCrh5L0TXyp75p10j3GTbqqknXWmHw/vXDHoAdqOVDM6XPl+QucA1/0J57Pb
D8t05t4AMGBVFi90oiAsr6m11oadrBtR2jsECTJMf7MJowehaqPs6ooYcH8nLbvur9H0R+4hpv7+
WBhYvuxZo/T8TcvRbNhWID3o71whqe//h3OhASMufKxaWpza3mg+dX6LjDcLvOYuscabdXv4gQNh
xx1KusyjtUgii5s/nQHmyKWBQjOjdwt6WrgFN1Gvw9yaPtZwXr59Fdwy3IzH0m8h2dg9lDuVnN4w
70iFMyDoT2a7+1WiQrqEoQ+hWPtpEdv/Hcp8YypkmJhd9xkKbWeN9V4yKpq1kX9J0KEJIUXt1b42
UCy7PyVDKjOX2w6aS4KoG7i0JiesD2E9fJ5A9zdwVKqHgi+4z+9pCQdVq5PgKyFuHcfI0yEkdCfs
Pw1tw9PAiSz/9fuiy3sFHvIKZLt+OroTiiLyEKGmjwDN8Z+WRPITa6SyyhAmb5h2puxBuIvQx2Qf
4T/iscA8soGTNZU5zg/irsxMoLFtl6Ak1vTveNMzxorIKi6+6GAsvdONIopZISK4mwe5C9sIbgcm
30dMrcCjh4+lUVhJVnjCZ5c1AQbmFqcU3k7gj2IK1Uj2iiOKWIdCa06WebTU/qvuorVLRiVh4kox
rFiBWT8pzCLpCWe7tlToxcWYxkFb3Ckil/fZ9Z2yWvR/+/PP0rCKN6/eIK8GlF75kfTzzalUMSJi
ZcEIpivSp+WPBF/+8W6DAV86FK0F7226jRBpGU/BQ5XBBkQeNUWZ0bEVA16+M4vbiGn7ZscdjMBW
EDrulXo0Ll0YCFs8vP+9V8ukkp8VpP7Dxlj935vBBFukHUlFVcKD5K5IOcW1FJ2jZjguk3acl06S
1tkcs4O1PorwGUnj1rueTJyB5APXn/MjnbhrlBbuQd3hAbI/Sm2y7cojvmq84UHkzkEFgsFnVzSc
3VMdBfiDU2laIiPwqJ2OuWOv2+ZjakHXNfk7YIvM82Gy7P4/g3uDcts+aRDavcRPLHDN6QNqppyG
IqKciCfOiF+yX/nuprTRtDAJZguPQe9Hf1pNYenNqJzu/YmTYdT6fbrMFmnXm+yfQItjZqUNjcpa
5OqppJq8zN+3AqxRSM5lgl1qVJsWpAZbWn1U1ajeXzIAR9SUexUDY/T7Ax30RZKESViBCwd1f/ER
IMph1uqMUAcxe6647CclQWzG7MQftrYmvJg8/LQPDaSH1B85N95I+JrkDzVn3/HkQ+gXuycsWo5w
UTdY9Cw7qNMqd3XLbvKp00UASeS7gRzy353SuXrtyAYFbaD3F36qhbTJMH8wRgIxODGYJoIjfRQC
nAEZZCMbCKj7Tu0gjLC7Y4R5FIc+GwRQR4HnyDXJQP2oWcZyuj4snxCkfT63foc+r/ZbDmXSb3IT
YGpyuOHqlPzaN+UpIZ8rtVFrUEFscv+T3F8h3xlQYUy2gqipJihUDAH7+akz2vItNrerJwSeLcDq
BhuXsLLr9OVPSH/KLuG3lIwc+rr039fGdNdUWzE7MP8dwD6f1iIN2sHe+yk9RYbbGUu1wr6Q0Ngm
0A6hbAMuDTwUhqEKweZJIR7Ta/Y9skIdfEURpsm2XEQ3g7KKrVr8Gf0u8/cvtsdWFRfV7rozzIaG
NUC4DShjkZ+elBT+cLbltp8ZQrb0ZkHIo9tkvVs8x4fFC/xiUBkwFkBd60ZhLoZE7zH/hahfbSU8
9Vz6ENZ+hLh+F/kCdaxZ9EFGTK/Hsj+pDQFKHXtgzjH962zoOUXoJDiJrguXZzR/lWJRpZEUzpx1
rBnc6moXtu2J3hfPVHlD9OGKt0lwMOjgqUIPgl5Z8TuRRphTUhlsc7UP5UAXJQEYDG4lXQ0hoG2v
WMHLybOuWMNgTXaLQbkTDWxm70YLmkZyTJ3uFS4tMd0Z3b8onZ1sFH72BAZReB7RML/tbzwgPqbJ
+DdZhJlfXA7u6k4YuHLF//Q3ln0jTP/n5Q9wavo9ZWo/+aco9++twNdQtfnsXDcTVjIDiabyEMAB
dDhl0N/Bk6zdnsDHW4hRbJzrgJOTL2Oa/dWH4emYaBMIQXXg3fngvz/rYdtcC+EgaD+iljEZcIeV
aba5TQTIKDswM5DsvKJJAk9Zw3qjo6XZuzhJd8cQ/yqbfMeWAYUbUKN/kg0lTGEw+2SiYt4gZNUh
m6N0p2RXdbjkJNt5LRHX6OWUJ8KDCfZaYjnvxx6X1ew0gHRrZ5S/scBJSlU91fJ4mwXoGGX+/0NP
WH9Vw9B1q927bcRiKS1o8vVb5qbiGQjnyd4/o0XGHd0v/SYRabOnlT5QAQ5FmTifDFru3hb6Xq3T
YZE7KjDuPkAIy6sHJ/93URyDnwKoQoTn98muw3UNmDUGgxm8ppZDGPWNVygg1lHvQbDgkrk8JO/v
3NyPSwwSIZi/Q7YqVck8nqJ5YXV+A4wniEkqCQg31nojUw+GfbfdjQ/+KdXTFgGokee0qmsoeJGP
T/ELdwLNXzkC+qCNNn21gMOt3w2GnyUcKrv4HvWprKy6wB6wpnCsQ3tDJ7Knfc0BsvSOpyr2WDti
LK7OoxwH9PaL1y8EE9JDrm0kxt6q/QvGJMgvlmv411u3exsgFzwpPC2CrLKywHBe5DfTH+MAueY+
dAZtKrGyQb4SJgEOcAsvtH9LqUd614SysSV7Y6t/KcR3FUaSzGQ4+pU4DymKSllYnmws03LNo9O3
Bf30adzKsceJk2HL+xvIHdI5a5o2t1I0tvYGcwrK6zAyh/4ee0biFiZZKQSX61aYpPm6MnZN0cZf
raexSkVZfwAvBzbCn/rmkX2SUY5wYYkieicrQqCVZ5CInII5Tg5swX+8RtKcioqBI80NgqmSHtle
9rnb6eebLafP8Lvs9eZJPW5uRNda3qrLmMmtBewY3PtM/DVmwdACzKqnm7eFp/PN/XhPr5eAVPPa
uECI7NBaIZradJLkN5LsZji6ktFSRMlM5L8P8EqejhqRRiNMNWnItJMQ3OaPoZU2otK59LEvp9o0
QlaauXo5TXtTl2P6IvSc6u0zKCnpnG+X23vi5mMmA3cIBaqJLxII8V9yy78dL10uhy0JqttpwnYE
a5m2CUjFRiG04reioRXa4b52oM6uyPNaQIafIQhCnmb1B11tmqGQCvilK7vLdhgX97CoLjBtsoEg
1EdaIItlP4ZI3XvUzLdA6cyL8qrwA/LwukLMHh27aeUqaJSSa+2x32yxfAwFxXui8phx3JqsErbr
3JxrR9X59ksXAKC8xsSCF9vabV7eSsAICE4UTy4RvD3VXXFW/kpMMv/dn4AR8jgxHb29w6a9lqmI
RrEF8cyw3Uh5m4seJMEziD9AA933GZ1zJq8UrID/Ii0kvCnVTUwxUJ3Xv1sNKW/hnCfpgOoDciB+
hWRbfzegPaR8p1Btk/em0RYM7oKOe7I5l0XoAtexptRIOqcebG9WLteDkammjl0lSzUlY5An4I5U
vudZFEP6hT05V1fuhZmXCM7g2cPipvuMc18dIuHUTWYh0OeNcxRhQXV/z7O2PrsC4bSpct5LTDnC
sOS0vWaIdlMUb3g3fW5Jy4PcGp5QuIETA07U/P3wSnqTh+yK2PG8fDwcZMr1BtDiqfwyDH1zqy0Y
XMjDdRqdunnIwbU2qPfIgLckFYWzYCMZwlMSGD+ypkzW9DPv8Gj5fG+OJ7/VGz7iAN1WWepUBUuG
YYGjXfeiCkwVd3c63se/fQ8wNEwoTf4Uyt4woeD3VXoygZKfG3X98L0pbjwJZgmRNClF9XmLop0M
fgVLd5lD0665S2o0jlIdi1B32QlE/ePhUHRwjQo5cBMBZxTgT5qOS3DBTRVATtsv47ooI0Q+BvNg
cpPTrTAk2olFT+5ajQxEwQoBDkN487F3waAUWFYibRe54cag8K3+jcKjHMZdNnYxXK+uAKSRYD1e
eo2HB59bIig1CHMvqy/18XgZw3aFm5EABcFp2kawYRvCSxxQWoQGzqcOV2Mh+W7AIwg5/iqUQrFI
RIeLmZVa3po9MIIDa3ooSG9jWROxJhaM4CsgHHx9Sxkc1s1LBi4AUuEoHlWwp+14KmBR8pORRoH1
+orEzAiFxgs4mo2Hkd4HE99TXZu6pvace0MVNx0mxPEtuAjJg99z6yAcdyKCoKy7scDezJDeEsXA
MEcKIFXtEcJbWbcv38fck2shLw0djinkiVjB+VN5xexwdXLnHay/XhMR+449XU5/VaarXP/OWHNF
Vp1xEl2jGayx9GYHR2IHh9AA/W/w6umzhpQj4WjZHlYYa9XMb/c0d0iC7ILS6JpfzYXtQOhrON3k
M7jfT/AqpDySjqw2ZOb2iiaJ7psi3rx45yuTtEO2KZHcoGtzNWbH0vz1zH3DZkYJ3+dYXp51f6QU
ckObt0tKkF726+1LdGyQgsjxvPEKos84APGcrl3WgZs8anCFfuajgba/VgzQkuxyXO8/+i4gwYDV
9fcStgsUzFpXSx1wHpMtf99EzoOb23eNSiKicEDbr323JTmk48DuP7sKSqlCy534t5HEqKLU//Xj
iqDgXQr8d4BRVEbyMHu34i+wY2wKBC11073JT3zUG8DE+RSZPyLdT2K1b3vSLDMLP1IAGGx0tPHa
+Qq5nHti/i4EysTnjiMJ8GyNzgepb4VmpFdn7DMPtUA4AHkWzuDxWn0NkDc7B4JU0HH3wou2LNaV
JIhSAc2pUP+NmjoUkkva8LuSjz7ZPdMwHcH17uBgwA+EE638G3yTZOCqjUZ5S/rmAw2DjSLE0tbx
C8Ce+qGyPoypXORPJl2sU0QhPV+GuDkqVaXNXtlfcPhvt7e2khcN8dc5B/Mxt9a8XAwbgWVLLGl2
m6IdMBUrwJHPRQKzW68tb9bwqKe6r0o3qA5Pr3IUt7Q8ZpFrzF8MGcSglqrLcCy5lDvHiuh+D/Cz
2k3PKxJuz0FRDf6vtZ1ndc75SvIwE8+Hp0gFjKD04fTeUJMxiJoYJnQ8ZcF42A8Th+NK+yCzO3TM
OSORSH9nODC7C/rLwsDEx63eGa4xBYyagRepdAD0Pg6jkYTgwqUJ5FS9rTSdqgXBBKAzCjfymwSV
4bbxYYkvQlc8F7SK0aXOxNnqS6NakuqlWSgbxTaTHKmzZlcdt1/bvKJ0rS0MM74kn22zZ0cohJY2
GzKcHIXPdaoecWpfrhF6Ckkfp7B0SNFNrCM4Av1Mzs/cJeQpHc7xcQpuOxLC9uwGuNGC2A7408LF
8/dwRVjOmiYvlHo26YEVCcxj8UroEHGlQUD0L5tJzX5EdCvHA4tq40sRLu3Hxl/JLinZV93cJZoV
cZ0d+2RHJyf0+DBedz0go+myeyj6L4WsVr6O1Lsd4ByKUl086OgzAaFepGY9rkWUaHU87qYJG7nM
4276GBmnsmZAmd6oY12nE5bfVW862aYmrmIoE9c/mxruRNAOz1lw/vu/IT3gjrP2PQVdc01BO2w7
1zQA2xoxgPyuVVNJ7kQNI837oxDBst5FoAyoolmey6LZ699Sm6CTSWugsRWQ7rdztqBWEnp+W8fi
BjJkNi2d5+SHAhEXcrJEan7aFCLb+J0ibLuXrCQb+SKmmr4kO3ZcZABslBLgm+ObFBXW9c7kHE8a
veFEwEgj1ml3v8d1Mb7duRW3EVeNS4TDjgZ0s+doHfFm4I1F2CSkfRgScMAaqSSCVDKNp1pCXgBz
YNtSfTv9UfuaAke2t0VU9DRee/0iXrq3Rm5+OOcR5/kzsKLmTYt9oeI14ansFhNvw98GSsGHfSqJ
kAvWKW/ufpsUHTvglV1k8dAfg95IZHiJ3h4GmPKNkaSYEtcyVpk6IasYCcc4iF520Vk/qPiGMYPs
Wg57YKg0X7SLPLotpNEcDTCgkbm7mpCdc5anhtnoXkhPixU3AqR7ufDbU0nxurYT/rSxA/6hjX0k
YFjbUKxJf23gJqt09w29LeqMvaCuHjTe8KcC9dbK8WqWd9RTztakdYsTjhJQLWsd04X9c10coJS0
4ZBvS1HA0kJktvN0XkV8ur47/0VZPAekqrrzLNFLW5M+anEPmH0JsnuQbBQ+gbr5dt6hIbpsQ9Ul
Fegtv5T78y2wO77eRSyx/s0ceFGAKdM6bvzUtp9h/erFYomlQhusV0gOwIh5oJECAztIHjP2WFCq
1ykZMwuGIigPqMq2KE3yOkBsiIPugkgJqH/4DgX1RGSZKDo/6BplJlNIL2XflIDBlr0OZaLJ0dxi
L4NPzWmjguT+Zw/DwyIgAI9P0Q16MygoubY+bQbPcvi0uGPdRO59a0rgp3rOc8X6InXaZwI3ZxXq
jTypdVcTaIrrXgfz13R20+xW1+q47Q9lLpEbc98IapMBTNSoT34Mk6WopBsh7rUPXX5qarPWSyox
zGPVEmmUIKbQFUJBBGf9jZ1Gb3uN3fXSTnWBQdjhZuAjkAnvXBoYvY8ni/k/nD5JmDJBWcpFnrhR
COgvn0A/M6YW0T86nenZENZUJ3uUD4HVZWZe3DGUSOGzftZ1ou4X6zOkNRoRvfSLW8ovBaDsMpLy
whMQcxSlL/g8sEZ6nUFD+9eqstc4UnozMVhJIr1ws1ldnzrZkxXyqhzhLiYKy4NFn9v8cugLnrRk
67MWQWTmxlx4ibtTm5hyOCgWaIStU0S/aTr7eYilyj46/i8jg6mn7kMlQC97k7Rq7RlcJSEqvz8s
+6b1FiEg50Z/yXRAFoE1P4mARvREl/lvFV3V9xEYoXJeHaUReurOdcmsuFE7EqjWYRqS79JNkbUy
MyFh2SwsSsW9GQlH4EevH0RJpAORpkokcqjuaUb9fNUjJKzBgTuauCZ93FFIAkEDYenBKj+0g4hO
NETalHXlE5GLhBqQxbhBhh2kPzmpLp8BWAjPUn/mdUWCIL+L+VYXADhkfCiNFnln15DHI2S4OtmU
P47l4MYLEvRJaNLm6iULZOxJu6okxkpsgiCS1Dlga+oaCfTN+JngSKqd3Wt99GGhYMmqT0hdp+x5
OImV/LNxB476Tw0mi6ChegLSRpRJpCO45WMesomycHCy29XRVzkcpnnHBAfx3WlW1iMfYUutfDi/
yvUSTjBIlA6bxFGfHualekxzg9+aAdHO7ZebleWaAg6KUIpuzWUQUFgsS3QtjhjmmjZSZFN1ZJ8u
09HKmLNn4bj/M3OUqvG/GDgN/cbLQGvMROh9HYO3F+9GXZLuWhfVoPzP95+inHPKrpYb4q/Rk0Sz
CRtzA90Gpg5mQcC0ncgJvvKfE8Zz1iwjF07d13mizXZ+nouA341Zgt931d9+gdC6YqPcVB68DqR2
E9iThoP/Ykuph5M+1Q6pi8Qwys3Wo05ZcqsLj4AWHi528x76OVIy0z3IUHakWqLygNlRH7YyvmFI
JtWyD8SbVKT89L0+vEN1+WZAzCuDxjTBWRahdEPqzTKCo76QNImcRRNl8o0xzAomH7sYpu3HHIVl
WrjEZZwSCAaPzMHAT7iXZFFz2E8l+8n83lf1AaWvxx9PXJOQ9P7lcx38w9eUCCDwGM4r9sk1gqRD
Q0AimLGT5ENsRceTA2gyP79fXNEMLwBD0I2D1kS8DKofbTCuiNhGasGvtrSzGdWxenveDnU7lRxA
NNYLUScA0PaJaa3bU5AQTv3ZxrfZqy8M1GJRDlWGBp3RnQ0AbdskEdOdciYSkpdmbbaJUH8Wig0S
DHVCqdXf3vsdiB6jpwYmJfFIZ+agDakBqE4UjS2Rs7giqSJYKasAqwZAzP+TRKZhoIC9NihenTkn
6MRp0B5mq98T7IkWRqSsxqFsb0s/oUcNSw5wcO4zJJC5Z1viwdHLJVSNg/3HPF3vNIoEy2EZnbI3
/zLZXCjuXZc8Urgsvf+mKNrbBUu817ScYeTvm+zDghQ3L7Eg/OlPPRn+Pgwpo3jeKD294rOexKO2
ByseC2pvUBmj29+RlumtXDiNH8SYajjFnVCfnyyPZQPk5yRzJoIUtjqG6cT7hhTKhMNyw6dnPRKr
QoS2OmTo0Pfn7V3peCmnKMLVjyVTZNR8kG/Lf5zaWDUMM/+3sYI3ZPAs4gM2W58CB5nYc9XusBiw
XqS7CpH7xhUffjlR5iahg9NINyI2JnTQfcfhddtMXVXQWfac5X3Ue6EsctFgKFiJFYOddiae06n1
wKh9UpZXhuIgUIizrfMDbb8H6MOHJRe3+bbjrpulKM8QqVPp5cU3X05XNtC5wu0UN7jQV/K1B6IN
7lB/KkL4q9+9tmSihtJ10Ll+M7stJBNXBMZ5YPmZQ6HKUE35Qus5PoJZD9KfFHJwqePvU8mHKAyY
s9Ty/S4vRsO55K1uBrp2R45stLDvQQhIpI5Sc+tPNhPTxXgAlATQQFNw/5Mc1oEQnpye8h6tHKdx
b9X6Yvio4EiL/iuahS0W5Oe4T/5A+AhRVC/YKmTWVLnzv1U7/t1qC1oLZYIh6lSfusabg+XVsp3C
7TCH9Pxi7E1YrnAWzsJGTXj3hkqbIzZUZ9iDdaIKzd4YtjgZqpSmqa1xR9zXKvRPq3IS/+bEQelQ
WTsht8eBGsajNYJYa1SZ2AyeIqluzhrE08sTri2uNjLbH+44+ver5CKUIxaWSYGG/BdSUun+kqsr
pat+2OlRxoz2hH+Ud5DCDGPavYxm2n5UFZXgFwxqmH3JvJ4VW73t+tem27s//Ax0yMfnK2H0MoxE
uSVN48I2VabSWgsZg0/2yjMRoJqWOZ5vUlmsYUWWytO4lGDTvB6mOp0mTMVmo4O3MSkZl8Nmdq8z
qqzc11VCIMPeo8Roh5iaHBTZB10eKO+HzR4oHQxeJz7lq3jwWKPLDLXWMfCNj5XX+O5eZIwSsLtm
m/4qccsdnylQj9MInkTj7nVOB6jnaKzicK3KLsn81QqbsBRbFUmAmcgsT3HjhzetzUaDdo36uffD
QOHvP/ZIaa2VZ/hU79Ijj0O0+oFbw1maSWtApbJYMd9MjuO4bv+1YdXWUi5IBWLMk2pO4jNBdo9j
wR0UAR8I3KWqOTvuWc6bXm8kqxd6Xk/ozSHyHVQY7wIOJYt7S+FJFwQvfLLuttK3FRFFxjptK+2d
gYs1mr3dPZkOWabkOU38GPn+MU45EwEbryDcQu3v3w5WYr0TGEglG+ZmaDthol2lGSYwJDC3n12D
lYvEragOrCj5Za0/pqmc0FqQGt76pfkrp7efkIg/BDinJd1dWlJGCggdRUCY54oCcKEpfh8KF6qf
eKVoe6rfHXydHTTpknqjNpEG+7HidpgMKHzQvqCUlVeSc2vDkPsqBjr37lHrgYvCypk2YzD1GFKj
Nvyny0Evtu3W/gVyxJvZDwIRQjhJezZtaOVJrKeleHlpG1eOaYdYgCkcaS+cY2+w2a83buhrML3u
YdsaKWSkOkSTCi5rGqN5Cr8UvcaUhcdMBKUxpUrri4bmwlSXTy7EdkMY+wnAjev+neL7cwJPw0sL
Kh0NY0zoEk9OeSakSaBKgtj4izGwJjmjOPv+eYdYjv8khTSGfO/5pLVhhfTPDEH9u7yUY4dxmzgu
Za4BikFO7EsyBKbkoDi44E3rzrvB7J0Jxn14soGWSQwVATpcOqRhPX8K7oHb9/L+ZHMQ1HECyoQi
vqj/NbmqhLHNdhiSsFaT+7M79jRTYKtO20lpQv3doIYoasdbTpkqXX3PvWYYN6Y704YHp894Aist
smQIhYaS9yr509n3l9xU9nyAecb+rqYDFPk5RQd3h2GeWSsOAQzcwvtEuEIDM5z93A8+XzZ9FVA4
LY7nK3TQNRcHRCdEC4x18nNms+vo85VA1wMTL3nuTHx53AWC5Tb4LoZZpIGW4hbLyKRPdN8LeBkp
Tq2oQ0Hj2pdtFIlCGmqzPNn9oe+mZ+RUykRguOdiMo7ZiO9SskmVjg6ov/KTAYULjxDEAQm1afAH
GQfQl4ykUSKsUICN0LS0MKa7D5sVwfuWNEGg9DBdaLHKLVUoS8nyDM55Ouh+1tL9pxkJWNwQvDXc
Mk35m2qyZ1yioQ21J/l4wi00ZRCrMdBTaIRnX69L4JUJRbC/f6QO/JgsauM9Y/z2KCef24/bUF56
B6IikxOQe+tumYDqWj8W8B7WsQD2hDNrigw2LeQ7uj8Ki5IFf5VGABtX19ELMwZcT8DJ1C7sr7EW
A8U7z3nd00BpZf5WE1NgTbzveimFtIl9rvD/YKzzF5aXb93ELbNmxB00fqT/tGRo62PPPiNVmyas
Lr7s2wzKuaZ0IWnSY8Kbik7tHzibtwR+XDtzPazI/vW2fA+I/klrQ5isNxiS8/ZOxeRBqBLKX0GH
3lU1BDmAVYB0ktmCbkBZ5Sf5+zHC8zwrWygrsUmm0OFhRs2EcNYCdADhYK2oK9dURp3tJcCya2lD
qo5r5y6xIDzSrH/xiTr3Y2WnxSXny2OTQarxcLG/VZ8Muo11ecsf7sXqK1/BcAu4YCzWrk64amYT
f2wepUT/4GGI9T8qvB1qsiRjO7HEHl1sbMJ+uCx9XxWYpbdSQ/E4F7oUqVslpuZy/D+G4LM/eT32
twAHiLp6aOme8C7kCdWA5l3GmI1xWBrou11gAiGAePxFMarFjDQvgn9S22pFh/CtLPDa/iGqilXc
hHDk26AE7BLU+7xMWc+0ZNi5U8pl/8KC5AYicBXfPGz9+KdFEzbdsmyydWyMoYsrwsVaSih21hrI
0kjnOBcMxG3dRUECw8WgZF8m6tKZhkQ7zPOYmnCs49NofBTEktO8W/pRXw4IHeUOy4uuuuEzJ/sy
iACLRkKShEmI5kgh6LsnME1mY58el3bIG3vCZz1aYFn7mhd23t68aQ8U19LDq6R954zAFLxmfbgt
qN6Sy6581u99d2uAz68RZVpIC7DcfPHJGlc9WkhQms+7W2hvjA1OdPIdQR33tNZd8kViXy6jyEVv
WNj/HQDrSQlvToJ2OKrj0yb/zsrpRdCLRZ30AjscbK1HEPl+umOQ5mDSaubxfa1j+/EWX4ZruegE
5zBv7/DyRGlgqZWPcCGOMnE8iKxQN99nt3LJOBtMNF88leqquVxJA6Qys+AFG00oxQ5Yn4oVggJh
G6YWX7cms/akP7pXyJZh2FyHsOizpnIESWAZuyXJ2twAFg25PPhxBchT1pYicxCMBcCE96/aq4wO
jvrlhHiV+LzkwO0MuqBz37IXxp6358TvZ8qcsGeTUAV6a+e8r3fogFfHbxT9OOWvTJHabKAzRAf9
xncQ7jXocoj0NpXyNG7u+Rxiz/yp4CKClc6k0EymOsCbbk1IWfN3nuYnLoiz/3Vo5Bp5V9yiNp9Q
sGxJ9wLoS2zg2DQY6PlXEVREFOPgYP+zu1Gg9GX7hLbiHbmWR4wEfY4O3VASNhycV3eJCmYnHqas
M2qVbczhmOykqmIQDpNL5h/SI7Fo4PKCTEqg4i8ryOleF8usfB4Y/rr6AyteEujYh8lq+KiI27tT
m6J40dTm9Tq1NlP7gzCrRE+/3wfJwNkIrFkwVPSC+WZsL/OmWutldOLvsc3BSuKH4zCtqna7ueCc
WfQqIpzVWIoTvfFgbQExtMihXIOumuvuGRRqOe8QdMxihy827czZEKuknz3IOmportVfno/YHLTr
9ZCTfQS80WAXic5Ye6ZcA0jZqwdM3Mh+cAtkvs2Mvvbvt5USnDf14Pso0X3JdAIH33Xav2MAszvU
pViW9M//sWgauLU6tctkCM41Gb1ZaL0Bczi8npuU3znhdwknaWZlkDyPFV+6mCfNz9UTcvY73Ik3
RNrHByPiu/HpM1upPViNP661Eu6ucsXbuChzH0GezEUJCDHj7FZPoTWqgBfTNHgnVij87qdF1Siz
yOjs0qMahxBW9Bo2PEICL+F+6ZquDkoRkm/3DOW0VLdHUJjOlsd9G0AjiguU+2U9SLPT/xoSJA3L
VyRZlZzbi3qsjoqLq6kH/GykWXJ6EC1utuCVgJEcDnQbGMd9TlqjnM7zLPIq8A86tKelJKtwew93
8aNCdhsoOz1pmQNfJ2QLws5DKW/dm7u5NOT4eL1I59GkW0g1ddb4OB8pk7gOupWyF0APOGxZmPMh
G421o9adC2/h8iJKXam5u/+Gdo1X5xHLbf7rpb2UxSqrEBKZS26QE00wYKbO2ve0C9l+C+sPJVmG
ZNzQgkZVF4rdHBtSgz0LKoO3DeSkJuNdIcDP30+hETNMXbcuGRS311aCEoAodHEHuVDUlK5L1zUG
IwnklCGfO18IHQowbvekTDDY/Z3E8PtB4BNcx0D4+PuSY/8+2b6LrDLb8v5wfIxZXNU0Gv0xh2Lh
YMnw5AtMy8TGn8X3rU6jJcY0segeuO561+6sroakJOw+E89hBNCzaiMA32IRrNg7jyLrO2cME3Xf
tgWbXTi0LyU2lKVu8aYsIBZojj4Jjz85NU+Y2DQTRijwQypxnCcfPXEaCuGfndJot4q8jznMCJ2p
HcQzNTuQseampN0GM8T4WuKfMmr+YCHEfDjWiq2j3QJsYQxuLDU8y3nkwggUP9M4hzV1yc1B6Q5x
eAq50UGNvHEI/4EfPLRVRvig0zx3g1ATQtWDK+7EtQZTk5dACx6sUg7n2nxfbP+aKJcIv3CfNEu/
BbnwzwHHDzKcpBFTCfTtwOOlvxY26l/PjhwpBQ7r1N3dges6TBWmvmkcQa6vELJ3hnuVb9sARt2j
cReuxTwy/5QeeWpVKQ4lDwKNeQQ3ohE2H/04joTh4c+afTDfgqD5imnRGUmrCbWEMY+UO9O6ESYS
t23Ixb6DgiYOnXULeMvw/MGfCCHO3iT4vrn+h/n9PImSvjNiL8pXFOUKr5gW1QrFdCqz4WZBojFX
iz4aTSQn40VK5DWTidVu+1Hs4sBCRToL1478teeR5UWkn77sfb75UrfzJXvU2ZwOLhGUc7ympHEj
Tb2uAuUDBNeQ6hdRl0KgpkJ+K7mApelvHUEv3bE5iIak2IH/sl1sVhEJkXc1B3EbXwPwG5mrEbR4
T4IVtEBTMTTY4JI0MYywyr/VRUu5b8Sy5O5QfXkXnN0xZ0BViFY8OI9AcozlzzS7Sla/xaiEIBno
xmLPrLjCOpQab1dOwTo1vJLFN2ZjBGtSPc3n5rNm3LyZKqzep+WPft+7pgYcyY+Rp3Pi5lVAvtxo
wzboFUhPzt8+bkSqu/iP5ZuYbwuOEu0AdiMbL8hOlUycXO67aWHXn2XrhtyJaPMxGvHX2gDtlt4o
d6oqagugVmPjm3Vh6lLad/wm1UgYlZvY7yVBnBf3D9SBbmtc3ks0WSkv9vf4lUHvyfuRYglFYorN
iu0AcVxjyv90KzjGBlhIwjyfOeft/2YnlXGt0ocibRj3HP1o5uWopvVVGPTW3Xtn7+xB7oLCUihf
3IPJcGGAvJu/oBCM8kzB2p692XsXA1ea/ePOjm+iy9ogmCf5Lz9dpNQWc2KQwtzecrJ7fRs8Xw2s
vrWk9f8t6SO1UTN3uweydKtBTKFdJr3Q/K1cNPyxswqUeW1xdYQFwHJJS58nKOun1zcVbJWwlK12
Fpc42dO40Vq9xOZ/CQmw/TfdyHZgLuPFX/9X+ErcddPRAlOB2k6ulnKHNSEMVh4KYMyP6a9n7egO
oyvfbzRl+qOm4hG0rTynaZfiNOUrgbkby3XQ0x2tsChri7qeexFdt3lcmEPEfTNxjvZB6bOOYlV6
Ku57DKFneBivtkT0+em4nkQREnqJJfkt+X4th55skSzAWDNh8CKlvetA0y/LtRcpETGQhkh/0Z3O
QifPbD2mBBQDPVFIar9r0NOjLU5AMP1q8e+l67XsJ3lOcoa4zd9Ugxu38lpnQ8wD/4k4OuiXylVA
8nHs4EbkR6oUyIUxVNp7eWpaYTZNE2leCUs35hClZu4LgxxIRVoARGaPsxzHeDfrqnFzZ7AlXdkA
lmHURIlvJA1Cb3ikwdwYyHYUfcOK8gI084502QQD3usLDIcLMh9z7V+XlRXjJ8EcRRemaGTG532K
pxHU4c2z6FWBDvn0rOyH7epfMRsJvg08Eii3Pr6fkFnTmU9pu11Nj1PiNls/I1NwRhk9XTZGuRs4
fDnPv+rnaHsKZ0NZreJMRkw8Mrbkyj5SNuOY1z5LvPHoiz8KsvdQzAJQyNClRAjuJNUx9dhfYDY0
1/3PN7+VDcKwYnxlBufhjp1MiddYLN8fsgQ+0enbft9VbgjfMWqzPcFyoHxVdVnQcTPHRjoygwj/
O6sytplpQzZmObL9cgxbJmuF/nbyFExpRf+/o30A39QhM5PbjD92WfJ1PgBp24s9v/yT/yckYr/k
D83J0JZMADTkjOgNqaIuLEBCex2jNv8OCKgXHQ3bLBtvzYAn3Ld5I1kO23tzwhMy3E+e/RqW893M
vlFmVV4/b2NyOphPCuAFjEPP/SY+Ugz1l09jvIGPisTE3PPsq67weXXyoiTbxK6XkgfDqF6vUKaM
mHWtLzpSlOUakcCNTAY7eKQU+3xELy+JLXbuKoogiq+jkBldo/+gqagCL+uptjdmgoM+1ZHH3xpW
LvA3kNVv72Utol48miDL7zc9nVjc8FvZycb68UnKTUBpmanRGEvXTSCpHvnLpqhjJPF4UbVS2yt4
TdNmmRBmrjGMz3RTTRUeC479h9ylOVu2r8umR4y7zcZ8q0sM/eBBZoS4nFDqncuZZpajEhE7Dzz5
jfY32oYMB4fFrDgY5Ha+on4bFX7XMByTuJfUKBiEzXtAxsV7bBcOxcswFsXlx2pjSb6a3yic5k4W
tBvqWHAza++UhHEy5RTWnOxDLkKiGl+dyliqc7uflQDMlgVkOh198rWBBTQuIAWrLY6j+D8yJHys
yun6bKtlB9HGsL2ax8FFD2avJwbXmQwvvPuCHPP3Xc7r4m6twnY4GlTG7DZRlUaf38vvRDo8SLrP
o7uUhi5CIWlRrpusfL/VXU1xR1gBE9GcqgkEBaWBiI381ZoPuBkUcKvbLcNKziS8rmpFIsrNexjf
2l6HEyW0yx7cZK9bhRvl7b+MJgUQOiiPcx0I/OQlpy1kY10OXr/eIyjm8YN1pKGrfbgBwQ888zUv
8eSajgNI3m8NIbtQx+xO/+0BilJARV787gK4PwMv/+/0GhSFDLVSqqvz70Gz0aUVejkD34YSorNd
62onbxTSG+Qrsc/f9IXE8wH/0qZCsGJUCeVY57xq1GG5XE/HZl4Hmf40fFgyK9D841sBfnbCNcuB
SE99UAjFj/SQFDzDC7fu5SGd9m703sFVyKGlMBx7hcIbX888kC2iaxTVN9x2xDxV8Xq6w6vKPNZJ
2Dgdka2HlG9OioTzB7lP/CJm1P9yfRXAZuUfQMEFWrGgaDWtlQfnTjoqvp1s+FmytJXRqtPs99UG
4xNjel2ClYD/j3SJLOsS0hyDtd73gTvY8C6iFiy4P8B7aBMHV+cj3QQUx9Od4XBtxVl0PvfxdE9U
Wnc02L7jQ227evlDtDg+L7AI29E7qoxmEaW39syv+AjrKR9wj7T7/E0H+oyGIk9hTN/YVlcgHFCa
0BmW63rie7uRHYr8/gCSOMLoa/8HCQiXtBjmvtqKUTDYl09QB3jUeuMYUraEW4+Ckajvj66Sr9kb
nIId02BVVnKa5KcZTd29YSCpBIyRc0eOhz1ysDm+D7tbyjXXyc8tse9dBkRzUa+kI/adTPrJT2Qc
fDdoMS2Nh9Yx5lKcEFJX2SzULCg0l8gXhl2JvxNDNZQ6ebvQ7Q8MZ7qHdw2P5EJeChN4ovm074du
UhF0IiFyqcVqa3HwAGyONS5Eu1tQzTFnOcIAdiepxDOz/2W3mP77j0CgqF7ZDg/sTJ/wReXXQdy4
ZJO9EAuveLwCSq3OPY8zhSl/BzBh++hDqA1qlWvl+vFl4HMkqTkpCUEn85YGy+kTSZw0F7OHA02j
HRIRxQ9kStFiHAsSCY2I1RD2/8F4piX9GMWH+CfhAqKl+xEiTVusaE9HYN1OW0WA6/qUxV/8nBHT
oo1+Jt/0K+jJE2FkJn3DnQjZN2oQ+GCAMN1VMS2Sas00tYt7uLdIUSBA2ZtkesP6Fpd7kswH21Gr
hw9zi81Tiio7JYsFwsWoiTaJ4sJTEvZsX+3JgQFUq8qxmLHM5Gs02w/4AknllK8E+N+by2WnFOJb
lWSJTuQTxPl3Rdctg2NbFhnSGZCTZxg6ijkuvIz7mUjauv0hQq73t0MCJB/xdxvIdtZQR/kUtbFE
KaM14rXYoJq/HPiv8/8KTB6BlogB4KmoSsBRHUIZp0TqP4hlN+GiCQ77Tf37bjSzTIqzEe4To/GM
PEYIepfZBMi7UaXoS4wN9OCePoTGInXwN72fdT63mgSJ4pY5YRThN3ajVk0QTlhnWJ0QYr2iiY1M
l7vBwTdGcJKy9/vTihN0uroUVe38bIu8VURNi99niCdyFSNZ40mJZNXhofiOZj5EoV/7XU6rWaIs
oXxu1lpL8KGfVDIB9jeanpgZCrSvOfMcwT1lqDpKMpYOO9YCdTeu5Gnrm9md0yHrpJ4gmji8DVTn
OkaZWvxQMdpC6NtykjPWaCyh6GFEq9NhY4HDbawsmSGj/pcz/opzrmOMQU2166H7ntkdl0EUQmYz
P8Oh61/PXYZurJlZb/sOwNOSmtPhsy8MRR5fW1yJA06FFI4idneHTusZjkaoK/4uxOI6KVpQhCWW
WMyAKg/fha6yf3dfcTDJpY+atCYy2Km/2hcqNswEuH4KzU4GoaCJmQgIr0qsDGRvR/Y2M0AgZSnM
FbeKOxXiaX7TJPBM1CVqzvaP6alR2TQZeAIyaehIwii7iLlaRWkKsaFjyIgQyJ7MZy1PfvegDwvb
6z0CowLH0qd4e12GkmNJQgQDZeMeJ7rxyhqsIkGThQWXiq8feCq/wSJ98Ey4H6OLQEsdgoT3uM8N
UtkGtIkuGwdGZXzTKmj9cA9zR4f719Dt82Pq5/TWbJn6ND7uY/1bPkipo2Rp5FnRFsAUHGakjvBm
orUYd+UUEXZwH/s1JhzdqPywszQuiFTCKuG5gBRdVRAMNB11d0ej+v1Ov1mr0S+5ZWsB+drqAhPg
5FWUVUtl76X4zxlWWHhWIMU0nanJe8H/dwWdmeqWb2HvvOCwERSw9BS3IwWqR250vPiXc5lsczoN
3aWjyjqoqC21t9IaeTEs2dY6S8IHhfElXiZ/I5hEjtc5wjgNA0ruXLhFr7EFMrJn/wS2ONnY5rTQ
NNLDx0XJZTOsjgL5q1CbL8pvAqrBNe4z37tqVV2GVGQx11YwzrsFz75r5nzXHdl5SRSKGwzb32ES
NtpWYrGP7Uwr7hnIe1KfG0Svf/jN9SGp2uz8YRNd/bt/j9CHvQ0KIWQHk3v7WFFLNRshXXiQeXvS
Jzt1CwGuumMxdAJ7Q5j76b7crOHi2fQ3iLVG+jsJf3GOkk1SW4UPmC/BlDRxU86Obn+bwZsHV9md
Uuv80S2Fl1JHVNmP9ZMDFFj075ascT3LYRSjgeasQVhHTFIClfVI1QdNJEToRjErkusRwa77Bw0Z
YYXKxHIooPwFGmcnTg+1RwqzavMbgDnAmukkaBBYFaLm/bxOsVvJjlt6zmBYUkoGqvoeemjX9JPU
XJ13NO2dRkkafj2u7IrZV0oTmji5TPM1j1BEwLObqrUHbDoLyup4W9zcp8jS6D/lEEahYmWlBc0n
scg7e1iwpctFt8REKzjZPou+Qf0afcLYZqt2NcgkDH6H/sQrmMZDtvlUrGAcMOMccbGY9tEjcHiv
RwgDAsGdTKmYfGstsswJuD/9KM759LKQ9LVqlrLt57AM/tmbA9PR4EEOQ3t1BMa43nX0R36vejQu
IrLl4CGfFBG6XojpMZmPqweZfWMAZqGb4t4nabsgWf3VICffsT1X2dzYEp2+Ya71BpUbDi7gOUV4
5BRrVkLNewzN8E2YLQszal3f8bkKyGjDAKG31P2h+u8C55ngPATqVtGzbwkup8bSpDRQl+rMINcB
lFTqZhYJDdaNorBbDZCmFQCfIzf3ruAwZQxBve+eCnG1eyocn371qAEfCozP95jotC1/HGQ9ct6T
f2QqmC2tjIbdvKRQmURYf3JxHyJQQ9CgGL4xlzsIL2xOOWIRa5nDnAHCjqwhy/eOo7mCv6fY/Ztp
SLyEZF1HKid4E2ZI1SMWfUXX8TjIgAoBndRTwKbVlavqelDWX7wtwqjs1CELoKXBF7PP87eH7PJV
8NeenLtt2WfhbJEwzRZ6PpkhQMBARw4gb42E3E9bGPO9FtjGXHPMjSIolTst1DDqPgE0KM/jqGUH
g/b63aAie/IbVvN6LdlKvfCWyXtyI9unnZTbVeF1ipjbmjt1gTsxEIjWTcpSwn+jsty8hikNuWM8
C8XhksSHxLttKHljOTW8xRzFCeOVqsRZjcgnFVyjkOXdoYYGt5op568xiF0WlylxXdHezabK00dY
KoJV9ynIeBGX9dBnCpHTYVgmIPwUuXDdPb3dWTyCw/EawQt+WEwYBjVcAHWCIxpSWDFICfUMjPJK
m4K6UtBE3SEtRz3or6sbVyFpqPLCVf/4ZkTGMnu4emwVqNOPTYKcix5w6evCrIrzvRbBXthOdf7U
5rldGwcLvmSIoHgui6Y2FocYNN9GVyB3XA3iA29WUAI+T7/6t658uRXq6sgn9pBfh+bpBAShaJ4n
GEluOnNa63ZPD+IRcN740FNoAmKAz9/8HGfe6nPoSqSX2ClfaI3SixWhIIwKRs9bmBRv1fZZ7oH/
O6orVKW3GLrhsfH7EDlayvNVGcNvPRxhD5sXdqI3YRuJhjMQy2hZDb+PrkiwtK6UnnCfVT95qrgo
3ZDiRKJQ/+FfW0/4UMyS/Jtx831TYLXHuNSi6W0No6QSS0IOma0/ucy+AZ+1RvJQnvP2g8xgOdGi
MfDWW9gv+4aablEaPwXBjNBtWRjeslJQ/l0svSBpzTkoSHuGcUCXIF/WbJGkGseRK5gPwsUeLU5G
PPRTFSJz4TbMR447AggD7HCkaN1zGEPBSkB5doK9trGUY2yskhxgd64uKAK22KFdTvxVdqpIdXOz
qe8DV8N93hquQ4Q0xAxPTU/+rJJfqpUbrSZW4BWCd42ibzn42peU0hp4XkJipl3kRYInl/Ud99Jb
hs7MHE6yXpMH09Thyfb35LEqk01fibM07NoSlv99D9PHavgFkLYIjGGo4Bbuic5588ZDpqwU/rE3
FoUiUpxZgvsSXXsrkQaVKeCd1hoTEy9eL2A7U/GvsI8IRg/dMVvQayjQxo1bZuMJw1ssQm1kMSi1
crMbbshF+w68CsJOoHifSSxqgwS9rK+bBqCwU01yxnjIrMu8eiSGOTlFSQWPhZUDe4XFKpEcoLh/
hwuW28J7OnuSruMt+dK754OSeRFIwHY2UAXKD6vFvOZPt088A+FD1XMYOtYuF61sGigKA6m3E3b8
WhZBeyCDOk/N2OyF9Vj564ENeF3bnhCrogSCmBShjPdVDX59V47LDyTPGuoikqid+bQwSJEtyMgh
e7RvxZtMq5AJWn4I1Okn5USCCalLZCfe0MEms/0BADcM1anIumlf6MqqamvVl+tCbZymOLCtydzu
MniB64GMbBug6KYAj2etTymgyljaQQ2c1FrGLYB6yq1pH7BNB4+gWqunx/DP7q8J52thgGjfUyHl
PAhd79GZkXn535IK1ec4XTWss+A+Jl+3NrL/FhvX01Rzt/UrBwMW/H03F5xE9nYBfKfVvcEuz24/
K2mnmkZxA6NkD+YbAcPzFYkZ4jg/v3i9YLNsd0ZtUqyJcYMPWiJdJouQc72gx6lwVqVchPuB6OPx
LkEsUaqo8Mr4GFMPW3kQuAxcCa1DUU05lJBMml8UR2KFyHRNlKG+TyM7jFe+AQa1k+tU1t64Gqpu
Po6LiXhGub4jiWEmUHugTL4ny9AR/abX11krID0Ybzaw9Aj3V9fLaibKzrwJD/qalh4tOxo1f39Z
1+KPFlz18ewuroUKq6tfkXW2saNebLwy/rpSX3QjX4NNWUYHAo4VOcC5GeRJxC9sbcvdr8u7mOXJ
YF0ynKpIu6S5z+3kJUc1JTD/PKxgHtNOp8sOppgQrHc5UM5xWy20IDp43OJIIpyJYlAhIgctpcZb
eorg8PcUC0tAvki+uaD2uSKsBaLVZbVjBmXkjvnEBMMEXPSueNP8QDN+QiAhCgedI4jZXYb2gd/t
Vg9P2m/v9rXpSgS6x1+Kec1WmQvV2Pu+0KuKqJpoNeBJc7wogfb8GfqvJw3Vf8UxncIarxm/yVm4
h80RVymSWYho6y8UXSMLIxsowyuS60Dzn+cvc4uapLd9z/ipzz7nbTqPjjdbTYPRah1Gb719TWqo
P6m+d/iZuCvhT7OtDxzc9AmAF/kbf6uZSR4MmPKu6foPSHCY6cU/piMqsL0ckcjmFokbb0m5sIeK
1oFGxWKCQrCXQdTTbbmFlI0FGqOAjJlbdiphKUCl4SR5jQ8vnnsKLzsRdqrNWWxnSnv74ROO0A9f
zZszPHfEQLueuEq1CqmgkXAEaSZakVpKRQeW+Qv+zJ6oE8h9p1128MFWMWt4ejCDLfLvxG7KrTCP
BRsDHfcMa04TwY19Y2jBRHbcCVmTwgt1p1Kmormw6XopXtSxgKrim7ZZaJPs+iF6UOpqAwqO+soF
cTEG1Q9yzNj/Dp5ijToU8vjWzXAoZnUPDueddO1z6VfXIzi5W9Gzfbf5w2OvQ6dS/Nz9cWVbuYDA
b3bKsGHuliRaB+U9Q0kmuWSp9/s7xnYy2ofZamXzBEvBxMaiotV4HtmBFEXpdSeaYjDCQD6lv5HN
2D2ndJIgotsJZ0eqj92LjkLpXDI8eAhiEzx5Z1vedARiIJtxRshLPox040mUwD/0Dn6Q5cknvVOi
K2y3c4iBAUmPM7o27Mv4oInfpwW2p7043uf5SMjGSuOoDF2h/k5qopnfQXz0pUSzEQK7OaIP7u2t
FdPdi3FaMnuwwqke7ViG/pxbbH0JeLZNa7mT4rJ8rDBFd5itrPtbUoY15mkeEZGKg0fg5lTSjoSr
zLGqefRM+zO1xqbWpnYQj4L/fsfBhaFPot2jrKpoeABotE3A3PzdKLoZzVhth1m+oN12ZRvsiCO6
jr3UfCHpAu+Fx87QyUzqhV2Tmfx1NpX0O+jY1weTPcGnFT7kwHTwCyMffosvxzNn/s29f/K85/H/
iNNYnqpNTd1K46UeV4ruHXkLPs9wCsUPBdi+MOnsL0D/EEcJ6wEz5i2MsZa2Ux/WPlJ7sSOnVe5R
aJw39NJRAKoPDNv2168iA3xepq5Z3Kaa528UNr29zqypoiKg076Yy8s8Z5YmUNYIn7aUmiDqzZhx
MaJ5UF21b1Rm6AVnpB2gnhtMy5zYkFo6I2v8duhb5s0ta6Dmf3sVBx6DpTgCoDRDThnLswc/rGQY
zceJMj7b3jkjgJ0uTiGddfXDSdMc7960RQQqYfxKaQjhup/zi/tN0NbJQI9P/SyJlyq+Ye+UOMsM
Tc/kzP4GBGdo+1HbqwBQs7vTT8t9pyN/B2TMOINAkAifoUD0hLHtDn8/DVH4ojucrOpp4VGA4nEB
y/Lw1b/Uv+I1mN2g1C4DO88woDL+GTmwE5RjNWc9ARpHu1ptgj3SlruDg66SeEMJVo995fN+vKGc
zmK6mRi1TFERxbjAEJmTHTDV1eVsDEJDRT8WTBgP8VJ0VHyL4bnaGO7VaVMcU6l/0n/ux7O51DIq
j4UTom4xvuMguEQUpbHEU/rzPaBpbxwF6XTf3qdilqmYEYSVqtXkSsW/ytAX6vpZbULNXgQ4otR4
mCFRC+AhzsPcMGttfaN0+1nv38WjF1cYX2ABD/b/QRNp8EqzZCFlhjLaG4fpSlSp8HOkZu06t4es
s7UOXchXuDgjxPQdIIvToMPpk8nTk/NPdxrcZt3JM6KHHUqwtH9zMYoLfKp2MomhGlcVus7O2LLe
EiYMRUTLwvmObv3qITP5XDp7UVkNOujZSRwk9rQnJSka0yXtEJsVJzIdHf8C16oCPEybKIKYRc9a
a/BRWGy8hqOcK5NPdobx/yndbeVcHVaq5cSkhM3IfnoVw/St9VKtaUKcMQ3VC7gog4C9eXTYr5Iq
7yeck6p/klOPDAU74mmZ5gXTvqs1jtb0BhrbdS2vLnZAusyd04GqE9nsGgfi+RVr5KKwoWoED6oc
+88pzJy4MbEwR2zyJnenUBqHtibFYL0zTHlcOjuBLbUKl9GTiVoE4AQWB7XtD5g7J15TiXVhiBXd
8UpWq0cquEIIoQ7bR+2heZlpFSoDDfpbL/VdOMQwTfoEl6y/B1orsdpzbc1/+69rraP2oZ8Tw/Wj
SmFFp5yHSOj7Dx2ZgDvaMVCBEmJCzwP/7XSTQRVVlOIKhlOV7gxtClvJEpK5R8lBogRqXxhiJ1Ek
0Ni7KIIMchUJZIeB3fx5gOmBB0nrGDvgjnrS0dlcSaKPIfsnMd2+xugdoELEOX/OtONHm/e3rSiu
TU59SdkJ13HZrUUkL5HQ7oIO2XBoA22RVX3tiWgPUjmjw3ytovEtSp3SpENebpP2FEYMHg+pUsUh
zH9IzYC945DQAhRTc3z+FM1O2Cd2uJHw9FmeTsxTG5Ra5MC/g0L3+21niN6l7X5qdfQv/FyAse04
02l1WuFCnGukFD39iErnVh5+hgScFsZ/j0oaBGmerIeIZcxW8hAnJODFHtXKw3dnSXFGEQYaF8z/
qRnETcT797o4FpXf2S52OgtZTIunc0mnyiohmk/5ynDVz3EOyiMAV7KwsTE293TCqXaki/5xtU4n
PUZ9StIgKGlgPCHtgyjbLKXICBL1xVhNsjY7Lr5yBrPwFDIvKrDuEDtDVTG0hUPg+b6kbeSlmeuN
aJ1eN6xaDBzQY8V/AGqYFU7GWflezCS+cEzEse1QzItxGri48JkeWCQW0J4hKceRz3xdJLfx+Fqc
uUABKGTYhw4zUWyx13AriEydx3bhbgnVF8b8/nTrFPxbh4yvNOfe0toBsMOHUpxLRvCUpJVrjA+Y
YafYksa3G+nP6I5/tl8qVc1Wz6brWjjPsz2AWx2KGUAqsltfybjPo0d2K3HOkJr6eQ5VTJ4v5jkO
L5vijpfBuryhM/eQ8GOR5DDFtFje9c1AaXUmB12+n3LU9jgTV7oen+0+5xRrssB0YfmgzIuHIleM
puzqbh7U3Xp/fnwBRDLeuAXzyQITA/roz2b027mYvpRqhlx+qnb8XgR18lgjrl50EkPm8akMYOZL
6PKugkIJ8BOmjBxAGz1kk8Hm0aAy/xNxK6zua8O7hrl+YyGQu6vv4lORHGoCUj6xJBQnyMcjRWVY
odJJvTBW36168OOTi5eMRvlz1K9ffpXrZsa5jpsWE+pVIQlw+v799N/BB3b51cWDRr0jxqzRjdKf
ZzKoseucAKPOvzVpbCwkS9Q3Fm+xhuCzpoB1a/59MFz9S3n9X4BQlk917QGhScymNGCTkofl5TBE
XdgWAe5rqMdKV8TpnVaxs5N0NImV7MeA8EpAsAHjUQgOgBX8yKg6nLmRZjQjhePdT41pqZ+VLopQ
qMJuDskfHUf3Fau7aFjM+K8wq67d8SwoLWKtJbS6B6IHKVlO3XYoXx7beXbWAC9S7W8AtP4F2peM
k6SVXZ1+3NfFZX5NSHVKSNC7sk2Tar363fgiO1oau2mvdaOaXLWa4j5VhykO/ZFsy5Yd1xs2LoOk
P/Wi7h+r7e9rL3BbxqMaQanohaAypQ1mdFfLhTSPsCvmj3lx2Vl3FWFM32hYwVmCZDFOty5Rf+rT
dHUno34+jroXQLZ0J1UMRrd8mdha/Tp+QjEBr6LgtQM/9nPKQdAmgxHzyt02PdjBkzOqynEgac8V
3y5FTo6j2P+CS2rr6yISp2pYJ0cVDADMIU6VYEHk03rnlhuaXwzZ7SUQh+asL6VY3xYRYuoPjXx/
LP5qs3L6tIQMz6ut+Z3GT5Hi3ksX677S0XMcxZ002EgIJgNipS16CSTe1peTW1P5/HyVVO/M22ef
annKZu6corx9EtOxPr99/DONeakwMrzkgbS7Q9wXESRS7SnMFX6nld1JVwO8N7kO2jjCL7oRtXFk
AZB74D7H7exesqqcdM4SOPLs5Wpzg5tEKb7Gw66KlkbCJzRYR1UAcO8M1wc288WXye/U/f6uXrHh
bHPiGFDOFSgAe+av7CYI4dDq85dgeWhJIYpFZk6thxrrJ9S5N2sCALVZJbbVOkdUaXCHOVmar5M0
L8mHZYhn1+VIrDctrI6i5a/OqyHbP2+4l54GbADLAOQIZw+2SQiDKjCFdwXsfBAOCmrGgK4zsDLB
Hz8NA28hHlxxt3puzarSZ+FtC1p/UkMfX3RFICkcAa2iaVE/spQeBlwJ1iC1PDOmhU8wPH/IxSwd
syPvz39UPKlWQ2lBLxhfFPfYJOmSEzQw8TTs9C3wLho8Xc4mqSE8gqrIAI6S+TgKvxtlho9OxxAh
Ei8FKHxDxrk3xKJp5KA8K6ErcKqCdJNTwaWcTTEobzogSbmyJD61NaJYUO6pzlW/kdktfY6RhV96
BrAxAfubsKz/TeTtKofsL5W7us8fA3i9q63xUpO1SQcnLTtOcCoZTngCpPkMZYwBhlU9pDzIXU4e
Jhx06SiNDLKi47n484GUmMRhGrSpP24G8uYXS+I0i2YouH3z5OQv3xnGi/ip15UeCguLLOBCHj0V
AJFbayFf71xBh4jV0UdQW3TDdslQUtl1RAiQrZbWdNgrYOkzX0IxSfbzzX40Wp8N4aF8QQDqjdf3
zBTpWxgYly6/MuGf4Zlb1lsDhJlxOLYAfl4d0DYBzMQ7siHwTHVKvhmC1UBg5egqDrc3crvtcBdJ
wp+Jsjl2UWkHf+OQi72XQxF5aazkHNhvNFhrUX5Lv1Alch/Bszk4HZVIviZEpqZ9YdW+W1pEbzvD
qwelRmxl0BBw5vMHdMis3Cp51Iz+Z8JIvE4SJagAGVTbmkgIM7iJG/IK4QLkShAbbIfv0ebec1Rg
rm8iF7g2+Id8/vjVn2YFoHGgol7C/dzjuj033sU/mfqkKtvSta5ijwXqHpMVS0kL4PyNf3U+HaIC
b5YjuEYGltf9Ph5AJQ/Xnevq1GaDfeOcJJubP64SamTui0aF+q+Lk9nsYNhINRZ+giprbGrjqREJ
PX4GXPmUSUA8eyELolp3vJ8cYav4JevIPOk56XzNTqNcwOJ58MdOLgCnC11pPMDnLBzCLKahicIU
S/8fv65yygps/waGPI7GWqPZc2/CDrftB2angscm6oovLEWJfak/cN/qDUcRwEaDEi5CLJV6036D
LINSSWHGhhQFrnTmD/6xhol0cf3RPxeJB9ozTymV6xWo/+0BLOyEgLdahqF87bnBpUkoqh0c5HxL
BWlhQvM8rfXfUsYmA7sLhDH8StiXhFtxXacjtf5OZ9DtzMR8kXBNvGP+o1GsZvYWmiLxuKJ4R5kb
s+8i75vyzEGF7Yb1vry4so+HE9D9+IUXuueV4FNRQ8FMZ/hrET2B2KbDqmTfB3nitng77XAKdSjc
WjHEozHUsUOqYwQw4k7OZCoCB8YaxotJ+uPOE6bAjGyDUKdJo5gw7h4DLIghWA8lFk3sjiouW3Rg
ifAkIm9Es5xxoGnFewXnC9hEjOmVQUImOQA4L9I56jaIuABEBdI4GAt0Eaq2SQu64/yhpQDPHg3t
g4T1+DYO7XImE2Lq1DpOW4WhgP9zjqakxuOZfZUFaBEjZpqX8sQG4h8UFyuLEOlXaMdxWI89IXIa
/NivLpmrm+96BgBRx0thTSv4izMywMiVwUsSmbeZt8TzfwE94dhfJPiMdKrdCLKoV49hJdRRt3Dn
4XkoGuuuW8AjXu6pz/MvyX475tYQoar4viEqnpEpJjhNnbYleN2TMUdMhXBNxJ4fZ1kSceJ3chMB
0239md42joieIiqziI31nA/CAfXs47l1L8Han5MiyA7U3tsx70Bj8Di5aoQL69VhARMnXQfzvRx6
Ex0qbJ3Mb5pzuo/MBAcXmePl7PVfHX2rpCtMNGc1shZqL/JRGlf63qt+Tx69sEMfjklv8ynp7+Kq
9CbKiGl+N3ZW5at6/LrhFiB4yavK3gQ63aSIW9zSoF62r1Ogsz842REFaastmAMTaKVAUg9mKpJ6
FWIt5Ubr+44wEnt/DsJCxF+yZDPBiWl+od4G8DOA5g7loGdhk5CDPWQyZ2bW75QyJCcTCGz41dct
2c/X1eKoPpUiHheyJN8sIQLZOzWEQ6S7nFWugUq41bThG8ckBw79yTruGAKhfh/Hd1TeSrEA7Kbw
c5dS5+GB498Fius2vgSIqBDozVR4c64GWa2D/Hhb2f9ssUqrdigxeBlYDsuwYHmpxyQ6NRYEfGBY
kndmfld+3nqsXOQOsUMkD4AiSy/N4Mqxd0MCEgEds5noDpGNKCReMa6yosEfItIe1wq8dvlUgqlk
91PX4Yc0kk7jC3/HI88RITmdyeKUyOtMn564T4EXzaKBR9nxjycuL7ClW6wHyhPxlESrX809ingE
09FBk1HdVFcUc4s5X4BPdBT2iagqZw4Wp+GMeT0AuLlwf+3jJYWc31wBRHStE5bYzMT6i+xlEVgZ
CuJN8dH+EXIbz3OBIeGKrIcqUBpPn9ekwF2UgoXMRFsJYOfMLCyN+JxLvraI2VkNDMAx2GQ7iId6
9iZRcdrflPur40u9WPXx35kemW//esLdc8CZxGYqW8H+ZQuDIV/jbiElKAmIWExyT6ARwcYAIHhC
pyN/jsVsYlANMw/6xs3+Lgk42SR1Bx1qPRMSKADjDyWQNzv6ovofTditpHnKqJYL9w6rl79rfXwT
zAosEBK32Hga4hUbgnlLkmRXLy8zAUCRni6x1F87bIPwXZNkrZHLPNKbzjyZXnvUF+ykofOfHv/7
+zQLLRdZlKAAaljjfT8xwi/5Cj0JH9we553dPMaFhlXihb37QrE6uUgAB/t9N6UwfkX0nPyqJxyl
YrNAiF+y9a7imwWp50OxSDDnQN8L3dVolHgLIPoSxtL5GIFw1sVINylCFlUHrNEchXJWTz1Be4Z3
mvtvkDZF3ZMNBk5dWzPnoi2Y20RW8gwtP0czU/BEhFIfQvvc7fd+0OEEQ4gLp/crDf4CzSFLpSVn
4LBoSTSiu0WJ+HsEIRdIgQds1BPTcFwR4Y0fplxB3CfNq6rlZEr38W6Not9KVQ2r9owp37pgwl1N
6UpGisnW/Jj9wpWWOXxxt1xk174FvjhBk5e0uuHKHDZK7D9g1RzWWQD4kWgMDaXgFqDdzzlkvtQM
uH77hbpY5lLhNnd4A5loT5FZ/lp8LiLsUtnXmOo0WW6kX7s24NgxB/IeACHd9eLE/aA6OvZlk9zA
3dtkJ+Jh23NjBAFTIqjkrkpJu7l/EPAIS13Yz7HdRw8HARCjdBG7LWXG+fwRo7NVPEXhW3edfx6r
iXJprxZsV5DL58IYbijadrauE+U+ZPJs/EhNUoekWhz7wkg7QxGFawIxPk4yGosCKknO5rZU13MF
7Nt2wnOthsNwMU0y4aS1vXfXk6Rwcdbz6K6b0TlAjkQYLCFYOUebPahXqej5nrcgt9WgjGD04Lvc
TqRrTfiYfu3sTPsVNpXhjITgbgUZ80pd8Tv32pJ78/qBGAkTYgGaNJTITt5nG6uNUrCsEd72peFO
Cy/FJ9R3eexFe6xb/ElCKB9sLIkJJR3SSilKe2FsAcbfcQ5qBjn4O8veX21PvdoD77oL/tDCuctn
xRg32nblPchssum6ztXdzHCxfQ4RNxy1hxC/i8UVNg9svms2ZtuS9MBtWTK1niIpgRNc9RWEPDOB
1Zv7ofozsBySgrB2fDewtHIIgybnTUop80MzDkiEUDum/ibdwW22Ky4nprbghwMK7YIfeYAFY8v5
gar8/9kwBvCN8vPFhyqEZXCUH9E85842JxhGEdeMI+EI4qAbC6dRLZ7GkFRK8Wo5OUcu4Zu0dYGI
+sNouo3iLvlvLZmjQ/xIND2oKKYzeG5sZ8KvYtwMCrP6b7FUgjBdmOLc93mVNas6HUdAaqq/63vq
1s8N32m8j33/HZpVsr0Nulp42xv+YBIF6x6DNGsZel4gbC3IAlKG9qWtlxWuwi0nV/Q/CzG5n9Su
61owpzZTviVAb9A5j7WTBQdiDXlNxxKiNeFIOUHrvNSAAh5kUYKdNPjVCB5iC0nmMCZujr9RXn55
xqrxlwiriXvGrSDCCa3KAuv3vfJkVXokb/AfZXDHn/x1VZkASll+WP5i6YxfG9vcVY0Xl/xepPyg
xiZsiUVVOntzPbFFLCDJ5uhaFHHj6r01DeygsKoeFOB90vjO1o6oLgq5Wvk3Gg/MK16xu8Age4qu
HQMxksr0/Saww72dgr47nLHVgfHWfgAZl+bAE/Q7qkdGx3V2UufKrFHAbItwuolwwz8jAxYiuK3a
+QU0DdEd6Q0kPWnXGqfsy9sPeKkhXY3m2cW8DToKUL/IeqOM26aGsxlRJRbON88sZgHXWnvUsgYf
lnNGYMs+pdfC8+LgVHDnm40zg6AhXGp+F48PsnhCRMjVM4BkC6+RDUQHAOZ/Invkhnd4WfYSU8N7
CYNr7GQqlZshAMtMZRdgeVqPXlPaQ4/grRvGwG+ILjyW4fMtonAII10dnnx4zCaOFy7nQ+bqrZIe
oOnHDmvilbJM/aOGz+PxEEXubSqRqWJe7zZ4ZynhULFNja/pHap4vNxGRmGhXvNrT1ncuUlbhcdn
dR41cOjV5R3+uOEv6+KTNXgdbxwSz1qvTUf8C2aA+xkjO0YWDPCguDGf6i+QizLyitFLUuHdtog4
8isgG+kHduVdedxlHIY1L8Z6dJv5MqhUIXrlXI99me9ynRIDQh6qj6E7FQLn06Hrq6vkhpqLVqaL
GQG8S6NhoN465YHhb9b/mWBROm5wSYfAG44HbJocI9okdWxV5JgQLxHHk9s0BJ6GptqWVLWK8GGl
VKhA0J+hMgWIZZQhIT5atx41nDIeZCJIIlJgqOJ4Pf1xMYhQlsZ9x/BKy7H8VqGXMYbCtw5qZZmK
5EsQRWrMK+BdcFGAZkCGnRQjV1KDPYpVIi/U3QtOwS1RENZuBE9JMhq5pRDKTh257Vb/Snr5R6p8
MBXLvdK3+9Yg8eW0POKY4iQzfbcgveWhK2Tlsgh7sEvD2pPYaZKcca5SQb4u3hyhTQ9/3r68m48g
J1Muz2S0YQHTYveuYf9eOXczVEJelbVgymqnh8L72xZcZzy5pF2SmMLf2tXdFv+oMqOnwqSNAdNJ
m+GNG2q3wjya8I6IXtjR6GShwG3adEdmy0Oh9NJZhk0y96e8hAjaKE7dCToP94k7IKoBg3kLMoVe
CSIMFaPxtHTcBbRLp05RSJLmd5HwfJt/+oTPIqnLxhIgnFEw0EDQCAex1LM8OpGFQE2lrx2OZxbb
1StdNhl1mVwWmA/eHBQe4SJYoke2LhUpge4Z2RKJmSu30D+KYPh/tsTFvJAzjdJ1ocAtUGfu4KRT
toyCMZ7QL69weDrWuNW8uHH+otrNbDAa68bqwRKj20I6r/F1Qo1xt7UT1ijc7PJzEKK1P5zeesK/
3qdxhvhZxStaKXSJUY5XSuZFKE8HGbveucvBGMihSYvqinLxeRxEPG6D8Q9AhHYn9/CWlVH0KcY7
WhTWxE0TLn0ojN9DKDDHCBQX2bALMELpWcEUXp19cMPbXfb+Udwx8IROOHp2gDP3bBNs/GH1pk+E
UaPk9oQ7O1eT0cjpjVEA0KMMivgNZk/gtKjcJoULw1yr9WfXvkQsc443zmHC7XsdN/ASiM8TaN9p
aO7wlsLvfKfejnsvehYuz2rVRWmS90qZ8y7IbyDM6c7KguOwHT+oQXGiYshCkvpv6O+k/j7cwsB9
AF0bioG2hduIZXV7R9QUSY0Sjh2GIs6zn59py2nePy04UkRtFM/7RVdQjIH3g8GSkhX2j+YGJru1
fjUi7r+pnqn8A1x3cduhEpzoIYUBtWsAVczi5hJk001aENKAiPysf12mlphkcKEtvUtguQ3WAa/n
fyy5nO4XgCQzRKQ4y3Ui9Mw0mMiSuhx5Z0xtHQcKgedTLBxq9c6YEHIC/iwXm8LKPajgSUrE8vby
l1ZVBb0s53/3kjJQcs7+Ztoc4gM1M7bDNM2yqoU84T2XAj5KaRGCtfx7nqpcxw0CCxCn768DitB0
Y3brmM4vONRweFIMUpvqEgIqdLCPAJcjDP9UV4KyVSthrmgBRS1fuk1tmK1gAJ7HyKTMMYwMQX1q
U06G789LLqgqE35lGQ4Ri2s4UIaAIahDD8iq/B3yNUE4Rbu64vX/TrsUm8whSPrUg1VFQ/ZF8xp/
Mu6sokWp+R2dxBm4NOcSNJwV3O1aJWn//ZMQa0KXS1xiH1ZUMsVN7w/OQx2qU685WLD5sTKPAd5U
YCpgUuAvQufVJ8BGOV8r6jK+2JSxnB+OyJeznK8OcFP+06CWeKWIUeYz/etpVCjfvpLuB4qaYcKh
w+Kbf660V7jDzxr+oVo5UvqkVAU0DluFWW9gcMKTBLYKYap4zX+OSd0Pc1F99MznVq6e2HQNUSpR
bKd6ojgwB2XGBb+bQxjy33k4Cg4CM2XzNgUjvQdhTZmweWwe/zyVagWK+DqKlzwxoRvqQl12tJ/l
73s57srFwkOuPvguH8VI6leHiz3Dq7Vdm9nzN526CeCej53HNjIiFhiY9KIDtSe2eX3gqzJyF0QB
t+s/C5N1EGItlUvzhpcEWBI+oMqqm9LOyn8dLGTXl1/JLV64kDy4w4hiwV6DtFG49vF0UmeUAqgQ
RjGTx8g1hfD12nglT32ovqT79GySWxnov6IR0XC7/IBBsxJJYTfJLp8H6fzqKH41bHgAvDTejGyq
87rGisxXXoKtofuxD4IM0qCl/TCyXd1Hak9WV9FK5rEOlQFO5QLUcDLAHrZQsnnDriz0YpQdddjy
6KcEfcvOWzxwi0vnm19lgrfF+lzmgc//E7G5vJbRK5gN6wVz7AjCiIWLOVsr6+zhfrtTwY1p6TW+
TYDfyl3svjy+3885QHSEM18tbZLOONkolfMEz3hxjoFjRNzqWT2tXgWEJYPh0VMuPPJTZxJS3r0I
D0GSnNE43VaTQyt6aLeTsTQV7xg76ppv77bi+0+Km1R/OSmym1Y9V+TFXuSQDhPEOPQkt+oK4yLW
01sBiz5b6kjeWitWRQGHPo7pcxhzAQTGfCxqmvXcOqRF0gXPE8eA7aAaN1124h3VKVx1YVe86nt+
z+DyJKthY3f7GOTkREaKyuDt7MY6urqhZj30yq/Yix49EqUVFlTfcQ3R2ilBVu96FcZGm8/rYPos
+2P0nvdkD6YajQdzMqkG0i8Amk2JuPWgivDCd4+lcJVmD+LnOvUW29m8WfhiyKPzRLOmlDHU+/94
avf8C46AAxvamr7sFNsouF9NK77pMW9UHjgOPIlb6ZcCgxH41dEt+/7lKHiw7CwytRPNAifqG2Y+
e9YBHhEhG2FoBJNHKlcmBry6nvaP2f/uaKRgwfESn5CQgcbfGDBJzflgU6i+mp3P+L5VOBlKZ13M
f5LmspYC1tD79Jii+dzpLcpMwfuWBKuequhvbWeQublIn7rObjpKZu0yKuyNxpUSu+Zxb8+KbtNm
0eENLoVUDEfmg17Ym506N/XmEOM8jqnSsAYfHcYsFS8Pl3kZm59uGYV3OEgkiKWuWX1OzvS0zrW1
GnDkDAixfInblikk1YwtEaqRsX7Luuivmr8iRn7whct1noMp3ojON1uDiYt4awCwr4yOxV/Bj84o
x0S7suThaGRF5fMBF/1Y9KX+PbXIDUqgoae693drtIBpoU8at0tjlviz4CfG6sYUiazxmJvq1aD8
MfNg32ainGY9PnfQ5xwQ3w+Kzyu9bDpBsgBDT1Fkssc5Os9gGW87CuBoBpN5SHmEm8odepsKltOa
0wODe1iPFguRqDe+zgBMLgP2VeYX5z+kdxwYJqIYpyBF3Ul6iLzjfbbEHjZ8X1pQjcQG2eCEBdhX
OaisV1vLVpxNc2xCPANSxEvgvBc8yEE0q1ct2UkDKOaxJf7sUrRzShSs8XdFvb8bwP7onjACzzvy
aKcOvBGq4JEBMvMVBdIFBg9y6dVWCS/zcGMrKI5YRCebG6XiW2R9YPGjcM9S4iJZ9bjICqTAhR+T
41xUUVOzPTcsgWzULe6SREuSuar1T4zcamiBQDLmsC/wafMAO7joc+hQIbFO4KXNNqxj+J0zMoKM
oxcOvH/CnG/as46QmfQMIp/x8U6VhJWuF9bryc7s7Q/nDapHBo1dn6XavlPh3nseBPgHeT9QljgZ
Yo4WBUTSq+NJaM3CCxbfqQzHkmvzGrU9KjAUA+TsNIThOG0+j/0x04CyXtd+LhlFeteFBJZljgkD
7u1gV73n1ByK0Im+nAwQsgUdf57xPrGgqOccIT++8529/sqwuqIhjDqtiUeiz4MwI0+TzpQlasWB
0uPtdGHbmF41vxqQuK9XOFsM1Fk/lCJ650xzQUv+HM+ebaGDpQ7fr0X4k6UGa4Dur1EWkZ8Cfodw
Cti1OEHlZSsjFkLuLcJhWHBzFuJueVxuttKDK9x/UkG6QxRyfo7LA3Ad+mYGiXTpPaKaqsgw0hSo
jaOx3NvCO9NZ9KBiPcVocA2bZoE8yufMe8kq0SQNo7uBdZixZjV2nH+W85BEg15U/Ww1jbfefdqS
yXmmhB8M2GEYBEvC7LBFUgd45KxMQr/lLt/G5VBKREcsnq+ThQJnbMDuEG2HBYaxztbHINE4S45e
ExztZuQRITFmD9+90wXgR+iAH6TnhHHNHYj24woAPp7hIkH2Dp3Q/k6DjrpKeiuDi4qdaKVjoWUX
Qp6XfU/1K7VlXyO8HoP56up+8x8BI+qgk2vuB5O7YMsO9ul6ujaweWILkzXWWn3EbyGBtWVWXSVk
a0s0rk/uK0fR9p8rEWuQg/NRn1WMCKTTc5aHylFp7269lr15Hc1fVjqjtBD/oLqIT5VY/LwqrAbr
2wBWASW5ySVAU2a3rRmL3WbKU7IwLcC+Uj0r1/xw50ZCTBH6UfoywOm9QgRj8rCgIkgNAYf4MRKa
tSxcWo4bM9DQ1m3srWjVXuOnQ/PGriN3vr4q+Jmc6fXbM2MefkGurlbVcqik7dFqFUS1V7S3jkkL
qZYGDETCgRMwFizjmMmzWPuYemG6oOQQZlpKyCzmRykDWhWtUL07uTpWELyq46N+MCCn7MkobFaN
FLTnSl1WE2zGM6vCWpdFsYMnZ08LgSs09i8oJllRCwSJOkCbyxWQeaGo8ackVjXfvdJ8+4HNfDLz
T5/QBQlYIBDySNMQbab6cX7hxIHlsABPwGWSg8Zn1uP7LMuF4i2u/hvts/bwwYSSWen9eld9Lf2z
6JkA9TzuRkO4AUs/aXDtz038S7t48XKi6A5NvB8cXH5Reuo48QA26ZOeWOHRoQToDncWEDH63kXp
3BHpZ2eLZM3RiH+/FNJJlvZLJaiteeqF11NMkRA64oYNf2DQHuMnzCHy7A8nEVO/LIlj85+97wnf
zfNkaRh4qj33KQqSLbR4QCvE5l5FvXX5AhDeBQdQRFxr8HosufJeUSYYNtnyzaOL+qWgzjCkgbHv
VNR8jJWD2e5p2wUzL9b5Lig5G/uJP53kV/q0t8FyBVox4/NgN8438KfS2BvTfnkZIzOZjSBtgXmc
FH5B11+znVBu88rfu9u03DoWnRW+qfhSEmAX0xl1Mtbd4cgnGjiAGXNdyxW1O10JtqYOUCZLgW2F
MJOT0SA9h2ZcRtrB5E6MqLt+cXnQOPLSNCgc7yqS4vPNrOMN6QZcg9E4LuJla50cgUFdL+EGYgoe
i1U6KZ75k2Gy1KB6pIqb4ndQuYKBareyTB5m3FFiIqIr91MOISCxJjFD5lUoT4Wr5wDp1Mp7RaHw
S8SEevn0P4hDgWKIpXVQHuw3Ya7eQgTYZHVlG+lSczV0HsBhxQOUpfFuDLVocq/vcMxCZj16vdNL
CiZurfbhblqJY3qECa+Fu65RJG5gzgZ++wVRNfS3wEAUZ9LO0bm5MoeXVn83vkDJ5DKl1fKGOSAp
l2HQB6e+BPEuGaEfnOFMyPnjGYal8TW5C2spgPdpTL/SaegmD18QYTsN2vVuFcKSLXb4nxx4+nXA
FZhxpXKmwXg695Of5J3Cat7WADveNI+3UMHsrkbLX2bBpfuDXViszK+NZkNNJXlmajH/DI2Dqaqr
i4nT2kQgFh4beZ1OCcwb3PL1shaIyEoVeM/JRF488+wK2D8bCOpq0Z3it21jgu39FUf5moOHSVvx
HiPq197IQ9eHzoqB24rb6voL4zz1tl3lxr+dwWakM+8OquNWGtDGldXYA3Jlbwc6bemWghNhe1d9
zO43f7F6IsSWrkIVi96/NpcC2VRud5Lvm/CFz+/Lt7OAK7pcTp82tjmBw+gD/D7l53ZujgnDpjNu
vyP6AfCeIR1eY7sMtZ07l50BSR9MXFQQgiTCXGdF658CpIVQ7n4Ns1yfjOIwII3iGOaeYSqlEUBU
ei1Jxq9s6divQ5X3982dFdDw6tq75h/usVFX1EcAZbnvXbV6eM3w10shO3bd4zPu98p+okrKIhfc
SAKU15dnLIAxn7knwmm4panSELclONQ+V0Oo0KnrmvuHzQd7WBIYi6dJimeB8FnltHGH3sPSiTxG
PL5CIx7MQXgd+tdBgIewRXqt97t9Sj1CqcpPQVtJuPPY2d+qxYcffTPHXrjgbW8oY3N5Amuhethl
co+mXmhd2C9oxjFpjJOh6L6HQsPQLGNXbfZEhYCSCzNuUwnXYNmjf0Fk+HQpb121+ymQde40gnba
tPp/ajIIkah0h5ip3QA+1GbkNEWfAqcrYXhws1LhocrNZ7uExHn6BwIaNJeiJJXH+5acnG84872T
/EaAphJUYwsTYMQmFegQeHUYaIrHZmm1khzjREYbUnJJjyVvMW69ba0mPWhfhbel/Un/QtmAdkMU
egdVCg//QmZ3VKdfMa3qawD6MMLus6zjP2MCe4mt6RriL5HKWVQRYh0CMbhky6/AWLdtOBB8Ipd/
bl8xQ5ka86KswHQEbutWhpGgEuM5Om8LK3HV0c511mGo+UNtzM/tyX1yqKm/bqw7BY8AKpr3lyM8
nIrPN/sUYJILBRE9HTQe3yE/eScsEA7/Tk64qlJeV+/tZwthtSiJShmR42nz8kuM+ogYp3hNVHIh
iX7gjxVFheUyEgNLKq3mNyx/ANPqHyl2fsnRec0cQ1VcrsnWn4uHuxEryJMzSRGnTaV8adL8PCTS
YRABadHNtdzS3nZLlCaOZoDX9d2qGL0k7op4LP6kjYB3hJqPFiD+TIpBmTgYGmB4gGQ6vR3oIOZV
6GSidcitUIDP3hB+9MANVgHhhm+faSTccRfNNtO5ThFjjdE8eY35lyQF7BKSpFqVanqHZnue6mZ3
ojfl+rGEFZAdn+b8uC27YAvGICBUn5xgZyHZ95rBFCCnDRH/ATRXgnFutOWVGTgxw1f4PJWE97xH
NDM4r/Ys9hwqzYGj4Lbhkq1r3ciqnEfwBjsBwPZDrNKMfZsxtbF6Z7RdgqTITDemM3X3I/eiItl9
z0DYE//gcP571oz7aAf+4d1sy7fpakvV7mgRvu766i/BrhsnxCjJeBqMwNx+TskDFUQEfiPEUV6r
nlaAJCTVDrbeCSJYSaikI8L8tKhSSVlA+rnvzGkkLdKN3i6d/1zzkTzFORsj5zRqDKoEjNMS+FdY
BVrPY+UTmSLnazCAolRmXTJe77UKBJxwZfdvlayv/76zWU6OpUdwxIiRfAwvtgrbTOw0cVNPuT6L
A9ymHMhuBFb0S6PgaQGzeZUwuTw10FbL36jUp64bMVvY8Sj7gm+Q03tGf+Kz1uh6vd6Ss2Pxj28h
5n755s15WqoPjhuxWvXTFpSWIrl2XXV9jlGrzjtEvI0ZOeN/L18Wm1CVvrSoOHD7BdIb95dbAwTq
WonvPyfU2Y6LP9r4/8nTmk3ymChTbeTYt5KQUmNqGJ8A478IeP4fB4V+YpGhUCbV2blBbqXDeVg9
8XNlpbm/6ht2vyPTQVjJXeG8PSpYG2QQL7GVlNCzWgcWDmfUuMALCFJm45O3x7vajpYWAIW348sv
lL14POroQ+cZh0ZjDhBe7KZU01McFWmlneE4XRJFPszImRWCqaagr97fntqnt5zBciCYvadNOsGQ
9/OCmhzb64h8vzu7MveZQ8w64r8DTvGXd1nLlZM7IGlYbMNhX8W99psvn3ilVl/fQI84bK49SxxB
FJUJNrJNQXzhD8jtuT6geJMWo5LRcyZIYpgaqB9GvLcWxINkGyn0gQ15TBMU3NRKI8PV51yx1Xwd
maEdLPBN/HI44UrJEq698U3+KOQ4blzLSBopImIiwVmG7MiNzgqUfwGOZq44haQRocW4zw1aGsqR
gutBggz4PILl9DZ4p/sq04yhS3qlBc7mGTmvQwEz28V4fgDRjOaGEqYtID99vVuDphvJruzpZfJi
k1OdoD2pRpL0u4vizRJMdZPWdUqkycgofjVMllrWlWq4fFIxpecetRrrUjbVPEw6b+WTrZ+t9A7D
edKVaP2PtaAecnQ03XVRxVopvi7QJrkcuu0gSXLqKO90fiHdMGepq1JgC/ep9JRgQztxYHM/sg5x
8wb1R75VkFc/Sl/ae78HhB8qJQGF+i2JNVSB5GFVSV6ArdPjHXHX9p+wfzCvAuxKbRnFHhOplfI9
1LSoj3n10qYAFq1asQjoAadWWHXncpkgB/fXyTcVFg2bhOaYkRfMZLUYCTfLAx5oF3DH42XSziz4
H7HbH2Arc8E0YDeZJdoom6rmfoN+JV1rItWzum4S2JzYhXWTFPtN3IcwKH2vb2R+6JoaHGe2hCRz
vU92+pocCHEvr5wgDa0iR+2yh0dTZgdb6jd+5I8OuZOcjjUsAvOFmcgFU/TiUVUKHTbyHW2hmVki
INf4Otje0VwLAwH/SW1LxndPZESAuHOyc+Y85BTQGgd7kc6FAmMpJc6OOs0I2wDgDbxo/hj8HJng
iNnnPyLcl9yRv280ccWX4fubVYcib82p4U9kxb/EEefKaAql6OIPpXhaLyLE4eHU56j2ZIxTmpxm
60+pxK2Dt1vI00ipNw/YubVzpQCbNOqT2wEjFdm0CjfND5PAeJPA9Xc+KHYkGUk/jZ4qR6ouwQjb
PTyRK20lkJq1T6JrLxMxGiVwGY5nXRKKk2hwb5cHh3Sr+M7skTJbzKv+pB169/dUaAN1R9cuWpOZ
J5jHp/UWoScJnt2E8uR7N1ii7uM1OU3/URZdI26P++gt0qGAvKxukTy7Mh5tlPG2V3PPVa4hLELk
iAH+cU5C3NFhjAmtroCUnZTzjUpE69MubJhDoi5A7qY6mhtwJgn98dOIvBWLAodhPzyLwn424PVZ
yp3tIalBDhgrYqOGpFrJIwUI1Fza5nnfcjOhV/mZ+82e2+FXVHtoZFMc+dfK8yvcL21pDVeBFFdm
HYhbZpBVT30CehVZ4n+KQcx1cANLYzYEpSMMH+HefwLeEewTMC5cWqpaUQ2Y719r0l43BFxRuh0C
E6tf49xzJHF6s4ItepMUwq68DkwwE/wf+SUCvFgxURFfguynj5K7LWAJIzcQ2v4bw6H4wlgHrnff
vU+/ofmaNMb3Wnh4aFA7RXhY1eMfzkNy10NnX5vwRFq/TSGQEmqgnXZYnwLJiCo1bmWdm2NWeRWJ
H6FHUmPI6zTTbLGwcj5mgDuYvy2jdeeb9b1QKrUackc9F3KNr303g1kOdZMXyek8jZldXz3VQkJW
2vHJuKdtmLtuxoOGHNY/nS5NcrIV6yqYCsP0hAUiZJbKLtvy0qodd8Yi5VXc6i6DFQCrTaarmC82
pzLZ2rCt18QMtFBA0oUcvLBmU7lOE+zTTsxe/+2bVQsh267sV/hkHLtyZXylYy0xotU1eJIiRCMm
xfAhucVxMraUrVc/OHwdAPNNq+FXGvtau/0VjMNFetEClZe7mGmliV/Mexh+lkLjuC8vSJZbD923
fiRMOF5HlC+n8ywm/jLkWM5VH2LF0/zU5fUWuRez4/SuhBq1ImSt3ybsKS1wc3g+iFZzp0G0J7+K
oEK4tvBjAYlQJgm8DRYO2yhwfzBAiV14Zh02K9a6PzL/MPPKuLShndiyIJs4XII7Kw+lAtaJyOIB
tsHO74PCHjYFuSO/fg4L1EXQfToeHGjCsvXpA5Pl1Zyul22v6OVe0lxxQrtgv5hkTUanDcY6ZTnE
HnaQG0QbSTbFx3FrVhkVfLfXlax7Fh84sR10bRyarCMBkX79JnFG+m4eqdEkaBXev16tIqB+i74t
Uivpb5mcj07d87ab0XkE1F5AAdp5gdgzm3UoTUH7QD85qSMwAel+onn2E/56RdA4PQXVItz7YsSR
qiBq2/4sjhpH4KjVyO7koyBa1zK5OkJZxOC9GG1qI0x0/wO43s/VeZ9rtZmiate+A+jNRgG+Nv8G
LvHb4LJU1rWfUSdz4ir+y5BQzjLvmC0I9/nKyL5bYMRB2rKZs6mzzlsLR7ZB8ay2diCLAivY9YlO
znDqk9WvHh3Zhy5ERX3WuD59hZukFmPupBKo/Y4raiVK5rXGawT16uR7lq+EiGQw6YZbnsFjAXDp
3rBetmmukjtYlfjXL2NGuPm9Y/JsmrUMBs2krrUvKlrHZiox6VpWa6Z8YjpSunkoIG4lhfEzDwrn
KCyR7DqYiksOk9L18T1YM/fMgOhCzE+TzcpTTEwSqjoVI+YK2lCT+YbVubV2b9kiPHPFfyWVQ1IS
K+t1a7vKMCKmFDv58q5Q16ZOiqRcwRQN/Ss9EDcy+ojTBhzSbxdNJmA8GJepc7TutoJ5DyvEBpjV
ePbOHNIbJ/3TExvOsNvTd+rFG5gaxHNzz53tzME9QikeN9+UMUGRMiN25R094geP3zdgphdMkKGX
j7mSlU3F/0xUcuQo0jxy4CTXvdXJNhq/yWr5Wo2LeF2klDxktXiPNSzMS+wyaXT5n49p7daoCE0X
4RF0WFG9EjdCiybic8dJTW/+K9abVRxdsuNLsCfm2A8oTDkUwy+lrC5ELeSmzSLd8v/z1yipGNMa
cTzYYt8W0T18UZJnn9eeI9yQBMVVqMMu4abtoYW7LsIrYBUHVQGRNKCSnLakQljgi1JqrJyGzv8k
BzyWbLemeL38tN3owDWGMM3xmtru6jtABvdYJ/9yrB8la7GaaRGCUHJjbWcw1rL4WKArVy87Oub7
6yxURG/viXu8CwiLR9H3oOHwEgCwi9LTF0Vs7NZN0RcatNk17fH9BvMwdQL+L6yiW1ypuEewokI7
pNsv4erjR8oy0wuM4HVsAcujyi6UqVmATRtykUZQ0neGhcD7JrXcQOWsPeWyMiuyab0krbF/2MKa
9wixisweLNk0SWgsTsaUloJPZdNgklElPvBBXb0mWIaJqYnD8o3FDID28c3V7Qau0Fzj0i9x40oj
AsugLbse2vei1hQjIl0vHMTW09MLbzvwEBd2v9EHqwWdJBiqtGNZ1Z4WR++izOWtbS6s81+COhoX
7tF59eHUnhfwV0aAzD1oUkxIan8F6gOwc+JW0CyBJ+ZE/oHKP7xmiTMYXcO/4UlsyU/43nlrmBk/
rJOi+5sSfbCzHKHsX1ol7DrcgRk24G4V9qktzqfk3BIC3jjSqKfElM5M0ZKBzGyETtoCXV+paKKQ
p0trQiMqWxO8P38nVDMNTLsUNEWizo3CJz9SoxQZ2rexwvY6hPSLi5XBLsf3gZGYLZULJsm4NI5Q
fvemgv+GTt0FYdq8n/e6jcfsdntPZ3LUePWb8cZL0OSX4nxEBmR4X/KcFRKo30pyCxXgF3fdfuMw
OROCOQwiKwIdBqcfMfQA0w56YoQUWNR1q2cBU6019vYFJehOvwReaXFpEyB7sP4QLRd+ldr0OXH5
J86jBzcrABNIOuOjpTK/Wcn4rI8hdo+SVtudrZAkaqSDZ0VHynEHmkapUxSGt+xNaaYBxHkbs+yP
292hH2ALOWGZ53aaBmJykrmvQBQS4iWZzWYRP4gz2/kJ3o2x46sz65/4mjV+JIBufAQDWkn3HNAQ
8bki/LKXZZJMkdrjfEtZDAPhBNKjhMlMs8Dk2lseuZpnuRxVV1sr501KpFguJniYxrHALDlyBWs4
LHt5oGSI+49ua09ElbAHb6hRpnQhVZa9m7Os2H3KG+2aqNfo35HNYaowecyyo6ZF8zsE703HGvu+
rc6+Uio8PuVgexh9JLp+xGgcCRUh6s+R5VHJSv6zFf3ld5OHBKALrRoquhdit5dmH5FhE4/pyjwL
UJM9jdam6LfcldKae3KWH6D8fvrMu30gbvdt4OwnCWKbiYbFwemQUPn6ljkDMxoNSdfb+Z1BvmHd
UhZmtYrIrUjfej55tnch3gbseaEZ52wfPwuEOpYZ7Drk0yhJtmLcKaShgilgSFKP25hl0RDi3NTU
VBEX+saT29j5DgMis/rApcL/W8/qC4JF0axm2Sr7u3cuKHSFbnkQid+epa3LVQcJFPkTn/BqyUxW
VEQjQjflaiy04bDGfi+ubm+iUnrGw5ETRLPBCrDBFZ1NLTXYWCbqRS0aIM0O3iHxQomg+6tdmneK
GL0YkYyeERmbWHwFoXLapGoEt+2to05ql1Lwl5SElp0sW1hL63nGrpy4Ml44gDOA7OoBClCWHK+v
qgC3r5WpjxypkeShXZaXeQC/Jbkgqxs2mCdKJxxC02Lo5MDDfJ0LXY9qNVq8cpEBXAe5IDWzje5Y
0E2AUq2+8uePgSJ1t2F/qi37lzz+jU4TMH9kRgKi2uQDL/DubupwIwHiXFuSSM7iyaGtPHSrjXdG
sHGf6LteAv/v20GFHUs8lEQye8KVjji9WulvuGZJgNnxSA/H4yTnpzBWjV4HTgFNRGt92NsBvA/+
B76B1eAKNzmnJNu4o+EQCnDJ3qC4vZvIqFwwSvQA0stbK6rWVOtzPDsR4vFgCGtbIf/gpzVCIhju
HOf0+7rGPnLegeDadVnA10c5fgv6TwmmzR8yOonf6zZEBk+HsVb0ilgqY/OeOju2NPceV7kQoJPT
JecNcyQpns+vVOVDSC2lGJ1mfnJanOfFc3ZYPC1RKN+K0sNsjfSUvlqE/CDIF7mjVsXyG24md028
OiLkest3b0AvrmTY11QwljAT7FJJGEldPmCdzGPwlLxZCm3SlgEZZULu3UWZZp4qOQbNDi2YQ61R
THSvsRWPgPls+D53PnJntRqVDGrUM5orR4FzqedBPe3dp8E80g2qXDppzp9oNYsRbSyAcNSEREFU
SugAq1F5GtrC6q85IOki1UHAGlSHW1QeQ0kgCHLdAjTVinV6Vzj52HVKku5H5rXsXOk4bk8WSai0
iR5/BQ7OMXfkq4zLi0y/oNtVw02mZfbYMA5eGEkHtwchgopnHRa6fN0oBqqm8KACuZZFUjYiwWRe
zSxwGdwKhffdWwhiRmzKEJJJbFyD+L9nkexwBJXnmVZXmTabNz8UtelN3ZgpwIe3aS/iW2e70WXS
GUXLD71oyhJABu1p8XsPE0aPfik4YHxOxMxsZac2xWRJiBOrXKVOz/06uXOuq0PpQofQP9st7nzw
rKOFkvDgahBNM6r1Gu/3w6eE4j5YrBqFIFfFow+etDUr2FR80RcgqiCaM8cGtEjrwYMIQFYctb6O
vEAFinTB+T8P0z0ajPR8XJdI6W2NTQJ5V/deAp9C5GjjvpPueDEyUi+VcSYzBWbODn0qM2Npv7Lq
9oq6fb4g7NDHv2YfAY+ZRA24vDfKsep54ZJlkbdu/0o5VOaAfv720Lf7t7aiEFyjjd137ZDGdI5d
ZYwXXC802GX91eduB7AANlelMrRQbQDZP5VIijx+ehC24/eDzcK0UibesoxItdgHVOhznsc2TLSx
szTXq5ERgQGnsg7MRZLe2AMDbj7oM9hHDfYQPrGuIFHXuRIxl8ncJEQn/uCks1/ZyYFqrEAn7q1j
k2vxBkamEu5DJdUUKYghGSjQCGy4O5/IBG3Kdtwvtc57VhppBNWvWq3pwZLiUy2YPq4mv1bUSBvb
3LtE+ztuBYDsmp4lUA5DxeCXIm7FkL93BnDQrft/rYBXkmgDTl+zHsUpX/JCliWYWjnn6q6SV+U7
4IA55qixvDy7ri5j2DloRb+Y6Mas8xxwYfDOkIsozVLfvRjFmLgi3Ih9XvJHYWEmAdOorvbnckBR
OKwDpeBwY9+LIXgWP5kcTnWCAOppHiiHamoZpTs0OaraF3mkHmV/vGjoKxslpK/+INRVJuzsXyyU
5u8v8Ql++nCjxEUVWMqu4Hjg1CJ88r8i3nIpX4+Olear52kDm6cEI0pKZJsDf9tqrwBmJZ0Br5YE
ijalT9brcUfLSU37JSjot3bmtTyY+M8vUh9mtITagGFFWvPlxa9dhHBA5RIkEv90h6bYXYPi4iJ3
gcvDA3aFi/+bLKKYnRrLZJNlw2HFOfeMAKoHTD37pb8ui48H3fyZumUFsenNXvgwqp0N1TgP09X/
A726rEr8gWAFxwOURgCrN4QjjI/oWOGVyemGAtY6tEX6Q8RWCP+P1DpN0b7JQCr2LIQ/BKICXaq/
+OCGopFJQ9p2HFMRlVagek6Roj3+TjaMHD2vdY3BJpRZ6SVShc8tYeXvivMC/KnBfEX6sHCdL0jB
3JjqpRWH1XolD27LNUuUj4gsp5FXaEiHQX3l2CgbICOZUktKW+r9Nppzt4eTzQmf8aY01fS7JFkN
4sDJUaMa71MqwqGMvdNZ5ajnKLthVQ4QpbXtCRr82LQBErRzcVu1YwZYy7gJsyBRw52B0FnmwE7J
lGxQuhTHB6ez7emGgeILesh5jzMfGYNQ2CTCsAnJgPxjRbchHrTK+ayU7kCzCJV/E8EZ7/bPJR10
016dcg3+eIxHN5GSYatX42fHlppV5oWJjLs6DweRvtQB/l0aTAnp7717UJaSRWyccCKl4x/RUkYL
ctFGOGwln2gpqFL8HAHPOqtzYtOexF8crB1hKd9rSoVtlJMy7g6CnoHtxs3uIBno3qLLUA4kF3Ro
V/Zda9pHewzax7qHl7aG/ghe5plvPihQs5nRvWewiwudRBmBN0Sh7c0lD27Knc9RKf5c0FJT3hOw
ngSyEaqhujE+Yp7QHDp11ZVywmiNH79Je9hq14U/OBHJVsgnuHY7euuTHjXylu4MoBtbsCe+nQ/A
G2Hg78F/byfPid/cV5JNh//nbohgNWCLDPv6Of1L9q4ocM03freCI9RFowzF+Xf9rxfcF258+E0L
dqhmSVmPunhIgMwv+gehFqXTqdnIKUJf5ZuDCAnmFroAD93fa0yRtilHIfkebk9mMDeZJG43mZyW
aevp73t7lmQe5Zvot00Jk3gXwFOPi4yHGvmhZKAe8gouRFdhg0HgRNT4aGnxIDF1jadIbudVsFOj
wyCG0HySG/iu5pAhVqen7GWEFwYgNRKR3vQSy9gCj50WIy4l6OTkHfLiJ2ARgIfp0BvI8a9eS9ls
UyCpuBmzVzAQw++E0sXDnOEQtI00cWjKGPGkrBPHnSs0CV1aN4u709TjqecrmUeNsK3+0ZFVVqNR
QDid7C0/0p+9TaMSBVUd/yWiyWHuigzD8Y6hooNxJhkCHXAlxD8e6VLniH7jM6r3VYfbmdtkNK4v
YW+Yp8KcLSHtEzL0r6WGrm/7L5W4kD9e+yC5OuY1lpdmycFGg5PURL9u57MsdcEWSq3NQemwx+my
npKrUjBoPKq92EJQL18HUI6SX2AaLvDVmpnRlHjjl+jaASxrbVbIkgIqZpxA7NYaBAUhz39xqXdc
yJkTpvz2Mj0DuZStYn5UCnF7wE2D5uyGNdfcuwYDL4V2y2j9Vgc0QkJ74Cvx5pKNTzWCzrDbGEhU
bkqNfYc2Er9+/AQZiSocnRkPNkLphj8lJLDGQtQ9SHoW9WCwCrpeOaQM6WVjFm3eOQe3DVK194zO
Q9BGkVNTnEtvOtIEZCvCbhfZSbsAzHB73ODVBXOyMv76osaAtmdZxa73h3D+o7WtW90TBaS5hqSi
Xio5O1//2tJ80NDZt7niNm2jLz4vcyUu+iHyshSoDxrJl7bv5rjq2sskSwaT6cosxi3MneRGh/uh
V2UzXZUh6XfyK+BYn7izeyXXfcycDjxoVoP1nN22z8JA5CVJOKbzU9uhuxqRgSOzkH34H+TfDPQ2
/MnM1guk29co4QviAEnPlOgFLHUiB0BMP+j4lO95WL1A73Cd4tNZWl+6gxMmwJishSamiePhQQz7
WaZXF7mmSkuUxD3b3I2nTrhhR1GaS0P7x/Uy+aerPGogRaLcZZnupcLaRHOUReNTBj/8fC3D+8y8
rWZEkKEoqEFO1vNSE/IOUlCvnHkFcbeUsP1Pigwx7n11cJ+3x0GE7YxiI4M7ByBsJF5NlJYHXTzP
oraQVFNAdTQxKx10kQ5sEQAEu/Xaw6wlMCfhLTbEx3AxQwyhgx3I04HNdbY47USG/fms9VfDonIC
Vx2Woi+LPnWwJ56lz17ejxiwctwxIrZAL8N1g9HwXW9MUPbLivNIsT6fMiyGZhcNZSqTgVW0LAbQ
ADEL9SCJdXVZOHaSinE5OoIDMptCcEjRZOZ4+ZzW3ClZAXXeXwY8Mnj32Pf4eI1jpS6dV32eqBvk
azjxPexr0ub86T7Jj5+TlsCrdUji0sf4qvfp15Mghdj0CPAi6y/+d+IuTdGFqs49lb84OOQs14q8
8s769oJoBcjXvssxMV1m2s+X52SixXgjey/iHhwD/boWgYwm5zObddS53trSpHPt1VBROW4fsIsj
nuGctdV07aZ/SnawackhugjJL5fDGEVd0AHwPXWhKsZoO2YlhEkTfcmKTNyzXk4zY/hdnn2AbaHk
eAx4Ujtep8Q6PlyvysPKPkR73y1ROQHG1nHb6rA58K4RP1cMOcto2vRbvCb7PPdkH6xe1tnPWp9O
MQcTZLfreDmgWNOFz0nnNlar4kqKWvoiW16Sbwnm1MzSLtOFKI9l6CXG/gV8TSp6vxU3b7bbKqrR
QzfHdC4oAWROreXMNHBjRu4zWEZwkNBQqBxDDGIli/FuQKUkmK31dB5KdDXPO2YTexJzC6q/FdBb
dmakK6zI/qXgaIKk7gkWyZEh7TUXdgUlClDObiptNV3UBC0PkF02YPMcLasFbPuICn7IYo9phWz6
LMfuvwDmk5GiGX/QeeQ9uyKSQPTQEYWzueyieQcXlaBmz9gy5sAXHNuxz7IZ4/zkQcb8p6ZE2cg7
dttzZtylZRj2N/4PxRgz68JFkY+mDFfphy4BPNCh6BFPcnxBPyZoxfEpwbfMg763c4pH11OH0a3f
29Jcb/ZVhdMxG7LCpzOMoRHyPXyeXXNwz8yPEbarztw5EdEWFx/h/a5d7btxjUiotSQUDv3t5zXb
h0qsi3FKG2hAakEX7tTsKaJqLUJR8cnr5gyICowsESRg80qgJo5o9B1097r7j5YgrzZtB0foCfXy
yA6r2dTiiln2ZJ6jD72hzj+LcKZRE9yuaaBpriGWYCVzh7JtMWGgUbn0A28Hs44FEqNNskoWiVXO
oFaiyswGObySrGJG3P/JNW8kXKScYk7AInXICZZZdI+L0Y5knYVWoGu2tfAUgOLJYLiuOz5m2WcP
ayQEEuarL9ykCiFBNhGXXMUBfD6DF+fRV0uutqKuYVFnLRAIEZog/n7pBcZd/tl+Q0KgNUtf07rY
3C5YYac134UN8iux62jKurHlGJBTN9tTKdtty8DzuNBe/Bk9wDWkbVPy/IEU0E05i0qT7r/oNy6K
8zB5T6kCPaH58rBguKeHt0MoZpT7pd8v3/flMWEbQhE4GAzBZCuYcNko8cqyoERoKjlT53k8r3dC
IlHD9ini6Yvz/h7ctBxoTZYQtwa3XkOJfonvqnpzmfm4MYWl5BCK86N7WyffoyMBXPRooQX/OEZ8
BkFTzNG8n7P2PL1IfSrI9/H2B7BpGwKK+oI/2WHrtH2J7khRHyy1j/pdJfepsOAn+J0YzZTXVnAD
zyjlR92vuaDukcNPUM3TxJ61VcAt1VvR/qyWsx4a0610aMMCgn5OyAYYQ4YVm8FirzSsjVdbNFW0
oEfZ8rnEOQmvJdqkJ7vN11dpT8GTXvoA6GnS9TBJ5dPctSPzxdBwG674n6XWeuKhlWJ+00nOzL7n
wV+WN440BSRXS7atPPd/3EQ8AePLmGySILOM2ow93dE+TjJ7Nrcf+/E7VMhIXBXRbPnziO9BmjtZ
bXg25Nh0PCZOztU4Q5mQ5F6tOG4QCTZNRbQO5ZchkH2tS8cVPS4q8r1sdgenwTBPDymAoqtuj8Co
Sj3BJFZZWVaf1YPbYSqbC2zx4xL45XhWkk4dlI3w5zEFxWeOeWGiwNsbwfNc7HaHE+ShTn+XeDDQ
X6oWm+EFS1/nz+9yn7gigqs3fOwuYXKg81NDjccPaEayFXdkP+Yxrez4eteF3A1kgV7mjnt+aqy8
jRTiBpYid+m9gAWdWBfAzEBYoL/8huHlvJytoG1TollUEqdsE951sLbHZEKHRCaOJphxkyarGjM/
UMvVKNgfXVukf+7gkIey0kinGku+LJ7eFdjVo2u/nl1/QGvfI4+ww/udjJneoY7NhcTczpbk0f5T
vCpMwGVu759RuRDdFMMCBcBktqklWWUw5M+LCSHLk/G9eYztR8x3aHOCOcAwpiIqKPnzMIX2EehW
AUF0md8C9aXdh3M5bZOoU8SqgNq6xa9YePswD66Lb3TQYPwYrCdIQyG/J4lxKmeHdvODWHsjHaH6
uFvUFOrFA2qTxT4p78F0VMIZYNirz4QrVDSGcwk2m1wmudw42Uekt0i5WYJTxbSFIqJCt7FJQR+e
jdR43PUwjrcykqE+nsfjmJ77BMDuNEmh57UIa/WzQR/EFl/xwo2zUC1Pmag2N23vc6aOeKQbUr/j
3HRaeOnLgDzfLj2BbMwm+88WJ41YCD3v2sA56Uuxvwh8bTDjt5kWUMqSdOYQtzQqQKnCY8cRDmuv
rh2Kco2Yr0+Aia7QfJN1ItlZPU8BbbrACWMw+Ce7n33aXwXnV9A1mjNTmkq1oWhgKRVEsM/N/Hez
rzmyQ1nQuUKcLF1CZPolxJPWFZFJZOx1a7Kdp8/Ib8F9a6h0DtnAYSKsvhWD/mW+y19DAsK3M7wk
c4T7do9q+OQEDSHabGzTTXog1JTu6jfSkbzJMd3Rvd0Y+Pi4okXnbT91F3MVHcL/cJy43fnU3Bjj
V1kAXe57+ao5J4OOkhWW6M2ytk7sXaHAr1QW6vETYw0hG/zrbxHZWLw4Kf6nMVpqV4O3FJAjvh9m
a/YnoIphJOVgaJ4tx72EKFep2q5ZOm2/KDyP0nwyw04bWBzg3YhqRDFSPvCJLPEGqU9W4uXcpDL1
uIhwAl8QDl+29aUN4DS5IgisyYvABPgtJvwoHGpCS5BGdVGYt5ap5Lm7gBPCegnpWFUw96HD5v5/
77TS15kG0fFl+DmRw5Dl/MGnSfmt/Xmo11FRiXXsDKAXcjlaaQMzkF/7K3Qx7bJv+RJ23dzafPur
XJo2pmIELjzRfhfLVsjz9Mzv97tws02jdvhXFN4KPRVCNhsE7hMvi3eOUw9c6QEBfeUnLuwl9B89
C+8ybTkcmCVNteuO8y9Wv9ytJ+PgNUDkmwCO4BHCsq7Lios/TU3hQYJ0Js2tPLO+8Ekj44JFKufL
JSCQ9IxHwWpJO06xDXAMoT1i1v8X0RNPDF7QWBTBabGLU2VAXv4rCikZmE1WPLi0tFKBVBCwX3xb
bKdmPLyd8RuSvN/q7lJKeuL7BqmRwfUMyQL3i59kgT1lEVt7VlbxfoKoUrGPyb/w3x69MGSwdfOt
uNQ1hxHoFbRCGpSgxUAcivz02RRicwxdYJ3V+uboWLtTf1viL9pr4Mju9ij3SeMYHrJTL20sk6I/
n3yzVaeP4INitnvKVu3QjrVQ3//2xV/SdWwDQnmPdUqaW2rFDSG59pBmtLAjSLNyEPlAwv7ZkFH1
YVm2sykohwOUcWd0PH+9nsGMW61w5hQKU/k/IkPgu1K5BKUO1bQHtKh5UJOi9pMiEk6pwcPO4quL
A9sjcei0uUcOAj0+0Y38o5kWE8xpHe5DJa96OcoxzdVBZGoUjQNDWiSe8P+W78WIa5GKufVuNxgS
0M3+aTKVNA6Sh6IIW+a1rrmTNPdaKA6LhjStCjub44MQHDwUko2sKMSxHB5jsUjev9qlQSK3ISQR
vUKZP87EU4GGmr4txVa5ykI1EqeWN4k1lWaePFISM642J7YnMqYaYxT7vAX4Iq4mLOIJCb8jSXc0
9cL2LFqZcBzTDK2tNeHhiqsGzu7TTKZVZZGWmJD4purMJB1pZvDb3oZgEpuyxHcpwEwCZrgy5hQb
rr+HBm/Or5MTUILwnlyi20vumDwKDEpA9BYhBKNYlwhJ78fTHnQH9cahxoE68eJYjzLwXC6JpI/s
URRmYDHb8DYME9x3rNPHq7HUc42b+X9DiTatOGRfx/PKeQetkyD6yNiMLGS1z8m8+6d2ZTiFMyzV
1AKUOhEQVReB/uSyWD/N2mgBpNKycPE7PwzSqVUO/yHr8nXcKjar7QbUMsyp3Mwf4PzSYAFLzCWZ
uJQt8qqRo22FfyUimP5rRBuwlGKkPqhCnk1AlPmZyzmaa0lPuiW0c0ZNxRF8Xs8YU7Um/r+QUx1n
ydszwntZW0PAW5pfAGnsTnYQEFVGL7U/hmugwHXIALDinSZ5aACXazo1qsZhajATzZJYJkvD+Wha
j+8jDW+xcr6BHvDSGXJI/VNO25fKmjXIkDVGxFN8xnreRbenTYwCFickZp/8vXRBDjIchUEbHA6m
5occ+276bxLRkaJSS6bNJoqtuWVi8EPFCfVbbT8Ig2i7VgKfc/uy9DohsBSQVyFdeD2Q0s1B5Un9
8w8HUKIUClMxGyCaCl0saJxlxvGMaUnaN9FvzJRd97rR8IHhuQzKysRK6k+wVBlvXABLDJ9XTw1F
m4nGpj3o3qVlFdYcqsiFqfhF3GkshrG5utvZQtfT8sUmXzf1WFhtPulpep7TGocz4nZ88uS/gYuX
PqsPy66ZjZqDSZrfkYzTATDbe8FdNZkW9ya/MBdfT7eVZmgAn5AcAYoXHKsNI1sHWm3+bPiyx/wu
aBwG2bhiTddNbm0wLCFCxp6I5Dz6NZ8Qq4a7z41otl1VVjcRrJo/1iRdi5drTZ0gSzxBlC6Y1jdC
3lopAT3YkDQwF9GQEFkX4R5kmVjlD3BSp3lohpuJIFc//OfWDznndOiCpAEpc9GIhenAEfiSi+/i
tNbl0odg/GqQSKADqlS9yoR1cJfBPLmJL+lCx5AnwlCbJFplLY/y4aHhiGFht9UuMR6+WNdVs8zq
zcvzABuEM8KnKrGUmqohDi9SLAasZPFCfO9/BN3OZB1OnXS/dM/3d3VNnsINFH818UI2fuLfb+Cn
/ugPOfMmNLIYoccv771KNU5WfnEvBXzv8Km2v9xtPI6s6He8bkJzyLsrC5fPgFcIsgyYiv+ymW2I
0Vvn15lsU1l1r8bLsd8OXmzYo2xwPT8+DU2xuXAciSQqr4ZDPJxMW1MIPQ91ZhJScluB+AbSQt3h
ltZUHs7YdbmSvZTVDW9D4thoDj4QFyXjsHt2/Dd/RCvM3sMqffDP7dkAEA7ohPKae/4PVQUxLn7e
CqINSI34YdBAaqV5maBrndkpI4eedQ6A6eWd9g2zV54kR9LyrKgaXsxcFaBR8HzwfbEZqFTHurvk
1d5L9pK9GdW0oC6TUhafXoqdWTYMLhfvQ1daVEDHwNwfIaNR6VOxQRxgxqaNYgrxP46yMcYZLGG/
2jdhC2iS1u/3ZlKCST4r4dhPFz14tGqwZJU+denoBIvlpUWDRi5iX7zEvp7sT+XuY+VWsIg1LOqO
F7u97fmYFjjpI1Onh6FwFec4Qmef5La7ygPBuFQ37NqO8jcrjfUokiq/W0Tp/EImJMTUxYxTzb0T
SQDcKKlevmIXfT5Q93JZ9YiGULDcF5igMM9QJFigYltkn/4+D5weju3q6rkdXiZk/GpF4KwkF8ss
ozVFS22COo9yXAcRzbPlzNQAgp/woqTGwA60bPlxFmqxHPq+eHX0Pre6DqM/HgXyrciC+Pi1Upqt
gsz83mjHz4lm7+28WmoFSXMutXsLM/TiSVcDO9aoUBS1DdhzaxCpsQAK+D/Lc9EOTv1UG7/WycZx
x2Zfpnd8xH2JfzPWcRoebuTsGJrDtv0aiKuCOO8dxPfyN448GVgWBbORJ3Bv+qR+wIl8hUwHFZ2n
aaBf/VmzEHGW98h9FL6ZLbGzNB3QCSb12nbdxnPE3Hl7r2a4rYBtuT1Fitp7/wLujqtAchr6nmRJ
Pp1JO8fu/6PDaCcGmBwkp+cVQKT36vMyk6l5bEaL9zP3O7GI++A5DsoF0ap9jvPlyfsCyUBwEwj6
0u5zmnI+rzX2UWzrtdtBbzfVBzAd9JugHfkDFKvEDL08faE4oQpgdA+SsTb5OLTNGevqDzu1Ksck
c32soDopThJf5fDqdMFKQXXdgbRj27sGy+SSoU+UEuF7X6zQdx5znhmZECEpus2q/4/ReyQbvU9i
sFuDmnf9pTKqwHWJnxEPAGSM1xI0d+Bi4Fvq0o0OcQKe/GYULZseTs2lTRrUcNVo8FS67yN36z40
nXhulj9m5c9R08opk7WN/dpEK6K+GWi719RWpMuor/gHo71Rgqwovm0oJj3HyHxvWYm06HSk11lU
zWYIQPHx0eU9v/ItHWh18/PaAtEymZnCnZXBLkaOqdLZLdhJdDRFHNU4JX3sC2JuAq8nGjBtp26N
Ef6YAigPIWahyOSrRNRM/d8NiCvqo9grwipHqrs7TpkNyYQDalbRnPOcccM4YfmHE9eS3vl27Oh2
QnYzR3XDUelrLvjpKJu1+7L5DGDDMAgsjzEos9ZsbQk8K1dQO2wl6VjRFHTYAtJrTJLcwfZEFNXp
sXwlgAT5enWDRUUNXdAFXbFrfhv7Sq/jDMCzp3wO4R9ibWc+XfUVIpE4sRAAdDV2J/CVDeG2aQu4
g4VJ5FCOYlRzNQr3rCQeExl46oiA3Jhz/P9zOqAoBh52ie1a/6xW+pVT0ugll6fWdh3CJLUgdCOX
KBqs3gr2+9mJkSx1uA0Ay/W+EoIPAbQBDtlaEj+4//zcy+TTWa4MySSXdEyU+ywkDfmIJvD/o6ER
4MYYw3KIs+eMxN6u/ueR8c0LjDHZ4SjjtkyYzD0kq8l3EN2yMUsuqQjpRMzUSIeG4Y92E3E72evt
tX8IoYKt6Rc2oiWjgDlJA6kFLpvtG85quaS6NYdA2J0Ihy0P1tCGBVqXm1UC0hF/zTlwmKwp58gs
uLEJ33HpGg93RkHyf1mqkKGqvOGvxmzAYmyOf/v1MlDeMRJ4ijVm3lAJRP+ISzSrtr+sz+xw3ZDZ
sNNdNw7CLV1peOnrHMnKJISPHEXJ5RljlAjaLaB8oHa33wzFv8RX3aiqh6mS5tIac1JSLEALvRE8
BcLv9bZ43LXU27FZZ+Y1Plw3Lk/ZQYmeUcDXnQSD9Vv6ATkstxI2SboBtPFnT9fslq+y9TkViJAE
pbIljFoxy2HonbmTiCuxUgS5eVwENXigjVSZo8e8wMGaJ8TOYXJTWDNHt1o9eF0kK2UmMYOT3/wP
jAS+hIfrJN6wUYppk/I55b3lQt4r3Xv0qUdCJ6/kZolRH883RxGLaVtRF6KNA+R9wRmJhTWOSsXq
tlQOMYl/wN2jtM3cS0k8gUpLf1cOFPMrYncVMycYL50EBMA+5Jyxb1V2U4ybdGJ3X2i2cGY6vfRK
k8YW85Hegb3wG8dQkPgELMKrVnGfKHTifOjZMPu2vmN3VHUHa3OIEgfLTXBOyQ7wLLjNiVB77nxF
Z+iB5UXx0gZATbLEK2VFB0pyec5OCBCbut58tRbqKAzeX6xLipOH2tpHTK3+V0tIgB8dtzg67dbh
O8fkbjGrro4uXR/mgi9dVLuLgkgazvndRRRsZecVmPLZtpNpYfgSTRNGk+OyF/b0GXRWA4IPyxlc
W0qH1fQSZSWS6Gs3M+LyMNFeK1emS5bdZbYUGYvDnelVtTYhFjb98zNjDsNDHQFBsjjlWnNK7HIu
rvYGWjLYKnVgWZw7vnGWy2b5s9sQSB5P9mPpTu7BOLHDYxxGrlRwpbaRts6brtTWXx0Y45yg1rFG
Ht4fM3Q7tnKNA0BMHJkLiu+u/oUKao3HPOyYE7i7f8l63fbTjDwrqH8A9kaiF5V0qb3QL95r/lE7
yhW4XSyV3rB4hvul1ffGbwkkd7J1iFYbbfu2SBWy7YK/DMJDue7EV/W3EPfYe7FStHql5/Ts4vtZ
p9WZ5alEYh41aQkh9+o1sQIwd5poztMiAhfsL8UM4m4LkPF93TBS1rJGjjzkbHiMLuSzZ3+HTRiP
zoNU10fYpJmdFQWkzPCroipaGGGT4+Npbf2UxPNaKosQ2ZBstHvyu7yYOwOkKn0oBfyuXu8t6WUj
VAZ3BWKfqbRANLldNZjJmrUX3B2jdt6XsW1EUKfl6/1Gv7iejm/p/WjW/hSSwX8FCPOZXx5dBbka
oSX6TNEs0Y4lRRI9pVW/b3FD0nX3pcADmM0bxJ3Helo+2zhuxBa9DIcg01vPxZbz6dLS8XYGnIYk
I4e2IJLTFxX5EFhi6gDIK0X1Hf5t0xNdKq1MWOu92HsgZwSU2hkTMki6/hEGQu6SDKw/Lsh0ioha
0gfCFbSnCXkqp59IW69Cq/yAilox2BNXGYVS0U4PKL91K3o5NPGe6T77DzgciSnL+xfn3CDRhO4D
Q7bLwELC8HoLobCUYxOFcfm7NCj2Fz3caNT2NgNoHgBC3gWpVPTgDaZ6kc8pwUiB30P7rNo414ho
BfJdKXJulwAIea1O19pTfMdt0khCoVrtJkBik6nfGiVMTvv2CljgBJY9ZA69J2T5xsV9xY3EsO0+
htVn+0Pah1QJxAKYcNk9sxWSnrtGYJygW3E98JfkvWeQML3xOAfMijwHuE2uEC4WmsRK82p8T5lU
bHyV10lWFD7SZZR4KKUt2WeoVycFKzHnOVhGzrwKROEpQnoIkSJWxrAV3jhVOP5upOFaxV3TNRAJ
bAxSjgPR8XgN8jYYFPhvQpPDbqwJg86Bp82zhd/YTv+uD2Nyeqlx5KcPQvJKOJUjWg7bWJzX8ku4
LXDLD38a/u+4ElKJfP1HrOGHz+FZu5jAb6Ox8utyB1gf+qFUH1B7qMtmKAkYZOrreitZZYJC+nWb
Y7y7132TIj8L9zGYShfOhAjWB57MnXwlEVj0NhCoFUuHyV9dTvzycLRFLTaHeoV5R2DL+14LjGhH
3UQ3VJzqCi/rRUApFXayDji2TdtOytwUVwU264BHBZemgxlwK27Yqq1UZFt0no8jIHuYjlWv/zk7
im0TifuVDvCKhUSP+1kS/57MhcTOmejJ7TygUZVI3nNI0hzLEfktdI7jAG9andRF85MmQWFI47sn
5oy3boiy63TEuhbA1nwPPHzEKSlAgv4qhjahahVhJSY46sFX8/n7QiCxQFVNyEIbPB9KgviPCOOr
01YydesFc+i3DOHxgTsrOuOWP8Fj/p7dMY/m8HKguoKxWi5G4rTbWxF8z9mJh2jwkPkUTC38xb2Z
zFD5LujiHgGMZwOmhonecZ3CcOCcnXFux/TT1j0Aipf82cGTm7YNp1G0slmq9g2HTpA7QiqFeKpd
4E2AulgxMk17Z7Kx9+N7JSbyiATdhVC5CCXDe3hfq6FvYdCLvlhgjY/UDG6/Vc0yUKNuJqtyx9WA
gvSepwO3uzE3e+Wp2kBO9Lnk/uruBzoZT9auWlyLfkErAEbBs9Ejdb8UWTUxTsnCzwt013uRBcZ2
AT5uar2e4lmXHkrMBvf6iypnRjaAn+DBC93T/5SuB9JSgPuj1BcV72FezdKxC4QWkmm2IjvXf/np
sehjO4hG46ZgGv4izjJ7eppAGn16eD1fAkgiwKlPvFhbwKPmysqjkLHoTTYt1xxYjbhn/i8bN7O0
kel5+QDlTein+EIEQ2AQLexYj3kLNr7k+F008dAP+y+fatUEtQg4kOVcazXCB/74j5kYdRRLikaR
FQ7PEHgYdGGFCD1aJis0D6qeIDOgnbHbqN8z7r+mcsgalSO3xVgwPW8H94aN/BGPOvdF3AaZezAt
Bucw7WKP118dRhKGSu/6WTjD7EuD8SHrP7FILP1YOxceZvra9NcSbxXmT7Tc0/Powiz2lp7SMw0x
pg0S1yqXnfIb4wTT6+V31A+K705VnSdaMMK3P+xajrFEwoWMY6zrdkV3nAyblOOXIiRgnpXEkLkF
aOnSmaYifddyKb1KpTKsequLVBx5WkW90nd91Xd7aL36kd0xRQlOexzFH38omZ85Ay35200E94my
iHY3yQR9tGD+rgn7vxdFEaXxPdUIx0MdcFSNAJLiIPwinL5awuF/LJwmMbbuIQ4Fv2L4U7mUp4oW
LcOkfl4AhyM28CdAfTS/TgghhaMPDnJ1jeDhtMXrtohkGvdQXIwAcsxTHhUSOQgi95XkRxeu8AML
8siObmHXfUoe4d1GcnzZjY/MJRP+zVxWuRbC7g3zz42f6Ky2Kr6fIBl1MBXPHvO0TdKdy6N3lL3N
yQzUZpoVqQBZjyBTwHFaz7BweSPhxntkRa/lDxdoCtFpE77douRBSL81iVaPOK+tcBTSv2506Z1t
KHe4Kynsvp2MH2480u8n/KKRxrRAD4jEif1HoYSgqI8tz5m50jpfJQRg46USZxelUgwbp5X9wkWW
UobAuYmVCB5cJP5g9nPRYGTBjqt+vPq+NG5QpVa9a4SNl0eHyKBMhk3fxkrZkp+IZQOGcgwoA0Xb
/OkObGQob7rjI8mYbfJavYcsuc956TJz9j59cT9dRzKNBLdzzqPKwRtVJHrNRAFTIMUkz0vDcovZ
TDrV7kCXVxQE0xhJP1KrmurVLy3k1xk8h8hUb5CeucMmGduRXHDEhzi1UdCorvbivKshkcT8kxjS
eAayyY0gRw6yWOVSKp77tul2hTU6AXjrxRFHcmssIeggbnTWmlYY7tOHo/d4Pp0QtsD6SsngtD2X
e4MKc+hCZSaDj/1LvgXi1d72PkNWdQMZn0qFYNFaTPgvYHCKVocVkpA7fMZgWEtoDPXPEvjEPKeU
01DmfPvJvjxjo0kxKz+EOaQ4i0CDzjVcWieYtfhw2jaXQuFwd0yaqRRK4NrFIFZPHECi/udf+q36
LQuSp5/yHBVqrfYfkv6KpEotKDs+hsoSwzDGvziJq70wSQ4Hm2brF/M1sGSKRXFeQ8JPAZc/PXv9
L21w1u1E9kEYZCwWsJ8mb0QBfuofkApbXtofzssUQal5ENb+Q5BMliLVqfo8UEgpIs9bNMf2HgI/
p0rH3ndIXZabOb/r+cuMAJEr7XAyCSCkILbx/l9D/qZihcahxLBsHeH+VxW3tQGKYROvX43SiTAL
MeDnrEhh4CetPiUJwR+0f4F+sMlv8mKCBRu/MqjfOVg3h19nZd2nQWZdFvP3bw1w+M3ZKMgh9oZF
3yvtbBs7m691rbAd3yRCTqP3Z40fcHL32FCW37oGKScnZjfjY/w1iS24kmOD3Z0wGz87AWLFWEdy
Qo05FYJ7/C1LX8Io70pRWJ+/l1euxPVqk6xEg4gxihF0//yuRW2wTBsigVtaatQmvjIwLt9+7AVe
D8N7RsjV9mvT5R8zYqND7rD16Ckrwii11IoXzfBRXfS0ZqvAT51E9ISDLAK+6aYqDdoW/Fn9KT78
C5zbAsTEfaByzFYeNjJXo0zgsJ/j1sT9WzExJAmI3SMexGhNA9wdKGmtnRUkZ6FmVWS1LbgboKrd
w745ejQYkBmraY5u0w5YaO9crDdUrOMrWOl6RWc4lkbWYGxYpqtpBrRSLZ2JBa3iHHPTzum+0QSI
55TFZUBS3/V/4sZfs5rEIHZkadwh4UdPzo7SxVMocAuZ0Q5RdIcP5iR6GKYVE8r0LmsVBVMY8tIN
CzdTMbsjZJaNCg/kw5PBre2EZ7SVB+HyKffAAcNXv+tpXT55wY2EFVz6dARVuwy9CkLtR0dp8hKw
PyG5kbhP8xva//l31HBLjE9VbqIh9thAWy6Wqekk7WEpPEnkfjb623KDoCTypKm5YD5DTKtNK7wU
atgGLSnU5bb+b/MkH9fbfVm60FYQflrZyKZmlkXZFmky/cQp5S6yOfJfFKNvDrECfxk+jbBJfTyF
3cpVwHbRA+ujx8oTRsS3CYceuUNUYLLU8oO17pMNWdjeULn6jmGdq4IHbTJ4PdfTBIYTKcuZbLeV
Ps4WzHkfixHnjZ+aSBu2wnrktMrMNh3HRvzbHnk2evSmFHsoW+g7AMF8kUX9DLDRTN1magkJgsmc
jW1d//TzI6dJ/1gMvp+BWMZlIV3JfiAVoyG3yUWEWxydPV4KCsIQcCFLtNSJWxKK3jHVWnN8WOG3
7P2YtLL54q+bvUQBCMwN1VJiS34tCiGYpwXPVknloX4D2fxqzsXd7pCHCtp052pOhdJqmfvezsDN
GO5S+T/ZRWMlkgU5/6sly4SBw+LNKEcTMDR3X2Lox0lsdwdRnoyt5G+ckrU5En0flQcmaOEqeMWy
cot8GoXdVc7DIeTVv206DYzax8IS8PodWTjYZ1iOUXTVL/ahyva3jcQvDh20mSwA90RNAgaMmDdY
ySrlZL/0VZiQGzjrWIOiFky02dkjaCZD6+NbFnpyRYedMLP5zDfQ1+3/gjpGteI+KRIsum+GV7bA
EFuKeNTQqgnm+b4WLeUvWnZ2/0X1cK/SZRfDh7i0pQyZcSFtN5XoNzqwOtuxjr7gr731XqEuDWuL
ZQ4FSS/YYCQkyeB54rgeJ6WC3MA6v3+EFK2Y3qXo9iXZSLMakBCW/qo9t9wSi3qZF+wyF5+FJTWA
cQ9oNrRSpKzecbLYOsl/I2iqq2xeNeqrI0DblzBVFvI01KppiK9Gl+Em2/N6E6PFbKIHOBdm5r4L
IiJ/aNndPlJQOrW17H0I3bb9ucbqkvBl8OX+lKU0rlLd5HqgV+jWGazXFEOfMlmXk1CfYfeNcDTB
xc5SXVyrgCgw1AG1yqtktg366Ip869U7QMkRV0/aUDBr8GVVk7abSxurxqUU8It5AJZZlMSKdUSM
Z2tQmlbSdUB/YcLnj2iPrTjHQv3597DFu6P+UAY7DJBMMnA/OqkFgYrXzPw9ANPSRuVAWvCN9Ue5
sJj8+s6NKlnsqs9Mlwp0Wk15Q0qhhDfnzjSfLZ5fszU6bOFsMNNlpLGlLZqHAWx0tXRog2420OXf
B5jw5Ft5749R71YHNg2FWlct3Ho83YVEDziQViH5xTpCZwi9qHjj5r24DCGNLsTvHZTHoDh4RXRs
hZUIV+jgIsuzE1AdsLK0vMjIBAGHXocZ+PzuMvNe3/x2R2I/mjojITPjBr2bDvWDjKq1o90TT1DG
Q6CTBwCV36LcXvvrfarKKSqnbFD7uKdtu45WnGhsnNOihD1hlDUQLOohcd9wB8BB2BbB/qBPjkci
Cc9+YPs8OgdWSy3TX1y9pBI8/626G3Hc+XIUO92v3SReN4xJmYY3KMv/UAGiO61wEQ/+fwWxkyQO
5QQ4KL0+SUvqlFINzhxLSe9Uyuc0qjezob5kAC5Kyz5nI6f/2CUgim6F43BOoHg6iiKYAmDKMs1y
jn7ueAqX5hXHvhbj48Q+odyBeZXAIy6I0vSC3AIglOvG5FzX0sterTy09txPdD1rzfnA9aoqz5dY
PT7gBBKfDbeLEI2F6H4YFWU23C5RPOkVnI0hfDWfMPCRQJrws3cLHomM1LK/G+YAikuKQVW3fjbV
bEM5zN4sUll4wtkf+f3g5ckNuo1mSzibqQSZoDmNJITfPtzprDxe+BEnbX3Ea7iXfqGjZMlFZCdV
vRly4TuysbrhtZLx3PBZqjpPlIJFkaRISIiKnZpxK+cISNYJaXfy5LCbuP8453GAJJMkm65MKui8
Gkeh6JoOJrtpS5hGutSzqyAmPxKNpNfRKpDPRiXa35vTjRpPABpO/K24hVnCJHa5L1CiuSTcNWE4
wClWGUGQbwgd+7WL5bEGzzmA8oJiyR4kGnHPJWOCG58gvQnFK8VKtAj3nyF6z4sJt9hM2+zd+loS
Gi8CA7V20Wl+Z+2fraPq3zH9s6QR7X5N+ISOaJG93EYi7TNQ96E7xnLId3S3APvPecJ56d9jpiEg
EmMbiVShVlrmZJ3HsEJ2Ch2vChcSD7lr37nmTwNMPaPxnvWlg1xOvpq86V5o6WOpMd7WtJUerGP0
SW8HtJ/zcfQeUc+cIntleIUiKUztcIwDStYbdP+XyFTDm30BdJO13mK9CMUhh8U7j4A7JzibMvuU
Y5/oTFuQo4XJfSOtVrXCkFj/a10bmEbrxlDBHomF5hKhCRsmMfaeds9UYXsoqW6iomVk57P1gEEy
d2q8wq8iCXtc76vW2LWn081NrniTKJ2y+xOxWk+Y6pRq1IOigdhk/NAeGtIft9FmotTrns9THTNS
4ovgFBgEwpeS1bMzhSPuVthVbrWrkd678Q1IYgEsPKWRmPX9VmJ1MBD+IqlfxjYS8FfbQoEuc1X5
SQb/idCKszkXYNJsBxXyO49qnOkpelNzfkZqZTYMoUwm6/iGxbRar6Zz8gOqor0xzP+0VhCmYAif
Toi+5KjTsZTHweTYPx7xhy1iSOWzATQyuARWldXlCSXsJU9E5OfT6dueexyCucBi2/QbUNsAjOqr
cXnlRlRbwyTv/itco051jV5l3Aw/Df8bbJJQdumON/onAhGi0Lsd2vb6OqSdMDBmOi8aeo8BlmZ9
0zpR1hwHolr+BK58oOxgDbqJww7aas0CacsHh4eyqI6taK+gqsIG6kjKsnY0fkJYlKY2/7P1cIV6
tbws/lpFZTNUKtEDXXtwyzkNQ4eLMJNFLkL6x6TujMb/ZAOXUW7d2hlnbPe07dO9IgMyOdIOgnx6
XpBqSor78TLZkTGdsxlodqUIi4h520Ee8JwUWozEgeA5al74NwtEARYA2Evix9PdWPmiAamabnVA
GNs6XRNshMLOFgo5TiKvA6ptn+R0MirUNb2UF2PkkblPI98MTqSnrJeyJhMKl9HvZ7ShceVT5lKM
j1D2mY/JpQqfEDbjRbEy+XpZhyfbd7VkvqlqMPp1Blm0OsZWywLlqNv5Tca8GrrnpuSxJP8TTqcC
52ez0a8zRFF79ZT9Rruq3i/2tY8bwSIx4RUo6X08Q183/a8LOmrLiKvgf7z+kg0i/8TQf0pL17gM
DEDeTd4bd2qFAGY+lxVwrYWyme1WaQx3HxtGFApoosOP3Fr5N4K96eWqb6IMAGW7vnQN/enCEH3U
P1yYVPe5NTyYSJDCbTZkg2yVR0Vwl+WGgakvhydYlhx0sIPNAYBqFdXVgNAXbisH4i6nM2HpUXIA
PCUNWGkwrPsoT2oPcjX0NjqgB+H2VfL7qR/z7+eTvYdZxz0bbVw3RVNA5Prd3okcRlwoqAjaSVLP
aSWhaCnE33chB7/7AuMWqHHmJ+wQfoDiUix1wFKxzd9Wmkj06Kp9oyZf0e2UTxaZqkM7jz2h9E7j
/5w5htaErxcoB4D+cdVGyCgf5tB2VnTeHOGCL3KRxOPFuqA/f9uk6422T8qy/hyBpNyeMDHe27db
A0MUIXhofZHD9bsDlRDhHNNhOEToF5sVG7DLl7etxn0U9wWqBD3MMH3U3aetVpfN102U2suwkF02
jNXxOLhsZg6IAElhXv1DSRk8boTUiIng7VsF+J2DMYefK2IdYE9D+g3h0fSu7mhjJg5me0mAf+Tp
2ixEBDadL6rGlB5GcN9M8O5yZtcinSAUAIBhMdKha5rrmxfvtksTq7FOFXiEkzvtPFRQjA1qbJVK
I6SNmNcmYShFtCYfQrVZ4KOCrV/Hq6Ymk2EXqMS4gjJni4BdsK3xAXtvfTmecTs2RKVrc+pPcfGR
fYJ77/JU0cwfRBVkaAW8Ef+LRBQvWQ1Uujobl33/g4q7j8rjZPyLnvjaZMuUkii4gaZCQEj0pWE3
nDE+arq0yicn9gclPSpCNktbuWJN0y/z5BdNw5cbwADgFnFi0bII/4gSMW668iNtg/Oz56ZE6H0+
eRNdU6fxHYMjDA38vStEsVccLG3PU8M9dEnCBHacP481yPU2vkhrvSvvU1/2Qj7TTvkCuzZXUE3e
OhUC6HkNXXIJZ0susIz9tTJbgED9L+FBG5jEcodfga0uEMw2tJ2EfNvXs1TyBIkxSuroN60QKwDb
ZP9IPgIsc89BNWRmvalolz/rZ53MuobKQYORVuP82EA4kfwu2TmuJzH8aAHVmyrGY1iMoxxakoiQ
cW27I+VUiwwk8pOt4RoOcMFsYFC9tt5OUawU5Mpo+yS1sPEFIMtM40+6Rt3SpNLX3st4JzmkaSWd
EVzUMX1q81wdFkAQOYWuyOflSwoAKFf0BXvbFn8idd/tSiEwzuZVdZJsDpCzc4FumckoLWS02ydE
lsy2p9E32Ns4P92S/o6ic2tz5cC/bilsOSiX0YjwqoXetf8ZyY83nO4aTVtpUS66KS71eNZN8T+8
yNHZP4TNYFhvoO1rV0KpckI360bY74Lq2IaE+bW9QXmwDJhkRvk+Yd+G6L7H088LCY7k2eG+67CM
o93A95TBnKy6PZAUV3dv8clOAbezLwL9s+k8LVAULxgHhvGtr+HsK8PMcLPaN/Vt0/twgBX16tep
V64xvKRLa2J8Lyn40mjCJfSAY8N+yFce1eH5ykhuvhLVVPKBg8d2Rje2wqocP02pjMT6/k5oaLct
40snRkAwP1lxDHzcIYP4e9V/HuJlu00Fk7PquG/zauTl+zZidtmg7hfOPW/SkUncPrmfLN1Fkn3a
sTTI4bifTWJOYXWzP/mA+KFrmSLvIwGncFNG8qLmcQLzueltkG66/LUe48FE7FA4ENefq8GkbG5u
+hi+KRnDCSvxnhk3MFxDmxDomwvlx7uT41o9t4IfEdNlpTU8tWggj4QYNN96/enW9zwQFb2soeDZ
Uch+sZjotc2igPPmXyByF+fkkslpyFPw3n5Px45GrqSEd35r320NzyUJ5iD7RYskw88ZrAZUd/uz
yHYVPpnUA3rg41wh1bwK1x+cekURTW31x0jfWG2XT2uj04O5Ui2NVBUEVL+Mlp3fX36vB4KB8CR7
ioug4/6rjmIE2EnRt+KqevVNy/tyCPFymdiJ735HrknsyyEFvAxWQvJ0t+3tMNs8sdgsBMiMvzOg
0R8ZXFxgYkQHvEKBOYW8Jf3IqeGrysQ7GM6UCie0QTFTT7SP97lEtGxTrt+l/FuMRaOZQIXAWK7e
Y4EAU1GJc7e4wz/qT+/Hjfnpa7GBPnPauvjszxk6RSAfbv6vrbM3I6vbj24M5OWwP1ajNbZp8pON
NoMv7H1XvwC06DSOmGhc+ez+CI0DcaLh0+TTS3euk7gHVZFMWQaKNkN2HSgPNxcuvdnBt3A7AJ24
6rhS9vQ7RuxwnewCj5GwLwBLWcpwLyyLq9OdFrFdeH6RxS0zLPZoGTQ0Q8froIVFDuYppHUmObiP
KPhc6wLyQMY0zaVqAJ6iyZMLfJ52vzUy4X/hogl3NhCwepjARaT7n6swy4z0nZt7LKH5aTHKMbZc
EWQh+VaHlEmsdirFVzkYV1trzZ1fZmT7LDiynIynQf8axHEfLlFwN7qgN/1gY2RvBsOaoGyjmq8N
1IDl+bai/6wZRTKwkYnkPzBgNodHe01p1ha7He0dBjs/bbzMl/+VioCbObyAjtP3DoKsY9/DSIYx
4+7a/Ejhxq5/EKUmjRY1MBpw5ZPjygHiIDyaM7Ughc9CnXrVC6bf6NyfE/W8PWP+kO3VkJTNjId+
Er9Sc9Q1Kq6c/Kcs9NSJQOF3RuUutPuYeueixIB09CQj+IR2Gqkmpc/5JnvMsh0+riu5VfTMe3RN
d2SHp0M6AcetlrCCls1UEgC+G59zt+x4D3VAxV2VFHa9hB1R43UyHhFpEuBzMEKL0Ll2oEgRUYaP
FFXJopJrOo/6Ze1GDUkx5QBZRF7Y6ovr+NW5irnY1BTeseJYk7zxeOE6TkPHlYVPqOmH11CpddFs
J3dXusQAUT6YIs7Grr69XUiYHpwGmGpw3dcdPgLJp+U68MFYiUKhpjQX9EuvM18YrhiuLdsICKNS
QEzELCTWKVJNh0Z/63Qi769yVd9iC6pttTM7iMO3TpCf7TQOZ4fVyLUBvk6Gy18cr3oeiCXCsZKo
KQlwItXcHvnv3IHaAzs3rtzD/hzIbYNn882gXvrBch9ETasb8kuhgvNEhPR8RvV9v+TIwmBniCwP
lh7lxUanCRApHK2bsoqkoNPEMInlVrGR7ZlXNy56576D4qgRTFS5Xb85kr+WNFS+Pvh3UDweutXE
f9tfwnWzFWlP2/bi4zcqCNWY82B9TtpdDEqMwC8L8IeNL6t6o+aFFC6Upqm4GQXMpr9wAcbbDj4V
f3sEY4EvgsAIHYwlfgfmQiC+Qg3DvfJ1jLggyX76kjrV7LkaWeMcA6pjxhTHxmpbpkHakeZGLVyx
eTTNt1zWRKphXOVxMEV90Hs15S2wbF93p3AG5De4aomxwA3YDty0cvVlgZdfAEE0JCwzjXH7WVtN
DRDS5FeFVX8eJnLPjEG3Xq0xtDqA/ycLRhTrUJACrpNVixfUzQh3cDMeXw00BPpJlf1OMYNwgD9J
UgKG5GXOAyiie6CxdltbjtZi364zl8K4kY3O4ToyoSkOLVlwW3SLVw8NKjXS3a5a+xlin83GDnJ5
uWuhFhtAC8tCd9AMINK3Y6PGe65T4PVkt5BCNjObzjJ+YLhXlkrhczBp8d82hxvgHSjgNmbLEEIf
9Gj64Ttf1ssgRp7bMZ5melNC+uQ1BTO6vu1ynTh150HWxUg6QiETkdSHefFkBlNcjESjaZm8JcQn
Y7hfGM9duFmD5brjoTsCUvAMmiZ5O0cHK/ULTBEGKXAx6yU1bKdENKmdqS9Bxi4QZfvJ396sfjNt
dcugpLvpLhH3F/2qOw/cvnny3bvFG7Vv7mlOhVCDGDAOm3+2shEbE0P2xLgNAlB3oPYNHyUyRK2D
KVBRAuUMWEkIVM6DTmZ6e/8eio03x6VOeYi44XCnmIvPgajYDVMswzVqDBWTX0LymNONBQdy8jgE
JNr0Yi0eP6w8Q5duuq+sdZ9uELF6RCMkoqxzZSWTLKvRm4nLrycSIv3ONBoLFtXmvDVZVIQXjO+R
eC0fJ8/yJGL4le6jjjKRMEwApM3Lg0XV+3SDVB9UxRXdsicptckpdDqtOTMdxGQYddJ9Zi2xstyS
yLT1toIAA2o3LA52hM1UZ8zX6ysD4BugkjSv0V2cXaJn9bhjQcvDwNRJC6Wx1FYKtrkJq0sHrTIw
0uPcJMHu0+p4dnzXuSdeIYeSHtkANOSUa01uCuJrz2jwNRMVeyap+1MYl8vXQvgdvBkjjbIxhvkP
cZixp/juWHylQWbN0oKbJp4uCRqCvO5Pr91VPQXxkJLgiheSWAGsPNGppMBPOGc9GH6q9OXmWLmm
PipEgqnN8Cvn3x23NCCjoumbi47lXnyY9IG3IjoKhZIGo9QsZYnAzZ3J2+TBgVTcLZHWDgIWID9e
G+rwim3VAtIgymEOu2IlSGoTyxccRcP//L8UbGreOwckMAZITm6UrUIw0qlQzhFxpAtnBwjEp/Qk
+/wdVtHKRcXmsX+gYpJDEyFFogbGZE4s9j51Vak4xU6NcE2o5cahzgDqpSdVZ4JAQsQTKecMK2sb
x4HTTdRSQlczGnxMasACbZCYW4+y9hKdcEvmxGfJDOQVhwqoos8qbQlR/uHn+OcbxdPEk4AYmpRy
QAfq1hBOQG2mal1vpfOcSjgmTQRRwpJR9xUrB0HQAqLVqqmE1YwHl0LPlwt/rNOsv4gW+JcxqZYl
KaJ24Yh01lCmpJEmTRcmlworF/QDWvUMvuQoP2D4js5JC8HyK3xMdsKEvCJmtG9x+yqn5tXpcjk9
RjlsAAs/09iL77oH6ACHZFWH2su7zTxv0mqJmURbMKwy94zCi592C6FgQY+EnAJriDp6lr2BO43N
25OaBDRsQWwpH4d7rKNK48D7CK5Ks9DWjjEQN9bx3JBSCtFCP73dzbbjnYM+3DM1KLQVcOr77LY9
mIz/zBknGiIWdLOhjnYufiD0LhcmwmDMLIYG5AfmKbL1a/6kHucV3GNZStfbTqJvjtPFyGBC95fO
JiohLTWlOVPRtA8XpyXTOPfZDUU56GTV17pwRhPPo/E0WNwF9fUAZ4F63dmUoqs1X0MzXM/OuTRv
t34A2PtYEOk9KzHQhfgWWdpX2s8LqnnZXDGVzxUWCiT6Yym2uotdBawJfKgkcDeBric8kkRKGoqB
gmPjhctKVayetJSkIKtp3F3c0w0Lvf3FQVTHKmeYr59JATkccM07g4M+ETTQ9c2D29+oZ5iRS8na
/VDBMi8/zUR2K/hRqhEX6xZgeTTHP5j8W0jTv6w0Xu3HBmRgwkbH0+Oju+WTxlPG8Yj2TilzAMoo
G3SmJCaq/BJjEcz34DCCrLLImeYt/hE28k7T1QNtpgdjj0RqW/43FKMfYWiPHYU4hjNxj207wiE6
0QAMhHVWBdtkEchTfNNqd8obS1g9w2u95o0XipvDAHmi7hiX+gFV8+VdPlpHlUqJXcT/A9WpZnOd
Q/Yb1+R40r6gce6OWAl/pWj1neGwgSMD+1tuGaBnDj3LaE245rtnfN7weLUBkDwp6GMpcD27xsIr
S01Oc3ma6kRbhl3SM7pzGvYN53AygK10X7BcCrJGocEUjufMzYpu/aBoUbbZ2afQtX+XUsG2gnW7
lUHKZoAB8PgDbKCBWxi8bEFg8lx5R6FAMjsaZv+sn8ZZim7OIPtEadZ/8LTkwNpKdp/0QpY2xF5y
dVwHvQ7HShTuKQvMG4IZYSX09RulGGd6T2BcBg8N5m6vZa39Z7qTN5TTBBmASrgMN+LBHCdGx3gw
SY+HF++wjn4jSSUuO7GVIMrO8PaNFRZN9VN0Wkb2EGqeK3AvaWfBTu3A1tNOMe7lCIVNknVPGiMx
LuPEYPlwvDmS9HVr67WqpkSCCVxiUGVOTGKUgY5ECxI7gSG7Bcoakxo1qxi3Zz7ymss3X/6gBonw
YjlUe0PRS3dTTzIDV350lU8hp2fVzAE5Ouagzoz+6X77fMVu6IoRD2sNcT3FwUaoiWu98u1cFayF
Msc3zYCJXn9Z38YUn03FaXdV5yJJAo+x4iAE/7gIGlowgy9JgdjQ3ZNGiw26X4IQBdQso94NraJI
hQM+9WjmtdVMgGywkV76glY1zYQEhcMR44JgA4kN5ldlh41eiyPCNJliXCas6yWudz4p0yAybOdt
ptA9qMjStRvi74YaLqLoDZqXbDX7oCBs+69vh0YLOV3zO9rY5uRZ3zuFM2vU1PuHxQlJkBIA7lZk
bVDUTe59skUCNPe+mvHzWBkC0xwLUV7gJCvOTOnY/lmK4BluKu+NSyqfNJTUl31nFPYgZ8Ugv4ny
Dz++Es7clnj3yb5Tu+PzhQcMANZ1KVGoaCW2GcA6aOzlPAJXfRQkSH/6Vb7Xf8xsN6o4srhSIXoq
FgiVISkocYvGGcWONf69y6WS+gOr0eVMqlR42yo4JsM+N9P1/GrZbIWJNJ+smu7Xmpuy3+GOTRC/
2p6zaXXxO4tsZ44ywE7nC7uLtolJDxYrkHebwmVXDW5QWEJFWRwigQtgAcUxIAMV8m5GHeUQTEs0
xXZNVuFfej0hBtAIiw3JwlXEeEDlg9S+Jf1mE7KjOK5pggp662G0mGXUPNHeG9mK4rWpxfNnCeBs
GqXx7SRXl3+VejT4qkdiwHAUG/8xK+/j0wCX5LM7LoMjp0u5fTO4/kTRyHtl5F2K3cKTWaWQNjlX
bDO7NzhS9cALW2K6uBaOhGpr/71fdyxDqvoXKCuRuyeCu8lEPn49h4harmtcKyv62JVuCaaEMQgB
qgK7PVFs+H6Vs2WcbfTQU1dhVCS6uzyWnYSOwAPX3VIsd9kFhkyAhTUfzZz124mBpxDZUsuYMmPr
pLmgoFSJrpOO6p2EByQJQ8Xo8bXuCha9S0O0G1mCkvL6SZpvDlZ9HIpGrddm9AWflNp2uwpaSqfO
SgNPFPpyuMZJMOX52MbXDXX/1U/KMF2B/8y1Y4cYs1uFI2lr/5Rff4ub10iqPj8rIU1d9oCLuVTD
cVDum28DUHoGrvnb/HmOHS0k806P7xNLq3ndSFwNulDyB4dcw6hG6SvIMrdENtGXSnZKDaXhnR65
xa4heiS602mJlk09l/T6VDSAPpkOWSMg9ZjdTfQg3MQnd981dL9VMEUwN8n2YtQcvJ08E8RZmkA+
8Vc/jEiQXTPPsBUSC1Qk15zWW+Sakr+vsleJt7xaHstKMU7cmZrdtQGhHeXzILu0KlXsLBe7N/Oi
xzs62mEn+ZI/mvF1xQ5W+icKx6X2jESVrBq6aljrs0lIzF3qvXAPskjsI9hb1hGg37z5oUJwpQYX
I1FCP+z6tRiO9kZNQfLEdxRikcEeDSN1PCE9mjs0MYOmZr8EBhchzO8fYtrdD4LF9CidrJaz8K+F
WwtpL4B4+G4qyx51XCzUEnnJwOauGKto6UXquDtmva6SdgpzGMdgnRuHQ8x2gFPTg8Mz3hVC8XfZ
rllsVNsOBC3UgEyhzcwoZc1vsofbOlYZp8cuCRc9PPPnXpl9Kg72z/qqvSxZuH0BAXt6SOyFs/2L
4o8mCGAB2AYP0tjFMSq5eYiNChu5bK8shh79fGuqSS7jPuXxF2XPlZhYI+KutRKVXTYhp6RDmEEZ
UyfXTbXojSI9y5h66Agj0s8Q9f+rfz/3hQtMfKDo1DLb6K093GRiJSP2bu0/fY7Rt4XMiAeUbOWW
5kJSDS6TpfwLpP8bMtDN+hbAGh0F3VugyXUFgFL+QjnA/Lo6kFPaEHb9gfIQt2xp7OqN/hTXQYKy
ko3RjvQqNDqLSK2RXOzQkqpNucoBm9MZlbDScHiUuLDvRwjbX8CfjUc/GlOxdGsrlpnFwVh8FpUj
+wX/ioOaae1/iCTgZBGF7k2fm4ZqHK+LT7LVNuFKuft3hYXQB43bJPMXnzysqbFXZYQCHhuqpWlU
hkro+uz3ewuOH5rQ+vdKera8mw6Ww+dhhFnl1QFZAHK6X3H88LothEl7RQXVTin5Ot1Jx1rhbi5K
cNO8euK5MtO0aPtZSRJk/3MCBhWs/6bGlre2AYPhbI4CY7ueFfnSIXtOn5Sxj2s/Xdio66aSx21D
dCyqh2SbZ3z/FHqEdGKj3DWM5o6cBpxsCFBCS0T0I2X8t8jBglkibd+SAp9isXUOAqRnQ3jwtQeg
nb2kSlEOSb10XGXLBIOZRheAEf/LTl7qDWAIS8GWvSy5ZUPv5wDGytRogda2HCpUL0bRK4z7BMFv
8+5+c2dr6eOqI72akAs5qmFsNoqPsK77znpE7lGMOMYpk5CPCnyOT1kSAgKGvMmjgGnFLfDb9XzB
USSWOXtIbTCalZpWeARHKhLC2jTmw9pGkqm0QEpkgEObztXI6hQ4LbC3v4ayt59JVEwCWZ1Fa+kK
ps0YevfrgKBZtJwHhU1OZkvsnuvVDXwONrDct8+IuAzdGzTCCgc/Xneddl3XIvsIFpEoXXMcL3cv
d7MoFJRnwyKu2FbJ3p5VQK+pBv3x5ymvnVTOw20NVvG3wXUXmf23dBGPQJh+LOy7q9B+mYcvH9GL
ku6vYyH/0uydSkCYprGRvxOEchVOqiAbPqQn08g4AEp8L4yktyB0iaB6a+2Lrr30RNyi6pkVN7wb
Hs8z3NdkN/MzMeoWpiG+ehYCLW9sfyciBIIwpXrGRydMoh0bhEkrcV3l8IXKmWl5GWb34Z5TFiNc
lnQnT6UY526VHzmnzImYjYl1zP1Z5vFp9ElPNuEDAuk2PpZ5+G4p9QTSI87d4iSZi2mzJ4sVwpR9
TRs7IWIsRfbFQXnKiVut/e5oaq3qBROKV5/MdFjJQNPRUmxOuT9e0dMffxea82JENYmNxgBnNcQV
Bwx4dSXVURG1v/e5CIuBrRWOMoPwmGoiUmV7V/Wzk35L867Zl73ILmln2KqFG6SLR8NL6rPg4iVY
d4+3e2tvYzbzkY+rsbXjYnj+gpEPPrvbt9yOGoMaZBKt754H6MEGQvdDSAUtq5Qye+b2m156njXt
e5pG+QqKa6l9oDI2bM+az3YRwUqlbjhXMmIrm8Ad8iD56yJo9r1B98CZaj/gbyxwVW2UaC6ys/b7
LdPrVCugut7oboRSepHQGjtwkwzT3VYYI08WKvU+tFF6baOLo53KeCVQX+0JBJlO92i0qWZ2yO7C
nFvKN1qGZ2QyrnIbNjqF6mnui8NU7PmIdnpn/i2npTJEYpjv+Uy1H6uBsaVzSQekNL3vamAmcSsh
W4PyusIPdxdBBhffoJfECC4sEMW8bShJq7q8x5Q/Nrgx1RfJJYm9ZCVzaCFwoNdQGX8A4Yajm/yN
Hc6zQ14xQj0kRJ7trBRdaSRcBeYkGXIer+ng7ZJLI9YCU4DmMd4oWbNm2+9gn19NynEFFBEw6yZZ
0yLFNsMGgpFbKSIpkVnldKmkUvTc5xQO2x2en9DOEm0ap00ORyt8Z+TkKNomgILIS+Ia9p/IfEJ3
aCJTEyIvh+eSDQlrLVKDxkUxVvQEJkomXmRAeEqSdVbbMnrLwYRCrjRTF2crcBfcDg1LCS1pINdp
ffTwpSFMzwbCIugy9gi1q66jq9WXmQD+DA/y/CDuT2BgU7GavkCDlxo8K/ugjAuesMrjSzXjTRLR
u65NG6mhAROI87B2a01XNwApBDINufQW+f8artENI7f809ltObTUuWBT8hrfQ6URDx7jbyVtQT7r
EZZm8JolbmNpNlhygyfKSCxsEkuI5Q2XyiSFEJ/i5DH3JP9FApPtpcu4XGDvfgZj013HIiINdW65
6IZcpoNt3orbl5dt2yzr7eGgglIDgzf+RLwpHany427t5vAi3mT2rsPKTX1XtjhqnI8lxC7LuaT5
W4BQSOQi1ZMH88XEgwSnJFZ7vJ7qHKkoXOPcUBKEHSuZvPdFIUUEq2Vn9GsqEDoYwoxvtG6K7Ef3
dSRM54Lj14gZKbEYwk988vOwQ3JR3xAEjK8y6hMfTUmpMWDgZA7HJPldTVGfJKSMN2a10d2PLVgN
x7tA+K1xZjOeKc5uF7pCg8GKH6Z5DGuAEmu/dP5np9I83Yi395mw8GBKd2cYT9uabvZhaEP5VS29
NhcgDs9kTDMCIWSyrwhGbUwzeXDC7iCK/bkA0ED6Y+vk43iz1ivwLUOzraItHTmKwqBxHFUQrL7Y
5M/DJaY6KXxiRNGtAgv6cyZ/UkNYkickKJmvq5AlgVQ8A90nY23m6JAQeo1oRZKGOESBXWuHqJlK
TgxeWwl/LlxWWW5FoCC8F2gY/0jYWtY2eE0UPJkBkAv1Llx32HwHFIre53/Wt1ku1WWrJw62F9Nq
RXylBKG7OaSYIw5SM9LzU1K+bv+nLxCbs3H3EBXb2xKT1NLLB0eehBl0cY8KKJ4Bx7kC1kIDaV26
Gp28oZuli5TMbTWEsrtoZEVvqOO1G25KVat88lUGS2ZI2xCAJngHvqbxExKl+AlJQBQyL5W3QgUn
sN2rqToFG9yhKJ+Z/3e5g5uc/wQpuDc+jwjCzKzMTHQu0rDoRkqzXH3wF7onuCYiInM0ykkE7wFC
i/dLrO5ptmllFvoKxqSBoCWwjlfmz3sxZUFZCcTZ2dMJbuRxlMDQymyw9SmSOTDUD8wMheYj6K89
yQwWkaM4tzIDQzr46ARRpPpxv3LzhI9vJ+IroooKTnvddIscBcK9wf4qqDMmB8wlHoC9pTtVQAnj
qdxwk3Hls2x4d2VdtQYCPHa+SeqCu9Me6wYcOxy8mJQL+8YyFR3LeCapg4SzTFu9dRIMvtL1eFwB
A9xMZnA2W5xwHQuGzRkIz8hq1KfKZBzE5BpJUGqho+AacFvvN6uHvKD7Uvbp0bXT3y1MAzYJq7Xe
tDmpPOVPg8LIuP6H6ZelCQOiYyr5aiVwFt24pKD3opt8n7cM3rtbBsiukGGhB9o3xKhBWkCnaJIM
LrZkaYYftWt9KxfYoQ3d1swZgWeQj/o9lCFKWLoSVd6GOvBwr4O2L4BEJHHOSSPhyb5k66X6fkkt
WQkkAuR8VU3iq0xeKxvZZlf4G5MBzCIWMrfNp3NTea6QByUOOsz3Y6Gl57hIg8HQLw1+Qw+zrmWS
gx3uAG7QPt/G57z6MoQvEVX13HVAgCkC09BFjT0KT0wKvMKrLie2mRN/RUAZxIogtuVTVOZ3UX69
nO8syNSgPdOksqLnUJoYPBGnUH8Yt6DjMcoP+5/A6xdFqe0WlUdqhyIn5B9j6w5wOGmRdpOk8bg5
HDpCV6D/EYW1jECgEmthp9ZX0QhPrLI0Lh9WOY+dZsl8FtnMJ/FhclBp+oTmmCmeTnynRM/3nGR6
bXW2hPSD/kF+7s3/EaE+9bllF41nUY/xdbanzgGaCLPeoSvX9ZrSrA11kU2PcYVhSGpnv3A7HC11
j6hS6EWjKbPXbUhx+SUgLSOeKzwGNIUB/oWhTDNtBPwQgqoLx6s8opdMu8tUBxJDY+SoXX6mavTf
ysNKGltQG/Lo2XfZQnesIeDTx3v22pZ0H8vSUAmLBsx5Mh7be3su+vjTC/lzFv81QPdsfuqMbJcP
GbA+Gbqf9TkDWH+dZ9SzHSQC/aRmKw4IFSWeSNDsoDWXfYDQHJLahFpy6G3XYDVj4lprkv/cZKpc
1JLWkYkKTxv/okMU0IHNouT82U+FAyJ/eKn9IgXHF49hXmXtPKaII/QqFHCjzgTN1t0TZ45tcMWB
/ZFoFOppLlhUSmIRXD3p7YIN7hgEpKLbqAPR3qSqOyWxl9Bf/Q0Wg9YjuOHeHgl95mEfh1R4G7pN
aZArJMzySuFIcORjFzHRNU/dLT2LFzu8P8L59fI6Gxlm3ScVT2oIkp9GtY9mITLP3RFr1bxmyGkv
z9rxcTSxP3Yp3HLaoFP++KE9ZQ/A28O9oGmsA5uR+25LbfFTdliWjcb7C1Bs6vHmVCPOOrZse657
iZqcGad/Emrho+x/7NTTv1kPtRKyjKadjGf15F93+E39L1HAJ4YfmjtbvPj4UOziptiA1eIdj/nV
BN3koR39gWkOeLHu6c6KXybt2Zy7OHOF6OW1B0D3nb2W+Wz2336bgYWB3oZgXMtclfhXC1F7S/+o
zFXEbJPP9pRCudaeOJg7CGTaXNCZlwmgmQdWRqu2mT1HGaZU+GDMeT6V7igr/a75DLA9Q0kjUx0H
xKPM+Ql6Q6WlYIrrGXo8LqTgxd4uqjrob5EXQafT+ArWc0Q0uYoXhxWDKyXGJR9hfRxkrG49fPgv
b4MSpNLSe7vfjAQXLVc3550VvV+ne41WU9faX8r9lD09NEM7RE6gGGHN8QLOEgOK53cZaDK0XS+0
AqKe8E7HodK5T8BC1NScIinpZiDoXmtwrgU07x5iH6+9WfDBuITAqP1QJLkT1hVAPbc10WPzgwMm
+xEhQkWp3cZH2HFNPsMTEK9/S3xefQcEtgEguNVPoMzKo0zhbu5rbr/DFD+5VFpQ1NfgwgoXHDb9
smf0+KAh8vkczZ0vRHqr6idIP1Ye7nLa4GeotxpvRcKnOEcOXiBeiEiqt+67ueRDnu7cQ8fKusJ8
ud1jtB20CuI9+IWXaWP/wBSv7q22vHB3pqz4FyL2RAVSYUmefpndBKTyuDrtJ5PZMg2X/oBtdCzM
MAJuacGnrZJwkbprYKL+etYC6XAwWNo+MJ9aNRm/b/bPBfTMCaPO3t8VBoRmKO+VaqwrTU/uhNDC
Umg+VTj4rX83cCt5DUH/YuRw/BG5haAwQtGB+iYtaOMOaMIoFaZX23xZ2FbPxijP+FUtgQmh3+Yi
MxH6HIqvmGri7hnA3W/EKVhgkJbs5L5lw9N4Z7diRnreyy45NWH2o3wfIvj8+/1L1pNECHUaH9L8
GEg6Ypj2wC4Ut07Udm3Lup5QlMTGaH7gfe4MsZaBHw43+vTyBV4nNa1GxQp/VI5WxYanJxF1ax9F
KE30G9xY0RFo4Zz1U26OF9Cahx39l2V52kDsuCTpu2rCofq0sj/0+IzKR5rbC1639VX4LoWRWFiR
ErMeRupKFzE0g4nFMBIJAeR4FvhuuSiAw/uzgxUNVxEWOtbX301FvbkFSYPToLGeR9u73CWTk8b/
9A5jRNoR9Rrr4Ov0eds+7HAnFYgrsD3t2cgCWTZZ5t5AoQLwlsldZcy9lIWKA0JidiNP4CsIE2vn
GIzGrxcc/JyAbpXeSybiaITrDEE07a4X1rKXABj1Od09DwIr6FSk5GWm9Gg8oEyowlvym2Nxxvmy
1AKbcYxzweBUsOYx9kUqmrqodxnbcvet+vjvEIs1LGhMn4fShtT7wQn05u71chLjyYP0QbcIweIj
KpCreRHPtA+rD+Slyumh3sr6A7cUzQGaAVWjiY3db9BowK5DCQxRHkpHOl6o7EuPudSl2W+OCymp
Swu2AxMVs5u78y4sxhH+1BxjyHmj8tbygMg3qcLnN2DniwgVIX0iUGi8lz9DT4FuqlaiDf6W+QhZ
AC2DX5qr7Hk7vZcKx8Dym4Qi08MY4TmVr+J0GGFFUocP3jMQb5R10THbXNFFgmXsG+Wdj/6u0Lha
hNjEx7fmylkwCzI4sRdgW9+tTANw+F9frjo6cFXsEJCMTbKj/IVGq56r0Z/HDApSe7f3F1OLMaL6
VXgHONlLsbU+GMqIhoglsBL9X+OqdZZmUFHuXczPmD4q2WcBhzwKcxz1se1K1Xe10imC6U0E0d0X
y2yZrDDhSAyLlOPruaWgw2BJ5uwRyPjZ3y6jI2VMfvMqXIJs9+CeMHdJmybqs8LYb7ewlaM32Yy0
b3iP4Atbu6KRWVN0N982sbEckwVlOzXMIsV93WFDZUTyp5ksPz/b4KdoN4xlaAPuGQNjgTeXxA8r
f5SYj3fhqbH0Fg9ZIRDZp9bed9cEX0Y6vXm/Gj14zLo5fPjtUawu9jVCzOtZxXfO+owjEb4RdkpU
3Il/pAZAu39WA+jwNbNEB3R7Z7Hmhc20CpIu+4yKA0G985SFb3ZDJsVgldVXIn6MCX+WzldyO0RA
Zi2YXhpkV+7cmTXuwLwn/Vj5PmvVrVjNLXQO+OK22RxRaKtWddbV2JnoWWCuX3stXSjkD1wQ4CQQ
AEONt+zl1uSq5sbWeWiuFKHV1ibO7m6HLobnFqHEdvryUW+SD90DvoQl6o/MDMx5wLsF9U7GXUtv
3ngnBGlwyKfBlHe1iwscQOEVp5U0jH1G8WDunWGmflnf8LeBJGgvSP1I9hmGPIYkQO9va0vayjeB
NGN4RZ/KaJt6HBU8UfmOrONrB/vtZjDqGaaGfK7vbyaUQtXFeKpRkHDR+PnXT7/TlUjflKjo8S7j
IkO1BR26QCOconmnAHldDPm+OMuZD6QZ8tZDYQ2Bp2CtDItTlGYVKLD5YXzW5oVI/V+UqCYQS/ib
oBVrSPaw3/GDA5ae2wimIPeNvPVtfabG9qiWp+VPwAUOAVKMmHrTSSU2mwA9GtG/rmGZ8uMyALDO
NE1CAABAGkzV2RY2xMDGTxtnpeWzuw1bVTdPizuCy8A/RNorQq+EmeFd03J4T3lMyTyf4ytgV4hx
1AYxe8RJm5Ul3/vNGDL9f9BSWlGlRxQx2zAi8AJ5MyHuqS4wxo1CJJ+25J/j1YhKaeeSzqs2wGQP
Ko6/t6GeTEX8CKoAWqyJkbjbSNl4U8AKQpnJmTJet4iKfwMdjJFy8ecZcK963BQdWcz/vLz9gbPf
KJBaWGOVjHO8vyrJkernxlBCL4c0bSnztFa3pJc43HJBWbdqVsqPBCDmdfHzslhSmtJmvk0ry/Gw
Ap1jmRWNtDsqVEn89iWcmnpg9gTfC+Zaf8GnLPTH4dNz+bxMLMthENOGmcByhprDnNhlGYteckWf
SzeNG2yuLfYgkdcdC6xyHUxBRLYIn5AsGJYDF0ufIJt2MxeH4qW0BGrhTdCHBgUR1Lh4DB26t7n4
8Xb0Bk6mB5jt+Ms2TFuGY6cS4aZXkybLjCkWjDj+KFjIZFaKcNkOjsOzusdFpZYO4QCjwbKtd4Gg
jSZV/6WYHQh0Oylm6RNR2mxfvhpbTNmpZdpubkzninFwJodjZPmpiZFLQSM/rnQFlGrFZNGEM7rw
FnqnlZ/2PSytqezMMar14IMrmWiGRvYz5bdLHybYppMkpZps+/f7mzeFghVPxGRa8lqzLUS1bf4w
c/9b1t+nXPBCY2i0M77Crrn+VSUo0On/niNXRONvyJgkadVOxqUP1hMB4GPkDAT+PffDg3buztpz
tmVZw0dR6R+u9Wwurd3Bf7WT+H41fs27ROdxdYN+CYikL1OKcmdr5rxcCOz3mGrrkrd4b2c2CDpa
Sf6cfe4XVspPhQoVvSmS/RCebDJ1VRMKSDaCZhz8guws/WAOnUFQyjCUa+tMj4wTBXP5LQjXRmhj
daym1Y4B1raSU6MQqLp5zpe0L7qCffGJaLJoI5LdDKODd4apAQoAJnQN+3/gCY1Nkro/QI+bhJ37
iZuGvxN0HYxudFMlWKnYEU//XOk9p7gbPyLKO+QsgofHTmaFgsy/VpRLtilLQ9xzbffDq518To5W
4C8sZkJOhJpW74MtSt7xmu0msQBBpH2B52a3vFC3bQjI36xddDqPiTGrVw0nbF6bsETiJaZXscKs
IKMWs9w5hfBDf9mveSZ6TIt/qXA6qemZCS6X29v+4XmvNRMSMeclinJ7708emEPDBftWe/1sR2Bo
o4Oa3xcwXFTactW062GAqdEbDfGPi43gxyBKewCssofEYawPNjH0H1RwaLTNEvpByfjQ4QBpsBld
OtsGcYNn8vqomL5mNleXmQaxVDVRV5uCo29cUSb3WoDCU/FawEUBGhzvuAlDLTc7a9ltqlgORg0U
YygVYSBjkxAkvs1/qr8qVjbqZpfhwKZkzt2QJEv96uWL+zwHavGwbcAGKOrXQHeL0BZYIPlq+jgY
grR63s/Rgam4v3yrKyZ8vUGLdCjfyeX7W+VQ6jVEMa5esNXFTyWUl79nn/QbIJXgi8C9Jy2KV6R/
AdQFVGT7rdLodoxjuEbJum8uL4Zjk4jyeSwCiseKnV/HpeL5jankP7GaBNx+GsbeBibMJsWSRres
17a0wBDC9lr/sXo+DSSbfA3LxdQWJOpRya8tFVL5A4at0MuZJx07tnCTOoSVNex9vskQpAg55Tqo
njVVfwbJHPzhnDVILSGcWpghUid48EeUGr27PAjqNXwlw7dkB9l9Wii6sRWHmK2+0OkG3FPOzA3V
MtpvdC6GjiNszCxhI4ntyx76kmXBNO/YV2Q60oMVY7OB+78cTGSf37kJ11Y7qtVXccMKg9waZk3r
P7Xoo/3HcvD2Btdipcd0lRRu/2H1i+iMvZy8w53KGuM/YupB8axmTLQMeZWYX68+jSETb5n6cvgK
mJ2CV8UPso3IFRw4NpUasiWbomh0l7HekuQWVRUyZehdAZkarOa24e5eiFeN4aQqopc5ebpbtXUz
Gll512oZi0B3ems4jdGBSC54mcFI+658h8GpqPqKvZbVZnTwIyuqUQzDOxVoD0luY0BuGGFc1FMb
/OY839xosbzyQvUK1l1Gox2SaYAnHSWFbHLV9EssSobuRWdlop/LUtCShQ77ah1ONmMyLYIV6BnU
D4ECuL6KAbyIqfVTUmK/J6gx8LWkdzrGyDxqos3V56B2PAwbTW1lh06DrJAKUg5RxZqLZYF6qdPi
hf2sSYoBTE3TuIdHbelK1LZ1snUqGMJTKRMUWa8917TsZoi0KlMbLNA0OG3H3eH7an2MFPOXstxO
LqcI0SnlgiwpQ0p7RKWkmDSSb3iV8T28tiU022xohHL9Vv612wXrHVt+8pco36JHRwZQtm+xwv4w
6cMJhjLgo9op0KMgUKPBWnJx0Ps55g3CUCO2YKm9HYDh8fP7gh5vrPetAsHf9S91F71H6iSMdsOl
W2lKnd1hn/VUOaDUucGVEYUquKxLV68Xh400k04UYNeOOe6v3DX39wyEvR61sYZyWoy5T4CPO3jA
7WOdozM75+5l5pVzw7HDcV6VbEFLxKY2zlQOCKTfrT4FxkDGMX5c+EHOEDWvaiGg3p8wqtWFbqOX
BHsAleGLSJtSz7OtPyAK+AP/x348sZxgrcsxH2vI7t2zpcOnXoUMUcseMG8O6Dk3oRhQcndFhE/0
zoHmJBqGD95KaCGHJUMHd5LnYpUHqMl4CAQ8xQiBAM1yG2xvQB6z9JgF39ydYUWVNNEcbwSIfFBR
XBMjJyHfwz2+VAHRpqdcJ/ijcvXRMrX49PDWuof9bZBsfUnULrC/dtAMTsUifB6RaVwg2k6/ljlB
5fBGkU3BXrNzCXyKYNOySnsHbNkw8fpIx9QpRIfmx8kK+jeWlclQWjeFcpFdZKB0TyoIQHLslA1G
WbbqNT2BDlcWGhHZhlqL+pY1rqI8C/6FoylAKILksrgHI2gwnQ3SeiFRwGNyvJghLL7sSrlt0kXe
+SDC0rtDVMSmHEeR+7IZ+ca7oNL82kTu2fSzQNvaacgWYWGUdYGKfG4y4d5MC4iA9JgoVRkMP6FR
35IUdrPU3eGSWcRXpkea33t7OK2bTSSSc9eydDfS2Q05uD2SuZTSLwGAdoFb9cSa//fYdALRbrNl
6EJdo9wr9UYa+NyCg8UnBdGx8iUVI8zagI/tHsCBXJJqoE1TkUctonwG6AcdbqQls8FkOIOkvGo2
tGiHGXIkwapAn3evPIZkkoIc8ldXcVNwTjNdGh1SSHkf53xFIxRhr6irKffKnysvYnUrArjVR0Rq
snKsCBq72XP1r1MKldj9oIF3JFmxRot2WiNNyPNeJg5/I5AkwViM8ZPYGjIXpZTL7mFwkp6Bj13O
FvlUpatBqZbW0XhGtbkyPa7AqoBwG+tMc5y5Y5DQWh0VSsvmCWjKSl7erVFedXr8wDcLYFJAxFv/
qy8PL/9YEvg9dtThFYdZxncKgjiC1hH+6DoztDNxTj8qsPNzwLVXvBi4NfUl0GGZgxxFTPgnL9Ow
5FpOIEt4cRELCFpVZuxbb56NgsA3wSJSuekmuFiM605TYtBWaVoooS/Nqyi+OujxCUd2jv0xXtlt
MNvRUH9W4Z3j9nXS/UaKGNTS1hNYPOJdZjY2xvoj2FSRsGCsYo9oIZSOf74CQu3wZbQbE182Dbrw
TkIuFBjsJrU10xZ7HX7Wa/F4O6ivgfIUZpjRXunJArG7oVAVySYAhmMHH8mPHk+aVBrHQ1Wl7qJl
+SHSvGqICGTrFR6UewDWRMt98dUCRFhlX+BTwxvkeQSuOprPiukJGFYPy5jdHQTACM93oZpBmvfe
GY3XO38ALRT1tPQ3TsCxcR8SVCbdYy/e+po+44rWX7Df+mTCiIn58aikk3wPnCQBACX35J10Y6vP
Iuo+2efxR0B5hnEO4nbMZ5ro2qDM+6ie29A6sS+52j6rAPJwEB3HERkLyx0ZRB3XGx9itdjoLOWt
SinWnhII7JjvpmoN8UlbTW27dO5qHJ0Z10/dv11KsYGslrep7xDOHOCDEZHd35D8ZFYqgi/27pUu
pw663GF2cYhA+V4ZSrOYglGL1gEszRKqd+o9OYEFBC4MQjDgjtYVvhY2yo3RPt2QcKnQe9hfLEMU
zRYVwtEdUbZAPh4tSPt8OIR0pX9ilvujwTyQFOj7RbTWkx6YkDO1uw+pcwA/C4bxY51aZP6csfba
cPZs9tnGOQTwoSfrnWQPhK7PDH/gQWh+XIM7Gqx4l5Jh85YCKvDGTlWX+WjZhFPCsfSeJ2D1ddbQ
cMVSkcs5jVnerISa/6I5HqwlZr0dH0/Lm4Ac8djFXdw7I/a2iN+U4ePe2HiPyUEgskVmwmOf+W85
+EpHNNabhGYyDqcCCCnLmezv9s2Rc93HYQVxny0F7w/1QYOeRMEwaJi7bid0IMueXb9nkASQlUt0
xBIAl43zfLmzaq8Bwtr7+/m/94FGlZzYPKODWq/5wPknRdYK0EFNAmUHZQexUI1W4ltubw3O9baG
/PZ5XeXJLp2AmxT9rOZOJFNAetMWJAYlSnr+tZRjbzXECCDmXTtEn00l3QCba8Aw/pC2Tgn1JwfU
vp8t+uX4X+gqv/iEInQ1nO8VzJApmC9M7SeMVtXy+06uQ0VfQ4tW50U1Bj+K2cmVpx9fu34eJDMw
+DtokdQ0UNR7VtYFavOPOSs5eIm0WbWb9DNfehZXbmlF1uSYwSuNT0r6BYoTsgBp+0i2hhMtM3fT
s1MXHNO5tYslGzEeikHWCAmWYh8n3vYvpwZv+RUGbuzVBpBXjYj7q8DKabFNFuc3KDT3HVy4CYdj
MCchgW/viRGPH26opu+F5SLwiOz8UmA5UZs2EtHmMVVeRPNRWJwvdxKqH1ahHsatfg3PWyWcqjPf
gq5hXYGJnhe/tlzi4+bAKkDMBUB8Ucxd3Zst6XBenBKN8kGiJ4bEy4n9KEfn5omyKRjk/2Y2Esbe
58Ad0kx4ulPBR9Fu2kTXZ/wuMcY3MaY3YED6Mm05PLMOvHKy2q2H3kAlGV+igheSPhUro3UQrd1Y
gVSy+DyGNvNdmMbV/uYUllHSJ0TqVsWTEN5PVA0MgXLGQWin9VAdn691k3HapRnUpebNErIpofe0
K0znNQKPcl3u4WYIBUKhu4lmJ1vUJRTSLi2n0fIWBpOuD6B47OKIQQXKIFPtzwFcq6T2UY2b+C5C
ph0tBhVZROquiKNb5u5AstyihA+VlIxuf7avGcjYMTyBdrWsyeJ89Ptw931Ul4USD24tdOYgoxZ9
Uz/bmdcceynnbGMauKzOUndTGl/Ur8R8MmqjSmRl48qgFyFaPlvVlXjNMLgE0J8n4xYiXORn3JDY
Hca8tDNTb218MCo2KKAOqv5ZqjZlU2U9pkEQoVQGV3AY0t6QkZr1Yxf8Jr5fPr+Tz2OwE3xj1/17
dTqMjAVSyOCmEQp5EpGj40E0q1fWLUsUihhetOHVick+UZfEIhMpOq1dtw5NZhRYmABIeBacrCSr
l+qF9miKmsFWIh/5dFqbqqGxq78TC7b5WrAjftRvkes5jNFd2ZJNsbZno3W/2CyA5ZUy3OXeLqX4
cIA1AYzfg70oQIomyB+UJ8RQhx2XQRMHlX3PpKzbloUAyIETbUhTYlluT7PiGzRXlhqrneRhQY5S
pzjOhCv/gW0RlwEWykg7wyFsVpkUFuSdnUGXMOBVlsmPX5/+/ZS1voV4xcaVCXJ3wd1B6PheLD7O
E88SDQ+hiwpd57DMF6DDRycGPEkxXZEobdRl2CkWyo1JljKZbAHlXX4uiJcolfKGJ/YwE6Abiak+
wED3yEsBtflTe+WoL2BB4+/oiVTnYO98K9mfPurv7GVBOCKHEIQX+JDvP309HWqkgqUsiAr0e2fg
6EtrS8l/Emp/d+YHEuwndNAbbSrI9RdRp6uduVMfU+XgBacDywbP9eka0yh00uzej9t+eDuRzeXA
Tlks69VreGMYTkyxeJhGQ02lzjqJqzOXHiqNURtVWArdlUDWDkRLxacEkSshlcfg/cxNb5ULszbc
6JwG67D8/ktV3n4Utdci/Mt2BLQRjC22YcfqYlZAJYYQXf9q/JbiBBsB3XcXzwqAHP+AOo9Dvq7a
Tr0gXtWwQzaww8uSqBxdjWrZro65IBb4x/nYbRmvjFtuQIpNZBx7qntupbAi+E9p5bPIWdZ6tnVJ
4iOAprmeR8uRISU2f/BWWgItMKauPt3kvD2Ws0q43sYE/YC+X0GMtPz18iHTRUhPKtlIpuQcy7jQ
7r6f2KhLhZKqqUxbux+SEKePZBcoFYuk7cNn8VZOUXx8VEgKuB7iNSuWzkzW+1QKg28ToGdDqnWA
5UPr3fkaS0Ary5BD7d0GRurt29aezjdpaPFkmPWTlc8tv3duciTtsVn6Yt9KO3Q4KaffU/NYfcvY
mBsNBr/iBLZyBEzDN5QhOQk8uk62fRMVscYPNEhxII97pFoYYC5IV8+G7mV4/SpbCT0mCvZRU3s9
tFtkvnFw+YXF8T1u+zKfl1M1ibvFVIgzH0h+rjLdtnMrKZnCuXuC/RqcGXru24GsuK8luROaYOnL
9w5Wc3YCf/0ZcUufrUm2Io13zK9VtveF76MnNZQ4JqA5Rh+g+lBBIFZUQHuNFkwsfvdnU35Jihe+
vaJx/EwFztL2/W/irT/NeB4IVmEKXG1nlllO2VobOQY8ONsNs1MaMlurWlyg06KQuyhABHn9r7Di
slXr4xP6/E2haj7kCd9428DOo+JS/Ke68BI19J2KX+s/6jfB0ViFGlrvft61hdi9dhAhTNfIWAgx
fmOrHgFU5rCTFv/kz9o4UXb4COUFBNs+fAnoZonRlzpKTAGLFF5YN8BoVMe3zOJXUiskQRqAclhK
kHIQWhppKDd1Aq74MG/5y+Aaw4D5K/spRh08GKiiWT9mHLGjAF9y+RLOqVD5NXDi653wVlgrt2mC
JRxbIDde4Dv+IV+s/1nkiFMCLZk5xFnBBdwrRrgyw3BzeARIMVHXCC8+EbH1q70R9/LVJ8aisSp+
Jcw2xikk9elJ8ueQcQ7T+q6WuRLvDtrRtZyxIWWaGy/C9qpsn0pCyE6594mG8KX6om4OBNx+OBd7
g97vGtYnUwcZIYJZHTY5I2cJ2twqF/PZ4KyXvq7j1BPCQykbL3z7fzCqV9kAOgR1yfiaeHmed8SL
kdIpbDTKpbHCiV8z+tiTHOpF+CPCpUrbbmI5dGxEUHaxsYgzNeEIev8NbiDSX7tRg/UjbS4y9Znl
rxV6LWom0M22YAmN1r+qwhXNK6596tpIF4z1gwDxTBG6QtnI7kow9Rvh5XbdDdXrxLbw/irPciMT
hP+ZoDspNY+ZC6GFQohD3AZOSM0+umBtky4i3bwBxp8QUr41GEoC0ZcC1FeCLAF83KmGJiaREucS
8EHvDurdcMepcovzyUrxP0xfNqqshS3FUEep63u3vwXsn+trbgLOLNPtWquELD4KtXM10fjUKAoa
E8JRsiYBkGi3F/i76Cv9Qf2+ArTQxbbs8qe5j9UoAawZcPbMkJUYsa6m+Pm83QPl7i7S7C2RToVF
2nKzmEn/bITL8yIPkGgztpFfJRQvG4nqNEPYcYPJRutGgna4EUKKB4dgxDRJuh2UmiYzz26b9KMU
yOCU+152ONmWqTGOE8RgkG7TxjXGI6rsr1hB7M87+24ZaJfoku60Xh1gvk0qKZQrAzcExwf9ko6+
e8uwKerL9TI6bMZkl9kydrxbTYgoeZEcbCp9a3pXAOAt4P/iJByHDhohSL4u3196bU/W1K/vqR71
fQDs6k8jGuOPGJF11GH7ZXFQi1BAG1gCmytMVZ/CIws/2HnBuQ+t8M0URZglFCyzC+N3RlT1Qhri
TJFwRh+dUvJpLzghGxOnm/m97oKZrXUMbrl4QX7YPieXxvaYGKsy72gtmkJRzbzUiO3uMC2bb/hM
LuWbhCjOT3fHgwTNiq6kasKlum/6owCuEO7KFxRu0+YlA5saHbJWaiyRRec66ipHYppIncC/D7y+
gmly6i0z8vB+7T3ZLG1xsFATHkDv2l2CmhK/2GKGs5JLdKc7yKRcT5Yt20BU1QdX6tgEEUZqtRNp
fjG3JYn8jVwAEbfo0mqk6q+ckVj0afsADWyd/9ZKCWYCFddT0ZYpVwZgdBZlNXCGiAk2MiFZNATg
YeDhI72V18IZ9Yk9OrJQEtZ1CbrwI7XAvcK2zaaFyLsmVmqOPMcJta4sCHjZT0mz/N09/oay7zCD
VOuwHQCtv/DJJByGWzEa+VGzjM0XLzL2mVd9EYap097wYqiB4w52CeENKGdMvFM8mAikpHeRQb/w
SX3GSjPjdIDN0mqOemXDwemYylFyAAL/oFcXkp346W74SZlTAyjhx8Fsy2H38N6mOIsErxJKXCwv
bQg7G8VDabHaCyRpEhii5dEOfdsPaUOSNY0IcASRp/NM63a+WWJbxIr6cOHuPmnqvNCGrSFmSHcU
RPyPGatXuDVaa5HE/5b9zQVwNkDNaUd8STZca+uCisboVgErddXnhVLcJCqy+OXkDzs+BVa1cLvz
MGjyMeXty+QAZReTYTcJvgsiYhC9kW1OOHliSv34JNggh93oc/49GIovrNTSEHA+dlOztN5YMMnJ
eX15fKy9neA9052eSP2HuFAlOGSrIG57qS/q4OZuaKXOO2tBz45h7N7fHopcljlNGlI2lgbhLQWM
QHzSEFhACqGPGDvExKZ8ahSNRaRk+KBB9s98IEDdq+BwkwYyOkiGovB5aR1sgqjHtcOtT0z1W0AN
puMdMpwBjYbxnbbkJ2cJrxGxvBM0cI1pV0Ws7mUX8ARXdxUKiU98+2yVIj8kWhMLvpXHWU+xAoeo
CCXHP9iybaYDeB1nm2t7Lf2b7+y/caGMnE2QcbPLHJWNw0I/+roBnmmi+HR7lQIXjRoVYnp/BCBJ
BPPc+iz7BY+qf5U93+hVHhjkJLg4yydGVvKR074NhmhFcmanGGaVSal3HoUeyCYL0ywKdcQm8PDw
qPXUZaxFq/tESATrzP6P8TaVaH1RJ0YqWDJq5bjZ9Aj4MFXeDa/GwgtXDOaCGrD4KVvkTmHUS2Y/
GbPBnFSkjluiAl97+akko9Ysk6ExUMuV2+SarWfnraJHS1vc2LcC2OqEgE3aW6i22tVcCbWjbMcF
67GmxfLOdElsq9cVyJqNd+efrqi1l8To7XRqGF5GlfRFAZQVymIvepUusvtBtXtpgoJw/2UZASpT
9hsrLIysQclkm80uHkzZFNjCpXWqqgejn4om2HBX9IdBauSF3dUb35e0RvIN8biUuBgb89P8nAh2
na6RnErQVoMcDJW5Kow1ljrXePlSLbnTt/oKlS5k21wtQ5TBgYSmqZDg1RJd4VtdbRM/l1cXQTVU
bylaXScexES7gCMr5g5qmIQ6np/COUWJ6Mqj8odc47bWJD88Uu/VQzw9LgwfwkgCYvinrn3+ucCc
Nn+U2y3KoPQZht+TrRXcjBLt4NI8W9WsvN6ykIeW/i4D34cF9mmZhpaJwD7UNoJRKjTEo2qe+naQ
Hq8iR7TcdC7zj1Q0Pno6pCTjY5TUWduG6EOWDtWdFiTh0Qm+WUsb9HM+MZOECB76ZrpjiqmMaEtI
DouRtgUF0Oyd1nkXf0p1ShBeGl9ROjCcOcVqUhVlHZivNjFEJjJOKjZnQup0C7687fGWAScxl6zi
BX7N9hfxeOjctS8Jlzsqgxz3sfjBLBHHak5mH5RMi2OGVjj/+kK0C/VFa7ciYm3o8V0uCn8SAEZn
JlTCFaVvthmqZ5x5avmO7aIkjU4FN9DJp/rVDH3Lc8T1ciPMecnek492rnycbqfrxpYjgO1LxiXe
TVbQ7tEBDGDlRCXOviXE2PZKlOWUzjZvJhG29k+HrDwfVwn9/zGaR3QaHAP7BL5Xa+J7YfWlwjF3
tF30/iEPVmjfFnwXYZ19z9xcJ5ZPFxHhDj2tOEyfFfiVgLM0HnvOAxXZYWgRDNQbyWdZXruHlvvc
TPfor4G9JvHW37JV4PvryCzoAqy4M+wgBDz2jJWRDAfZSi14nMqeFr3XzOTOVOhqnv4PX9tOWNHg
v8MrmHaA6WWDTrRMP8PYG2Si6seBoP/WXywouZ6iLc/4dyoS8TTH9yueGJRtCharDmxHmQe8TK57
V4hhO6JYXSmpC0yDUwaaH/dNae/qAzNeaPvAHQ1K8XL3hlXi1kxQw0W+6OlyxLUfNB91JudNRwU5
J0OjGcZJra6kVjP3rD/928ztkhB0QwfNKZl0amCSVKKzP1FEbEg/Y5zTPoYX7j1EKw1poFxpBrWm
p7U12e8ukoHa9JrgJlx3dWbQUQMfUoaDDND0UnfHHRnhtBOwTgNXkFHrKgp6T8ijrqomvSA4Xm4d
xo7knJAek7/XQ9MGysF4KhvKF4jvh8T2Y4xUw6c10ERwClR37FvG5W6y95mgGCMm2T+hqaq9+COX
dGKGB6YtyQVcso39wpweCgyDJQX7Fm82QMdAuA++SJuGYU8dbqewY/gKZKknBIMWYcljJ+E03PSY
vHx7cI9LKaRn4Vd+h9zJZYksOn6Hmc2Jt2IIwcq8Cb2ilyY/hcM+iDtFoZGG8Hu0LZTF7MjZfjpa
w39qUTi1KpqwWBV456Fq1NyFj3r+0v755PJHGVfuwaI0yddPMFU4/W/6tzNnVOchWrp3bONJNUQW
0F9z8j50MkgWKK0rAbGSEiMdCOBmt2mfvhAMvwYpzXg80TM+clsR/s8Ubod1iHDZ+e9iGxt1xWZ9
L67cmMipvib5pD1vmdrUTNgmpaqXlfDveDGJS8K08QXDjrcMrzQjWpui8W04On0ysblOVB+sHFaY
YCdDWRJtwOUZQ8yw2wGY5dW3RRnpwKfJKIkSNRgb9UaqCPbLCRXnI7foAM8INdDuDRC+y2C7X3G7
zL2wpAS0/KfmX9ndkbpQ0Dlw/HToD++eVjYvNcCaNwruZ6CTd3vXVvM9a11aIOVLt+YHMV28nCGu
Ai0dAFDwjNcCcmfl1ZZKlDYKFppZxS4GUVjBmrJxrOSiAM5njcQUxSR4RUhaTpKWjUC4DcUx4nnS
2fiUtJwLr9lkt+Wc5Z718yzK4+95ck1xAjS5mL9FvbDq3l25xRK3hOGpjSSc0QytkvXG1TmPi3OU
mO8OiUILrTDWSoyQzAOy10FyCx8f9CtBDS2teGqlmDmHh1mr3NUN0ouTOC6ZwQ5DkbYlmbbttgzF
V5DQRpEGMAeSlbeLXX6Cl+hv2mMf947AbbjcORfRCsCCvs7c1a0lj2i1Jo8E9VPargsq/1vb1Jzc
T3PPAU8dTWGugE1rCQrcU40cE9M1IlxlVM+JyRbGHFywh0q6JQVMMN7wZ2lqz/vMegQU/UCpdeZ8
xEMvL7urpAK2UWPFlZua7907JXvGLFdvJOgt0ZKB2OKTPHiXtsIIKmQMyO7eqdJRZPAXgNpT211i
i/u0YOVbHdqfSjPwjhqsGVk16J+3Ve6r176Tmv6U0bPLPxpTv9urcnFSlA3BhIHpkZJ3dhC5f52z
LOeyUlTGaTr56vnsOeWyYecgwh42rORnbBlrSjc/agzsxrZqDpettFF1dRz19pUjE7wstfUowTKN
TAG3PNMSMJY2dU/TzjE3MXa8b9YLYZHeCe8osQ2T00HJ452ne6y5BHn0mbjpSHB70w0XSFY1ovwr
HMN+DiQISY+EGUJkNP3lMwSw0QVGKQLx6XB0yDvBLv3fsBlJ/rSXJ7PvIDghigzOGCbnjQH5Q2Jw
QBMtFu29Z8fMVkz/XdnpBMqLhByzb0n1qKoeWSOcTWh9izrxwdLJHEPN85eWOfBeqmOJlMKnL5rK
O3hXEkqDVRiGSLCb9nHLP//LWL/0FQQ4/2im/ImTHpyp4x84uhEQQv59qQMBo9d19KvdpcCqe1tZ
7IzLG108SBB2/ZQ2IsgcQ2N86mwxUv6b6QkEFWg7HhsQcbBEOQ/njTldD2JxvmkusS4+fNdGKF3Z
P8HWDkQPHdc/4eQdg57VMO8WbTxkUhMNBou43h6aJQ8J8aDed0x6btXXkEEipBcyVkiGc+npKF4R
tZq58MCU/a3v9urOw1zH3iBEgqTjKlDMpHEVgwT9sJjLD841KrsDssM8oUsKEt5o6ARaCKqX+erY
nlDL9fipHKxQKEaTWm+0GeNC4wnP46zDCsUYN9goZn05MW5N3vFsw6dLT68FU6UhROaFCs9zfVbI
n+kRx59zrFBLUgwzsUK07ks1rCcACxRIRY2LxOwTVxRcRg0yflRaBc8l+ArQ+zdI6cr6/BhCdLTr
mdWhaYOFze/8CJXYqhOqTCHg75SnVujTyrh//VSn+WqJ91+ZQon5y36Q3eYpc/ylgzbnDePgy06G
TdgLDKszndAtFFL1dc5fFtZaSOis6JYB3iB1jSOqebK+azpOu7nr7QO2G3yw0VzvIeCv/Wu1KIPN
azmErX867JxHudrRESLpFwmcfG6Fx9rhE8yjtzGfMgLxaHcrP9M8jlas6CY74oitr823gmNELGcU
lbfCS0CLypbibNU2aEXcWYR3kliBlk3i1crxVtmoxON3RB/0HSZeVoKqV65j2WPc7X23TqUBgjhJ
jw4zw/RJcYMG3ZKXa3xQX5v0d3D35GYfku0bQhyVMPg5gvExjHMN8WVU6lzN7af3yeja0H7WPU6+
vLCLLLCInypM7sgHgfSYlY0iIZU4bHGV5hdGsMKpYUPJHC+yk8RsjiMTJzLdRUQ+uzWZQCDw+YRF
zix4zjfA6E8ZimAd1cQsq57c5ewk673BIR50j/AWjkgcb2sT1cBxiAj+DIqjpbpccilPjBRsDoE4
X9Gh9XQ9ht6wbGaRKI94fIG4NdjLstt6mVfcQDz5hv6jb78V9o9FPAm07RrVXHO8vydLmOVHAh8r
gif0FgKI7YbGb/+sZ6vuCevt5SMknF99HpT92dGByh10E0XqnHBXLjPpS6jrxiM/QVPpfCH8WfjK
T1FASA1LFO/5XLt7b4867HTWyfTFoUzYehJH/4CVVyxnisUBO3SMzvytsBXpOuYDms+21XUqpi46
wsmT5MxSv2hSYe5jP1RNbPQzQMSJHSte5TGjB+4qOx70Y7Bd5ZnSzbzyFep57AukAj28dQNlNFYH
vAZ0oTFeRCjsXF9KblrCLC2FVTYTMY/JKeHMt8ycZTESdMzh63DyhyD2uNfBKlV54lAL7Dwq5K6y
VfQK2puLjmu/fM66PiplAJ7H1+66b2TOz2N9rg8tHnqouLAqjpPoQBGcVqmquw5MoaJ6N6dFToYx
DZVzwOfIvzsmMKPVu+n7sAmpl2WKad9T1GQw2WWjv9mu3t+j+pxaR1ldkv03ItYFNqUGD0h7oM4G
RjSya17UDCJtqFmn+lJs08DpDuyd5+ohyasbbF6Utb4pS9KooxF6XmUzBj83SVS1LQz7Ljz0uw3o
HU5eDnBaHG45G0FcjvRmz44tQ0Embjh3/x54s0Bx0F+g32mDxwNSUz9P2mRRlHXV4PK9eqv9OkR9
LH+J+NSwdUFeHrri1u+c4LPbQF8h25xDZDjv/QuKsbdn1t9omglUKmYOTOh8y2cqw3gRiXnOhzXm
DkF1guVTFnDSxEpS2h7RfHYJBq3YnYWp1Y1uIpy5J7/n/P9ZYY6sj6O52qP1bX0x/f6cXYT+aoYU
ohwikF8jy/ZROla+E7JTLTzatLzn8u+/y92jpUdqS6RS6zaRLUyMjnV5N+0uD7hir5SM/yViUuiW
JktxoiD2r7Mh8iXB6EfFS92wvE325V3iw9hp/htJxH28iBlxCQkhAnQ6Z0fKYSJ4+g4tgo/MxPKD
+Fby9mv6hYcHmtd5sGosCIhWj7pyKiyT7mR+7/Bi1Gfg1I+TzzSYI4SPrl8uexRFZDRQ1B9/wTRv
p7o+L0AiYN1jX1eJbBYf4RpPg60aCkDDQkoPRnh/s716pD+MiA26yiInbjU7Pm5cMcstOl8mCNLB
WaGjwKEd4S7QwWRYMJs5LI+GhR9KfpNl13ywoVcWVsgVOpZ8LcTV2Ue6tbntbPUEb4ltZWjgvjb4
R0+tiJnninclMF2UDG+sV2d3q31B9s7mY/7fyQWzLniRgWobiaGVPzTzAdEHDXoUS1KaeCvDDsih
CUHMBD6rw1TZCaTsfM89EWlkbLu7e+n4VqqOD1ageboKyeUVPS2pgFZ4UI0R+0k2/Stndoih0Fql
zb7WocNAn40RVtTF07KBng9LDsl7X/pLOrbghQ0ONgXbxX+1cZKLr0Ob6qPDQrsic86xJy0132fG
B14kNU2/7gPlIYLGXBzzyiTCqW974CDyXiuojfXhiNCir0TeDT8AZdYVSujdMhLbhC4QxIR53cbS
v/4AkD8XiZ5UJ4vcEAYJFj0Pmwyql8gZ2WEHdHW7R4wvpCp319nHlesxWyfZTValG8jx1i329REK
gRUt1eJgkZ0fu9cG2O2qbVvmnErVddOWbHvmU+1kgubyDNY8qKLz65XYkKnqpMwmS+03Ni6XseGW
Yxw5QRkXUOXsl2Rrvz/Ix8HLhE+oiVRAXFE+SF6TqRkwLkRM4g+mXRp2I2iI/N7vBh8wEtJI50Nd
HANY9+0tUF50gEXYgSmukL/mPPlI63f3SRB9s/uNJ7d6wXUIEpi8LEbwnm1OlHmFnWytJFW/Zhkw
LvcJ3gu4zrhnJQ0/+Ubao5zIDxFEJCjnfnayuOdwEOfJv4YrlmI1lakXEad9wc15nAcs3bOeDhZt
1yGvQeitEFAEB/1jz2Kt/hL4wX5mhZ8GcAqx7s4i/okFd6QNlA9r6TO9gcw9JQRoi5b8AycZ8jei
gkK9e5DTm3t8CYX7GspafDZZcWmcN6VE6dn5NvqM3JzVfTZYdYHtS/V1H/NNeQKArRfWJna35xZG
kEqVGoVQTSnMOxVThXacwpsY+jZ0AFHaNRcwW/50wRKrjDZWehBoS5np0tNAABSpxxRCqQKkyZzf
a0OqIPNjG0nS4cbLWAyGygRlf/UdGhE8zMnFuH/K0GOqPV396FRiBU4Ke+bremqtT6CsmbfAGHF0
oWWqXFYYe9iTQuZAAWy9i9R+BBQQX6A9g5/IamfNhrYchgh4/MrfODQjOgHXLrPdZaEF2IF0t3gA
f98Ubb8EEPuxi41bFI9i9SjG40PEq3PiZk2I/ngWkDNZr7aP5MdL4DpweyfFAm4l16stN3KsNG97
rBXpV7fLMNSBtAMOXQqhW/WhfCWv0pvY8JLABnSmcU3I1W69r/u5ucZrBP3RqhRA8D4tztBC+4HA
mt5drtMzV3xsSjtIliryaSYCILPwIKghyVlN+D9Gb9g5Gn1rUh0PaaEGfS1/HKBOLbtBjLWheB8x
5DkwAnRkkTO8Xw9ADtdGpSiwrGBwXgZJeTG0tpBtBlI9cFhqVAVJF8vqH7P3C5vbu9OahqvTAA2R
UB9LMU0Dg8hhv8OnJVr+qHGJGb1USMPPnN8vmzGo5GJCWvBKrvTrMUjK+hs/k0soN/dCONoNzbmU
1mtbi25fFU5BxiF2VBv8/DmZcHRPZ1ixwtxPyzZ7k/ibes5JJnspX4wKxACiQi8fsPGKBdJxpBJF
xvlOR1zZcBAq49Jzim8ae1ZLVX78msC7ZA/1AetNz9CdPdDGaS58jlnNpi2wKrpq/X0gwtJOtsvo
0QFZVuRs/iOMvY2xNGd9fTAyeba1TgzOaxwDrvocyhILP2MQ7J08GAQlbspNBxCgL1SBJxdBVVWw
HHnAEAHNeO6sSQtx8/MUylUoS0lkO2CNJiXofRJXmjsSCaFFeZ1uk1o8OLAdsULZoUxIP0idJuOu
BruqEaBdiWLyHSrAnNHPxCQYDAZbsYQDdyE4a3Vd5nfImROLNvTPcbZDOW8cMv8TV9xBrjj0Kg0D
xU3XND4dD0/8GTQZ9XlqTDKbgx9uUYXtO5wv6WsY1M/NBRNAjx2IlXL+OSs51cM1uE4309qZWlL5
NZGkU3WDuJ0Le4+XfqNMaVYZaxdw0oClCyKa1nFlfuK/1CegNf7tPcHkqGi5hQ144dZOxu53ieTy
61H1KCMl5C6tQuA9ivU38HIO9Ive4NW5gzY3E+mZuLlO3+EOBtTysWqN8ve59F3AiV6iaLopv2nI
cVZN+me8JIneqE1pTq8Qgeud18BFhxTCfnT0L1s0Px4EbcD7LIu48ueLtClsZy9PAlxXDHK8RlYk
U+//gItlB/L2jEAEUXXQnYhRQj7NyExSM5HBVVPKOdtZqUijCdlnJsqya4XEwdAKoVj+UZ116N/z
y3450f+DoD2ewKyfxQ8S+kUaNgCWhj9uPezOmRTEDuXkmy7gxePL6XZpZ8K1rvBbyvII9Yllc4Yt
mN2tXsK5UVQrG5Oh7gXHVpGVy4TbNL47AYX2LJJEtCL2xNHJTiHN19LPz+0yR7mI8uTjXMGugqLb
7DRtae65nO3IthbIV+O4sChdAJWydvF6TEDZQMeAQp3/hPBKxgt4+XI5w3NVOnx8eE0uqXYMZenB
xoR1Oo5ITQ5Jx15ppCice3QLj9oOkdzTbcqAn2si6XWfF44sXW0VBYaAi3vUfgauGF2T+aIoAs5j
PXgD1ZXxKpST4fjYinSbHEUMGtEfO21QPMF5YRjpYg8Z+qODpAwv9aV7Ct0fwp6U/ofbyYFAY6tp
PEYzhS7keZECLuG8Jqfsm59Nl9IXuCc+CRIKviHZT0AEumnTdOYCqeGkX1/dL5w2/0NOVzRv3Iqh
rLx3A5dudbLtC9s7JSoEivsAVs3JFd0BylmXlsWbWTbmmTCul1L5vzuMa/jA56fwnDCasu2fKJca
vc3TchNIB3p4wSifBdK0oQ1y4fAW5/iIoha+dWwwsS69zkyyObeD89V2t38fC+J+cfrOhQV15gIV
ocLTunTh3QjoKwpMT+JRDjpPr2Gj77K3oGJcZGWacxaJGiL8WhxZSoewGzqv3guhUM8cbyVVgEQZ
ZUnS7EwxuVHyzWhepZ2VKeNRd3gCGz0vk2x8FSsnIkEJC/+dNHJgOusLtydzB+LuYcbx4cKkj8qi
KURy35WLS+uKB4N1M4hWzR8ijxRS54LlPP5Q+mMIcNC+ijmhup+TniPm3rJbwN/KyGYYskzSfj/D
w1TeQP90sNriA5YKqHKidwS47bC4a6LGMs6bBiASkFO8l0Cv4i7RRoM0qvtJyjo6dTLjTI/XFEep
4lfMKUtaVa3iPwpKPh0nqKjfBtwgU/w2jF5h0S+bng3yRCro0ydCotvejfqN7UXdyDz0gy22OXXB
zZimWZcXYZbvJsmaSG5OTpV4QVvccF0/U/ZS/+ZGEDDIm857GankWDV2nB4VQRyZnhsC8o9hveua
KiNcP9o0goqCqr24eaYGlZP64LU1LTE5u7jvSACCRXbXv8ROLDoLs3OXakYBhDxlCHJOXjMTYquC
OWVqNx98yQEAENYn0beeX35uuOVLm2xbepFLv6Ye/YxnbZ4K7Gz41hj4ffjS0dfB/b12xzoWNTis
fztfw+NIfI7AY+2mq7yb18DuxJghoR7d7WTqHKI1rp3CzJBKD295M1rY1qYhudVd2DDAMY0xJK2y
MEv/yiTa8x9kaOOP4nZbYNwLd0LzYQI9TILuYF8Hi93t1STk5X644AcFOvNE7/oYdJKrxpqrnZS2
OJdKjpugpC/5mmUl9Rp1pR4REMAwpro/F0kmG3jS/K0wOtzLQx4yo3nw9akTabVoTWmusR3tdhRo
MSGzCsquj7qD8wJngDv7SxsxVPVU0Dkfl9sftfzAVUqbsdun8lPvtjZVE5Ad27c1jEG6dujuU2TT
8/VpkB73NdQfQQYRZle40KTBLNRLHZpQrzvAK918lxO3irWMbFp9cJU8tryMqz8m7+/DViqd0P/X
8HI0EFCK/A5VwABEdQCRCm4JRH9PgHFyS2eMwAYU+Ybtd7yIRaZyyefkqs0UEdECq/cSeaBpAvrx
U1WtEG2lFiPA+xAg2qf9UowcbXPr9PiC0zEe9l07D50CbSDTjQw06gCLHG+9ozY++lOj+bq8qiKq
wGvdYg+/wHEe2srUNix4NrsSYPwgoT0kA1edpdwX46jWp1tiNOak8Anb4+N5DuNsMcBJwpoHLJUW
YsXha/BgRb6RC3LTBG29kAuQiW32FwG+DQQ6AtBXPVblT53BqHxCQ5DGBV7aNeQ9+M1d7PzT+7WB
NPQEx++c5V3+idDmoXMDLZULNfk55XUnOlktPxlF3VtkJzXTE5gXSrlX6jXO2WRXHUYk/KVaTNHc
wDfsAZSp+OcXyyenDeNB3y70UGldgd2plgpXl69yoMJlvQhzxI/VjV+OJ17bma54wlviyywZWaYI
Zd2vgKqIFT1z0pyS2CmSrokxXG2i383rfd9gW0ScagxPBNcnWdfztE1320k6TScBY2QzM4ly2//v
eytvZ+J9rQ4XOLanIGSzGpbN0ucnJdmPTbUJxXQQAoOLWqAmthfwjg+Skdz/gA1wfg086hQfFeam
tFWLlsENLWVUmqkEYps2FyL9ChKsUIZ0ZLkHzZVN94cp4drbDKwFgvpRYVC1kge/ohlLj2Qdwqxb
vwVJXHFqRaYGTEbxZyeLNwq727GAxXTxgjN5V37SWT60c1ANxEwlN7PFjiGVvjL53gxzDIvvdsdE
RUB/Jr5V7lshhDdMcl9I2BWwXas2Wckosi7m8G3IzkJ9UVJpagtVFVDmP00ZUdSXaJkeZBoLcJ81
ioKIigxAPu0oYruXC9wckzNjd4L8G7MrOWMiKOPKtQ76+d9Tl7K3jlCYNkFxWjszxuqZeFT58UKl
Mnu8+q0yyp/jOQsLA0jsF0zOWoLG7jH0Utq6cTXerEf9fRBcpnw8mvIxDd0BDe4AvN18o6Y2A5ZC
lcV7xBcMik/DSk+UApvUybT4hE4jn74eysQKh1VqqcxWYWwQ1YaP5r/JEJTIg4AD63U9HnZH3VkX
aNHxMNYOCv8HfXa7TPgQSv5OxYs8d9CIqmGznQLJs7loEtNa/tcizKTmjKXfMKMhFM930PEF88Vh
LGyCLecbuDv6BK4VB9O+bs82ZGhZAcOT2eNfk5tEFhmeQHfPZp7139zKc/gm+ENzICi4HAWLHr0E
yLlf05xcJrEEDqLxxYJpeEba2jPi3+MZFRk2XNjuBivEVEbcjRur4l7pdmFB8jx0uUpvzYdU+3HE
j4eHBmxtDgMug/qWCs6pWBzHLhB2sFHFdS7w5HjZsL36OdRv86chR4XiGzCIw81PCrIj6MwiN9td
j8QQRHfl+1YrqIB4PqJqrC2QmUVKfLkX6gH777CwfrieN8niNNmti33ibvXBX0/eaeThMzJuyhZ8
URf3a2Jh5aE/8I/A7HozX6EJd6c0Z5S2hNnBeSgrlLTSIDcXD15xIn/l9FY07WP/3zXEJ+5NnPm9
Jiufw18Y3I6X7IoYShSy8bG/zeM0kkhoHIS1PknCO/cO/erIDr0mBHhDg+ghat1xptyqExwzYex6
t4SUu3GQSqP3rA7nXXql2owC9QWV5KxpMnbm2f4+jTPtF3JyfZIS0RDbDRMnyiCBUo/9Cghcrj4c
fCb+ik004U17MLba2ZGFAHVro51kz5iinwiEnRfmGSmc94hQJQtSchNjxGi3UangHcpPen6sm6HB
OHuYqEi/RCZv4dYArKee+pEZNaD3uH2YfHu07tIxYfaryuAoWOqvasXhdG0N8iGOFvZiwUgApbFw
6epQ2XmocS3ogqyzV3lQkxVB4za1izwi96pzsT1hLd/5/HOu4R+k/G67RSnuSTqloDgl+YH9g9uN
i8IXL1zjIyvg/zjrdGn5ERVIOMyIY1G5xEH9WTP15caUaRU/3J00TU5bUJbckHPnW+6Q+ljQrKx4
Mvtwre2C+qUQkth+4k66661HFUBAzzU3AvhPOmeL31+Rgk9TXslH1vpIAKuShNuvNlPJSofazIrK
1cUUqSU94fupLnA4qLF7B1t4nxEI3spuxdthmt1co4Wgz02cCjbgi5TJQ3hRVAg64qKLnCrTikz7
RckP+AEuUgCi52LpPfMlLscUIHj6cS4kp92Au9Zr+b2VNxnRhXYmt6L39vrBbDV55FvPBkPswCXj
KVsaJvwbSKM+UmpXiZCK+O8P1qjU/DDFW46wDlYTQ/NTl+p03I4gu/XZZN9UpA9LBg7jGGLrUEAw
LAEyH1RmAClU83G1Xpr1sKat3S0oZlmmPVmbFMMdrO+GlZp9e/1Dq/GdRrhJZUij2slIgkILUaqh
YeaeW2FtxAgYjCcbW/4onvKR8DK7OVpAKJW0ry9/FUh6Viurb+f0WegIixN9r0LsI9xqkBJtgAk1
kNJAAh97VOmBJSHwk8TBQ+VmEtyBVdDfKo3Ud1tUDMFvBuVtfG8jlDyDdMzfzeV/tJSyqPP92FG2
v5/S86f3vmdegej53njI2pA0DE0+tyVFsaIOkseIvPWARrhnI/VwE8COoELkHQFf9yiQKWg2otMA
XbJi0JasypQ6XJD28R0e0dXeX0LolET/1o3VuwKHvzUU7MDLuS47qXr8mkpyyJ1vPKrX/pS/AgQ/
h/GVtDGu2iGZ4SrQfpp7NaH14PsXhyvZ5/sm83va36sVhY1qvMrz9vw93SNv8/vCpCFa5Qt7AXOJ
t6PBzw+bW1mpXXomlci3/zuMt7fUlHI9+WaO0uQj8o6FGi31BPUvTqoNkrXeyE9CRgqpdCr1a33/
QIYbmEJtdSnIIfH/L7nM78Trx+3aq3wYrN5SGgPYPmmUiPPEbGIDcck6dVLhB/pdRwsvRI6rksP3
i54M86tf+Ll2qIzE0FlE2CJSOP8WJiLsR5IlZt+ZQUoN7UpkRJ8/ue5fOwLWEuLGM7V7+ElWE2Hk
54w0lxU0boFUVndIDqgCKuRPi1nNJnT+eL5KfkmohdLRzYN2tCyHuo4nG8SdrGkLRn/P108pZuP9
ntLugbxL/dOH/EPzxyDuTnhb6Vvkc/tf7WI4rSODrD9voE4i5cVRE19VdtQtSpt3PuFB0d2KPK1T
2fx5GK08Aplk7BjzDTxgJvKFSIK4dA0fzob/81t1CdjZliGpMuyX4XGpV85RGsIaII/CdYgo9E1H
LbKoYtHXTiKDG4kJa4eeMkyOox8ddbOqpQuF5CPymmDTukXoiVFNbtybhO9d4G3/mVD89dzuSFTz
MPTrLn5+xvMSXJQkEVCLx3gjMON89CGvXAWnNfquX4/IoPw/QUsphVVpMvaXD9L6Tclv0WxbF9LR
MfZLZ/zuib6dh4Yq+voBMVxK/ucW7e6PveHnIApGVr0/80VrgPQTkzSDN8gTlipw7yMf0ltObPxX
3IWrh38Kxt/jZpysH5OIHVPVAP0HpkQiQOrQOes5HcN8FZ7sGbRKaulf1Z84QqgxERhOTgbuKOsD
gSFSAWXjM+4t43ydfoXXW9Wdn4A2/HgdI1heGJ3cdRvnZPWGv4f58B01blAzZJopUPHA+l5PhqKg
GpZoFMIW/7rtnoOyNtx1BxK5gaAVk0UZ9hIy6+QZ6EMAmiVOiBqEMb2lpZS+d+mAVbn/p2EhFqR6
mD78Os3C6IXns1hEVJOmigc1pTJBtpkVrsk6bQWr9QELGhPLAxLQncbZs0Wih1sO59LqGB4Q16Rb
TsFyLajL5Db87pN1o7Icrc26tVYpaXMM6s9cBkkVdcIZBJ2mZEmvC66JCe+EINibpyxB2nrqEQ0W
Lg+oarM+jSaaPt/18rKfunBsOyLpCOgdHwU9YXVzwalCXEVHuC1mNO/ZRayLTRtPn9UYW2sXS2x5
EAp5dQUEo4Dh0uwMuebfv+yuAb8OAG0PIsM/d19hoXaRdWGZJ6nuy8BcvwangLl8EYS1lHCFpKc6
2KRC3tYrv58H3zR+a+kDwfD5duSTjXTFHWpjAOqE4TMos76gNHDInd9AIP7t7SpR1K82O6D2vn09
BD0pNOJCR75Ep59YcYMAyX9DY0yEnUK6XIDgNqF3X2SFtfXLHZ75JF6S5rsa8glPBUQhGiHgQCUy
shQ+XODPvdQUIOlr5qxtdIsFGtrjPeb3WRpbpWWcZVEP3thjLZ2koEUQAi208cv66WTuq7gvolZS
qsCgJDuVhaW/KWrzxE7WDe9wVnGS8qdxio/o4KD6legOFQ+CtVutEvseag8xsFjHMA8z/5gTwF5Z
y6cSMyY16c8s5QLxW64cXpDjMK77meda0svJ97S1kQpdKH3CSxgy32KXaWsZoXe3bRUQvqmVYVXn
o0JAL57T/46iZQqdsCEC5ZNNvDabbKRcDxcm3hYMpoXM4S+HRlqJ6E+4gvnbIYfrt0EUYtI84pcG
01IddI2wmZborK+K+pXldWL21Q+FgFxm5M1/qzEia4zKTY/2KP+HkX6oNqIxd6vcnGM9I7ACuUH8
e2k2DmuR3YLHxxMJnLwM5bcv5IIrupcalCpnYaDiOwzrN3482W4EK0VpIuXWCWVOJEF2RnSwE5Xw
LpUBSH9Nycl52xWjPdVTL5OWclJW4jjZDZrq3jn0+0L/GX0brWCQ0wCvECgKDmpGkbpXMGxhArP0
BCDq2BzOdV8BAziqPJmqBbfWAcjYqXuN6RPdPaV/mB4w8P2UCf8yrhwtQcRDeg9OOCthclzbKsvu
1CAYSvfXH+jUiyG7ybuXE6PXAyH1TgF/zA/vy0R+5M30JMi5LM56SVHaEgul/FC6y7JP7fEYViuX
mDzGgB+FzQZ6Ap0M0K0icMUC6Uz7hwOGnnJRjT9jenhSRDm9oitziA65BO/9N9OK8yyIMc1Jnna3
qPR9bJBY1DppXlYNoG0kqgz/g5iSqoK+ZHemdsbbcJ4EIAXIuoAo6N4XV9Qe6wW0GdBCx2KKzlQD
Mx9f2BlmgQGIaHlSkP75UsaRI14PbWp+QK/HXF4CMRNdyUuewwmm81zfHvlMjcP5N/6GqU3TeuKK
XnaR6m4fYheJut9KbfWL63Wuyoi33FixFop93TgjV3zHRLPEWyJ/NZAXTndPDmZXxisT9TWN5bVc
WLpupzH+BAyr1U++E1MrFCqZt6uclLSAF2ErASPvC1fZ4Vt4gQ0No+5Vf5r6iMW6ZwL8NOBWrE+g
09xCRUmni3g6kJagvcWQPKP2f/9qu4ZuBOED7M0chl79rUQ7rO5yH7yE5HzUUJYBZ2G6+FWgqpFM
5yjzvPf0I7a/JEmx2l6eeal1AfQCglWvLprvLW7mLCAAWLJZYNCJ6RnGu1aPJTjrV6AWJAB7VdWM
ftwZquS9wxXwlyl8ah26KXigwH/ilmlM6Q2ZCj64vRI55uvFInZN8GIqbPaywhktbNEOFCt2eMMI
9EKrBIv4j2pw4+fWCEG+Vn/Au7CgKuR/FzNHWbXaLGuV9XEN6nyxU7MaXlDBN3qw8v1TFxZMsStX
SNEIM6tyKoKermUxtAyJbpToh6ZvHbYFCxKUWsURwDiXhB2p5CMUGoDGzDxOHxHHiC9NNwX2Y4JR
IJebUoUK/1tVmZuDxwYBdnWX+EkUZFkGKSJjTFDcwheWJ3DOVJ+gxYvh7OAhwb+uFSKyr2j9sdhq
feuMfmjMk6jxjmn/OHTwimyJYdOeqtDjaVopsJIsiyjlw4T0BtRRWEElJYSHmulEfHHjxQQ+o8t4
TKNcGhuZizjz3nRGSSpb2uXuZK9XoCF3W9DfvOyaBvow1ArqpBP7MD8e6q6ftbmQ5jjDyBa98PfR
yuCGVHYFyJbCDV5r/uA5em1uGbhe8PX8VwodzWnkDSvXja53xW3VMJ3GTFxHJLoPp3EUGe88NwE5
XzwJDDMyxcfpgdixUwj91tl0StTW3fqUSXon5Gy7QZKWcJRFf9bQvZTtMPyrn0wFHCbFznd5JqZw
myFwIhos7+oEWv3arTThoYxlE66GWlcQIcjNY3LRbwg5A8AWhD05G5uUGlxSXx6QZTXrOYCRGEgz
n0z0Om1WQ6HsnQCwc1p5kTNCCmnK3tUUBvOegWSz04HVlrJaO0NLh3qSJYqCSAMs6VC9kn9ksJ65
pPJQ5UahgcD0CoTCd9bG8/2j3GY2/O8ufg9dKUAkZ8r5bhkFYXNzX1X1oVaoupLHHRiJKv06/5pJ
qaaQSKW6bT60JW89yWww9PmbLVkuSb1lfq7cc9dOmTL5MuXJlx8l75SkEMb9yDMO/VHRPa0+5Djs
bpG5S2gmJUdoG206AetqIcOOVAjEDV9BgTKFpLLAuRkH8F8c6ohxrKaH+PsRsZujfKMqNj0zBi+n
lfWrOQhXAchkKYS7acnAIrGneu6l6YzPitRxyqp++6tvswzP1zJBiMZjfGR7YN5NdmGL8J9XNNon
gtSzZC4hKYaOJGk0iMppiWzUe0BeW13Xpv9p6H5TXmMItTCFZjMZ/ALSEZVF3FvvJA86qaVYbdlR
RqSlLX6OAYhTwKCKiBxCEL8YQnXJssx827nNbXjqkSVwYRfMYS2rzFODqXf8K4X1g7hnNosPoXWx
jmlEeFMP5oMPsURi+3dzQ3bWwnC1/wob5R43wiDCzcKNa+PxHuXN2vtYW5TyRrlrRUjIiHJARQG9
Z6fVELJSzi6sXON8QQD98ZLeTa1H5ruCzVPWqxuIqdpRBHfEeJB5aWPN/Olb0adAP4MxO2TSxsMd
K/YObeq8zw3WfpFUrC+L3LUzqQtokIt3xbCQgT7f9oV4lq41xlb0DEhghwY7DrfNm2ZvpEAxHOuM
keynlGLgzXkbAbLhNRJZIYPYkhv2N+U9epvklz7vDXBWvJQxzOslOqWGKkjxBDP7XR088sZ6Qayl
s81NBfjeI8Vt9CPwN4TxROvpBl/twLq/3hQGteZqR1lQXNVAPtVMlzQc6Q4XrC0S5pSNrN4OMOEG
aQKlLBq31VZokgWPon4/SUaOTmwk3LNF8JO1hixZA1HNuv9iHUM9VaOALljQIPxOE3mZqV6XwmLV
R1vsJbr/6h/0rtk17Oo8chRvCAip5yEbTQp8LfpIjfBZ6qbeDJFuCG2dknqbds0m5dQXOuZXNoPQ
e7xpa7s2FXB2R9JoYNhAZv4fX7E9BwdPiURHtvzP3QUYpMulGtjiezZbRaTZbOU0+mznnN4txYIX
2fL1brCj7Vd0hRVQ6dA1y5zKedTKD/Mf0X2PbFGKjqDXrJrGQ++Je2yT85P1DZbyPI3QK6lyPh/S
CrT0Suf1K9/sFrsijRYzvw1m8nQir8UhOyvidw21SQ8gjKvqbwGOsepWNJpfzG4fG9oYJCUExZ+o
yFjwURiQm1g3j9gutkVqTa9eVJhPXID383GN7RtHC8hY/+f2kCUvy7IgEvwCbX4pwfGrqiBDr0rI
fFUGlkADgaxDrLJUlP0v6kXMLSlc5YvtOXsSbShunKFp4xlFwjY0gQ3Z7StmI/sOnEkLpyindXgy
FkLnPvDqgTUnngkFpYdhWKUWFS2VsJ7gOtJVJri4fZpIEnFMIp8hDmpRrhf7KEdV8MWNtV4YhcP4
bHqf60nwRK1ss47DA6w5BEsvYHVBmID+wczw6lj6tW7cidfS3f6bEyYgNweMUO5aUZ6vazG8KHld
4WaWU9vTV+e0LVJADfJcaKWYK/13XHBCuCtVb85x23z/fIjSFckgQvuJCe0VHJiCC7PaAgOFZHzP
9jUetrbhVbymxtM0YatVUguGDN3QsLOtXX/JhtTuCP/murpn9awpPMMV+Yvgipp5cZkIsc6/dycg
XXL3uHOwwTNRr3a16FWi4UPIv/qPaZbe3nv2Yl2GIQYHICaPrrWP2FOTlIu8ovPNW2kYszZir4E9
N4Ezw7zMXUqYL22JCkYDSjiHPnrh/O4qzqh6pYyfS6pNTfWh/XCW6fBh6Y4Mc2zuy42m56iE/Ad3
nt+7+1hm9P9DnI7mUrV8VeogBSzzpkt+MJJnSCc0xVqW1Sb297NK4p0NXaiUtTtKexu9w7aqXVbN
7+uICZZw8EtxIKfmH1wfUDBx1KN3kSTgA2zT2vCGnssPUtqQ04uAyBHdYmTFnPlD5JscJiVpp3Nl
COHac8EENVrk5G+pVwd0gyOi365PbG6nxEUFZOQWqS5g/Ns+oZQMKiBjzS0D2oAtIkexmUmMmQiu
ySiWPxYZwpCg7MVU957Jjkv6S5kc9qq5mLe4tg4nd5nw+TMVtMClbNMYddAe/v9MCTaKOaMc2WxH
vEy0v0bItuLeGoGQkITUjFohy5cK2UfAeZvJwyYmvu8neFv1QlVUjuXfFv51QbclC98GosTZ2bkD
nNeeIRwzrQFRz9oQnFIWx9Mp54ca4hpWqJm/cELti11gWJlytv8UIS9Gk0duS2SZB02l3ZpZK2dw
K3XgmDyLUqv0l6afM4NJ15ulXcabjXM4y+ocpodBoVPPwW5r/evUbmK31VMBZE7NYovfi/A8IHaB
cqXn5+J1RVBtituNMAvGcePg1i5evtrjwcu3i+54cCkRxmtmv9A7s1WNZsFszukTymiz2dp4kiAG
BT4PSoZ8bcpXi50tUbisQN0uV4AXpVolUo33KTy7ogAXwKPD1b178UTycMU1LI9RU2J6Ci0Q175p
Bcj/u1nOZ4SB3HB7NyuxvBVVwrXgjG+MQUWSILQo9ShCtgudA2wdGTY/g9nPLVQL5S8l0/bKjHa9
cV+5i+bfEpvmPh0mcjQT8LoaKvlba0E/kt4lD6CyjtrmolsXUkLi550VRsy3g8PcvlkScblDvv2i
0Pu0APWs0EfjAY6c2TtPkMBWhinBfiAPr95+FKOCCchxWaXrZuA6oc1wVE4s1OBW0uXwQpp5/wcc
I1sBWGRduutGT4BpIiIWbwTxZ+R06nenG2X4iRjcFNjgRpz/zvYXh0WfCO7KjVrDa1OrurtJPC4N
4IFYHCdTkSPg1dbIbXLge9SMRk+7Tw7iTD4XwmEJkwFNeSkANoUeFQUv9A/Ic5fh1AIJ6Q25D+Oh
CPnR56A43J1BSOdVeFWJr6Wqh4JLdXO9FEeqwxWkrWJal90pmDZiPdNVNbmhdzYkTekKLtBhJu2o
+subxi+ZVACqFaXaT65qB5rpC7iahSslw0RlBUAR+Rmpbq9M/Or/UzTxHJj/W2R6bmmu9HqZfI+/
9mRQyXfRmntxaYaBbeXlS7B6su3QySJ+IyrOjZB3y5Ljc1uopbEecmAsT74oE78q6m9e4SWJm38j
0HTECRKgSxFIDJKre2J0UtViNBHWr/NPaqxeh2WxTTS3nsOsmIi6EgAhZScP76cXgAZ7WsPIRm/3
fnMuHB7xjeF6dlviIkt9tATuTX8/hQ8TV1X1RmliFYNvVGTMQnB7yfdiXv2l42dodeGX5Hox8apL
um/SOO9FEsWqOekjSUkUyiM79Rl9RfYo2OgtL5gGMZiOcWZqUsvf/ogYEjqwszGCLSKw8Xp8B1nh
R0xRlENpNdFu/o1lmUTMKziSisNdt8R+PispOInp5T0/UXbbM9pPSniHFNg+biCYq8HzA4BqSwFA
42xHTMYGCLeI1MRKXv/bNXMlcRAHU6RvomSeMmYRTFPhJ54TROZsppTw5EtFG4yUbkTKpzjmw92H
IS787Oe+iCev2ZSZEgXhE/7ZZzKFVu1eURdPbDRnqu9Yl9hqyiwGZBHUrgYYeNzL8+iVTbHpFabK
kFLtB9Nnkisvz7vtP1CcuVPcAzp1tCD/2wlz9YLDPBzR0Ja0LaJxSLlLECUb3Q6D7tw0wp4ewrGG
kVRSseiKJ6hZOxDvw13jMuItyyennjyXqGbY3yAzSI4THVrJpGnuA1KoWJ//hLTQwcelxlyYM1h2
UzywTvz7PU2D/kecs7g815XCtMY6I351EQb+6PRi79S+tKEOsPoJXjo5ftLZMwzhgxyXk5mLWpBL
pIDMQcSVGCGRTPN8MvSZSZ6qhQmmNAEc6rpnWg3l+WYUmF5WegnWyjw/JZ7qSDAWKQpAIGIMUFoF
RKM84BkHt6/JnQ0006Wf7MYs8uOubxuo1dmalX6k/ww2P6iT91zfGQOVkbSK4LckBk9tgsRKzxLa
IQNWpUTKQIV9V6eQFTdT9+0WgGLQH4+toC5SZmM21FAjjPb5MbrPNrixd4dryzrXXT7++ZTaaGMe
lJaFk8P3qXJmiG3ENgNFF3cvKE+ATnsZrCAsfVhr9zccKOLsFLTUSQbYobJiBfdJBbney7lwmcdX
wGRhze4ERh/VCmKaIm8mKbTNFg+HXCMhV9Bw/6lprcXu6ebZJGroRPMajdr7ZeQdYH8ZR8DMIdGi
RoKxN1HO4m9RNSNtWeGr6l2/CqF1tpDX5x3eTUiQXqcAC/iT3ROOPh83vxahG09u5D2l+LCplHwR
KeRv/U09MrQ3uw16N6uLuLdVRHrkvOv7e5PXFNL98pEEGulY+u2ifCZzTJbht/8FRMpRNkjuL2HZ
vsqUBb3YthpMZDvkuyDfSYtvdomVukfQpwiMq7W4dzeS5PSfQvLcq9lQ8Yq58pWbQ2Px+L1O1gVa
pfmc4Z3DhiLhkVbdxG4c4DqXYIMhKBWkFLArRpNbYE8Sokh/jMHqZTWmO4bAhbxkeRVkgILnIS3t
9uPmmBYsGShGdxTR9BrtA+9riMuz5XZMdIEXudfmvjjp1zn7Fvc3MK8WBcqXpbv2s81/KxWLkjdK
nS+vZ77ODbk15bsTZtBxjU8LZrGPOAGbi8QEfTwytrrBwrqHVU+v8qVfKACyhdueihU3MUFqz9r7
Tn/MvqLObKCM3HNT+qZWlDfCakXxo/u3UvmhQDp87mxURmxhZFH4Oxs92eI2edIxxD/kcY1cLxtS
fPLOfhUL2A6GIa5fFZuJ7srpTDqZvw+Xas7aQuuWffR0psvDwhDPKrL/Va6FpBGtzHxNKl2hRAYK
5PIZ77a9E6B2EkZ0QDcYb0ocnCD+BYFpUtPaWeJbu7DG4pgua5tkbnOqgztk8VH+ZodpXd6vCPKo
EVY1a8qjAY7ZfGj9Ks9qrG8ehpq+69P18S/YWOFIp/TXs3kHOLDkpiBgGLY3XLIRXdAiq87JF6Bx
ULwq9nIcUPdtVlMqw041n/R4pPlC+dc8CBq8NWaHGMwpd/VjXVzV9aS9tWZ9gOsLmBg3qm+jpyRU
8fdZMKVVzJF75T4BwsGWtH/fjM3ZDAykzWLEfvXkSpekUw4GrHbKG3d6mu7nsD7advyu3er6S4N/
SYZ2OSeAm1gjatpH2ozhTHq8C3Mp2MMkhbf7fs3sYaXx9HVtdembFb3ouMtE3svbuyTNUdus6rb5
LGwnx1THR7o8hcZgJKSP5rlKRDaIBjmlqn90fKw8RoSKcR0GpeCTzdfTtgXY3xP9AVQveIhrwDI7
WAdj4Q/M9tErLU2Ck6ZkpT47ZCjPZUEzs/VABDvnVuK90tP/gfQU8n9VwzvupjHnEm+nsLZ4TZht
8XaUfE7DV8ftssbIQ0LFl/VVoGKgVa0XiLUrr+DlrAjXaFzekIwRf1oDr3DNoKx6Ql03o5fNWBd9
E1iaf9iDLvI5QV13VeWk97W5eLscXFiAqqITfuyIvpuDr6qSwKT+2O8SGGAthYDVEG5eKUlNAXhs
0qyWgQDlczVHHibgO1nH7FzhCQG4GFR/svCP7A9+6PA/5HG2wE7SfgdVhTDHSRKVKVmYJ/0pFd7p
53MM35KeWSsOMW21JMFpL5g8MjSvxVXGvHbGp+WHHprVSEwMOWj5koBgyxHtVdz6YO3j57E2n4xe
C/ZVa7eREpzWQV1ts7P3Cdyxu3Zxxvcy4KJHlgBC63fvoReB6ywcgWJBuqA/0vgd9cypZ7SgWQdi
ojV82R2sI7gV4PEm4FWYW+SzRDcijeFmNskXX3RvLQ8GkIQxVNTYB/lADgqZZounn2A9DUXTJKX3
lMoAoWQoHIt+gXMmLHvuJEa8u6j4yUbgry0kauciCNje1c8FkCzZqYQicoua5CRDeQwG4d7MRt34
EX/l25kBMkuTbgaBziszuny9Nfp8E5PWsgs7T+QXwNeIklnJMD1a2PEow8YX6Qj29STS/YYU4Tl+
vXQe23g3Ka/mqJMUNtRZjTL7cNkKxY38f6qPnRuVlCi+2CXMn83HlkKuuSsrYiR5MwHpFgvxiCqO
NkQw7YyEyJbBZqhf4KS7L77GMUuReXsqmfLLlwbC3C08DS1QSHENhCiotxu2G9BEsO9ouGLV8bmb
M2itS9Edy4wMxTvyl+U0d6YMTvj21oJjqncawRc8IhXwqgTHkO7omO7J226nn82zLCwhlOZYR/9j
G5zsrvUekyy4/a82B3r/IFh+Qehb4Ch/gHsyBOiveWKfz8BcRT7vZCP/5NAmKjgwiBodWwtympGA
ri8iFh68EDEOn8BbKJqz2dcrJHZGYfvFhbHutb+5RTbpfD9fFh60sghAG9ZfGznLwnHxeJw59HBJ
LbFShHLG+K29kyqwXoVdrV/8pxFTzxJIiLnFqd/ntVNDzpFEtlS/ymuZCn3ruh4GBssooXAPCrKE
tsORPJfikcZwLB6MwXVAkJzKJoonQ01uoVqNDUdG6ieLz1QFJQ+hkDDU7Z3RaR0xOvdVC8t9VXMc
9mNAUR96aUd4S4FY3oVACgw/4z0+wLL26HY1jbIprwddyuZQ23lWlvwbJFTHoWuFrO24mkGSAUKC
3cbuq9E3ncRHWLu1PheVkIhoObp2WEbbQxAmdyODqLiAMk2E9mFxSsc+00f1X1sFDoOaD+SecNIo
Lo/RzXrIqHY/DHAdId9BSe/jxy3LsDOMR+KkGlqJDRiLQbLQkeARKHuch2yJzGVmv5HuwrZhbjfy
qJhFvLmihWVHLU7AoGCLtqjG7sqsjqBtwsdTubFPOgHw73HXKOXA/D46wPloNtAgdYRgLiSmqRlO
AuPj4kEElA3Qo60loXDgGmqztqfVokvx90t81P1c+d62istKoiVb9j4u6yx6qXp2cQq5uOFg9OMu
bgw63Jq2tvTiAjT8YHnNJjaeUnFVv8HNpQdtRGDzKc2cQPOxYCpYyX5GFOJtoa3aGJ3WKpKeYRnf
cyPaLL86LTouq3WFqKSRHFKv2BIzy7+7bGeMmKSFjZZjsrrDV5MLbnvVw3kFqtwsxFaEyJaKJgY2
zuiyJmRyA2hi9AxHw3NZalBXd/zjUGzy6rE/kdjmFSTdfyY0XvmNimXKBcYIBZtV0nbsCqGWOUz6
RbmIisEaPAkQzQRVhgicPj6zna5TYS1y4lthKpCVKJu39IDnj1AN+7YiIfiyBdf3zvlpx5taZAzo
QhQUjHt1WBLA0QspFOt9TagyiiizH1Xb2Kp0C3uOPVaU12v4iTITNUTBLNI1MXxHmx3v/d+TkXR9
DFFLcgRVld0iKYma84EUxz//lONVsY3bh4hTF+D4j3nUhUqSBdGqg7/OQRXotnTEZ0U2pt29rar7
/QYnbhgQzOKzo7lsoNnkmcgITXbveGieYLpMJrguFMolcZubNkXcK0gR4/CsnwfUFcmCmxaYAyAR
c14cCz5YdrUxfEDJMrwl7WaXg/ixIpRQN7920VLPalhtYsOM4P+1E1JAz3houhm/VZQ2yedu5AgC
6KCqPVZlJPZ38BYQojMcsIkOMd24+q2i6ssX5mAdOGaGR1+XV4eylGEOLXynYwaA6nShzZPJWHr1
wgu18z9EITgdnTNgzTUwG3TTqm9XORF+Hr31NkVqwn/jN3edtGVVeQhT9TuwKH7XUcV/0dmN6j5Z
ampWkvarjBv54zQ/gY2XeUlzj8eriwsGNtA0xXcAcv8moFFPY+vh4waGM+/gWmP434bXjjj5COum
EZGRkSWFOkBjF4g5V9q4CzDCaYjvPUbW0VOWK6a2ag5htu0BQIX8N9o4us5dr0SRoQ/2HV7iklQx
pCMuLjD3Q/vtAwElWPIbfziLGjsDUoQLaNGuS8ipm3yfaMU4TMacCEWnZXrvh86Z9u8Xb+ZY6F3w
le9mcc3sHB6VNCj54Lj619eGIeNVQ9Y5TPB4UXl45rJbemsBC+yWAwa8NgeuCi1V9Q2fY7NwiSG0
xVabOJsSBSIOg4r3uPR+JlhjkQ5pKDOjQOIWallo0pU40JeYLOmoYfEOzz0tQjmdaWJW7WTt2VYC
Mi9DNyWowhFny5ki/hpixYpwpq5z0BRmIbp5Bq8cnIR2tRvVzibW3KjVcEIrX2hobUA9B2fXY3PV
mEwjPKYQYnqe9nG5wLLfD/wR4phs1T2erQTA/b0qUHsyGb1a7KCW78/gBEEUEJqb4UhOZJlL36bg
4XmlkbExk7f+zftpR0cYfqJUsnDNuticitIpskDXtALruduLMy2d6m822fcy069R+adwXmn48S+F
imoDKR12hQ+KQ7KdC0N6KTa+Bidwta7LMr8oKqco38jgJqJgN3jSRWc9eMKx9gGW85oVVikLRKlF
K1/X+fw0Csoac4vjln6nY0vBeQvP+hDZ3uGAfq4zcTSVqQajpq1h3rQnIDKqr4dp9eCcjUGUFxYv
nqhbgamRra1RjacaumYxcGWTRnIISeZntfOYe6F02YZivB9uYq8Bv70s4cf+Am902IWyIHxkPwyL
6Ndyqo44YgI1c0zcPS5mN6onUv6tu7LheZEH5aYno0zInJUngWP+gPM/XzQBrSpBB3kYRFsuS5Ep
hT/kEpC0iJM7Rby1B7IFyWEWF37nz48oWMFJkSJNFu4Q4NzwbtJ2kfmjmqfYlo3wh1ie6eiTMeBL
Tz5HHzI80oQ+HOK+8rzB4h9/vH3xunfxBHbZoNFWhc43fCA1+mu2G/UXf1CmgZQypMExKi7cu+JZ
i1SjU9ZTuB8hRZ7Dbc3pxBkUUsg2kp3oLCzYks1DMjx9QCBmFMyJIpwGem9oR0bXManvNSzJgAQV
liFM2Gdbdbh8exWwtdzOlLjIcwZeYLFg3woyjaw3FFsGqQwqCJMM+5rxmI6E6SBCRHvEWkLQT+BU
lPXmRvkgg558baxkw1NOa/8MhnHDSYCrhOckt/xmKWoAuWySv2HltNMsz1SA8bp6NOsQw7KrxYCI
cNtYAyQaOjrcDmTY5SRVozjtq/+EZ1ycGRMPZdx/9ppJDGb92owLkdeZsgmrjoOOkpVcoAkCHMrT
laE+2budPLjX2FFcSoJ7XuQOsaEhzXB4la/QVQs3+m00aKXyPvUbcmyaXwljOBFjk7fNvVcGTd95
80ri5DWByxPR6XnN//vEKsbkQUsKhWiqA9Tb5i8yhfUQDKtxStScxPvxvFkx1DhlthF+owUSCdeC
XTstme1v8j58RIebVUcTaTlfTJODJGJirXeFfxhaNz7nlpwKD8Q8o+WtFQwlFLpBhJ8ga+hYw5Mk
SMP/dO/qjRhX/Hd9czBtBbf/6XPVoCTL+aNwSSVyuaRpGmk6Y03frTxQi+fxRv1PAreu6E10Kzo5
OzyYyggFGyr7XsNaetnZ/IV+OYnWhZrU1u1K8CSZzmxKAqb4719HDWjH4uTveCcEBBnKSmIkXuih
pmXER+TWew7+0rXmQOOZDPO0I8wlcE4DLF8kdmK0UC7F75CIKtPAethZBGiEEOFqSNdYgwHEZAH3
NHzLvymezuPOQ60AiAY4GEkSSOvHQ7miBDty5hObngL0Kwf7s2K/m5IKlk81+Y7LgWouPTarxzbk
aSlqsHA06hViFdZKccQatkpWutVROHLjVxMjwPGCMiGFI71n9LUK6NnESVQDmVcoxcDGlU9lH1t6
TFn/OmTyYsDWKpwHXGotKFT+1DdIFPLXsvzn0w7nc53FWEzayo/xzOzTGWzdBEGuMqCQy5bXXVJ+
a8m6b/BGEo5jtN1JgZe5RTwfmYTbbYv0SlsJQT0vkjYmXLXmvzDq5Ko/5JXVVm7YH+cfvnYfFXlK
hlU/+MstyjT3kcTdAdvhfIXHRzjpzLLyo/hIIn5cec/PA5c+vcLw1+gkdG6i7qGSdkoGfd/iv71N
8XQfFrPrx7ZcWuqyYM/xoqY8v1sK4pTQG78HZK7nsYFebrlpHpNgDxad339PQmMJcpScwGgA0lUL
sBfu7cQ6zY0neGkUNzwDNepXkvNBdwQjDKnbqvNaAD7MfVqr3y+FqLnqhCFHXs7j4Ybvj7dmHbpr
rOHwd+nqw7APsrHkpI/TwYfgAdRjY4Cwk/VqMEQVAgMmS3slZ7OxXw0yW5eK3fihrbhB6rgB1g5O
VrO1vylay93oztDf3iELKgazdhQ0xgehM+fkyc7yyk/mCoAB5KPb839BBzllhWaQpQCMPY/hAJfR
oEtnMQG4MM6OTM0pMgXFmvKMoBTE+mTvB9Kze8YXzQTaUH1lroFV4JioZiBlrsGjCAU2GdqGu1Of
jHkAeURJnn4gL8GQ5x4DSZKDwyhTKXV3PaJoOSktugJyz/JlWmQqMasIQGBCgcXn81uIoERNBPwX
eMKbgGmr82IOuHXT514+54fOvijMcS1DyhOOctjlIC7mIh2bI04g9V4OFkm0zXgCqkTq2EUt79MJ
g0RavFUxjD0F49V1dWpRzwvFHGTsJnxTmFPwtPlmqSnsq4DrgSK5Yv08t7ImGI1MF+qryXWLlmDc
9uYTcjpwOOMNzhAR77zUcFGb460tp5IbPsEFOfrr9fxOdAzfERZd3+NyYTGed61gmWoPqQttoEtc
cAwfgHk9vRoNAvKD5C2Ne4Ga25FKMnSPFTmiSrrzYo0j3VzA9f6bEjknXGunZspVHBmgkcCs7bpk
6Oo6F+DbJqUkEbUYOHootIqIEHjoxJSLr9xBL5RkVQSqkLh1/XJqC7HuqOeZYiV6uYJ+AGxju4cd
oFdV2IqAVE0e4hB8U7eOjbfmJ/gIQSKRo11v3+b8pF8ZwMnBZMjLs4I+8P0qf+axh8t1zuIeR6Nc
fNYFiA9KONh8ZRrYHq8OAtwJgAGGSMoZ4yEB3Gl9zwNeHRIMSZvdDtjUjiFMs4RJGUbP5+zbP+zN
I8i/uNm6kZc+4v8v6zgc0YxueMie3HOVAbetn70pMLR5H1FjDq6k/BG8EUOSTjS04g53KVOj8nv0
L3pnkFPcJhhe9WBzOrqBNYG+vDUgKdHh8HRhVpgr84I6Qz7geGbkcGXJ94j44fs6OP2pi+ozQ0YO
/aifQDUu8yzQsM3jp4ik3FehVTQbMj20FN8J6XSIdD5Qb0JfOrPXtg8q4tRdmLr/WCBYkWy9KPST
qkddCeaMuJbgOWkgzVl2f1AtkOcowqrn9T12KFhYtOvNE2boeNTm4LtxfzjA7FEgLMeGX9z5bVb+
CLo+RZci2MAsHWKzbIljXGK2DR1sCKAXINa4C1TobZacCZnikhohXg+IxdCiqcU4SmeFfXWc34Hr
PTML8lkWE6uQizoCUTZG1el2PGLhGt+UVz+Ijq0fl75qpef94rZAnYVRluYdyZJ4ni0/Ev8dwx64
MnU4NE3MdNSVFU+KQRVpiT5bEpZn8Wfe3pSxblNCU6LgsTW7FOnHdq9VWl/S5Urb3Bui8tSiHFQP
62UuzeSe4LuJMljaBVUB5yacmUtNPN6BGd0F+jgEJh3G0OzjR9O7/04C2GJPTOgYmmk6mZnrtHRV
vKFhijuoPR4XJ3DdnOmVCQbzNWGWEq/rSfcVIe10g44ftvdvxBEAbsjFhF8eXay+GIsU4NTQmppC
wz/8BNN8FU9XQvFXJN4/JIZgnJjN7RcFmUhCamLyJ+0g5zH5BRgkS1Jtp5dOXhPEGVwh1nwAgZm/
NURccAGonYVjjaKx5RAkDDAdD7FZTt64TeWS7+hmXJXRdgXcIai8NRm1VIqctYhgMqmPfBG6t6Fm
gUFgqgVaSmmeKBoh7tFTcejCuk9VIiwYHlMvroUVHORVOVWHObuc8hROfgb5wrKjQ6wMhoL/f+Nd
SS3BpPnzeurP54Nn2Krp0C+7GdNmcTUW3/YouxGy2u9Da7uMOA347s1LDnlw+WK1Lgk4U1g7a+hc
69EgFqOjVZvU48mH39Twhh7ow6Jq/IrDseXoFf1pOurf1lL0nXNmKgwSZ150WaUQBprVuHCGPHvU
5D/ytPijRawQbvFlp+7kdShtd7U5goIVThr4leZDvKYJOMAa2fYsnxCpjj9pDlWiwNK666pPGGuY
Cs6b2Ken/2P+g/S52x8KHey5lGpUfAs3oKfOuDIGCxs1lf1aPYRsCZxMzrLjEkpwtJxMy3Cr2dkx
HU2WQ8jYciJWWCS6eJ1iwZ+OGywPT6FXJtgvZ2IZUA+dvFAPw98Tv3OP6ebEjNru3e6W9L1DOUEK
vAo2rspRjfcp/3pihQKUVFWAN89wk5qjUZfqWiVCS2BP8IZoMRQZ9oj2mqPOmv2CtUf5W5RgW+95
7gCru/2WCvRWBSdMN3q392MhYyTDYAe5kV+txx1SxuSCsP3svh/wu25fr9us2nHCe0QsGDjGCTH2
vowoF3U3FMAMTZjdZ1yDrN096eiUJSrRn2cJxJE70uB5crHswCeyJuyAPInbCgwnsRbrgodKPs63
h/TL+gDqIm80UWOvGSTgG9zGx2jMcehAlcBK5K3eOc6O1YYlPuJ4DcXIWVYDcYchWdrggUwWUeSt
ZjM7eMrSDESObKz3lUUoluSaR7gdvl/wxYv5TWCTcfUElXccy3YbzLoenDsVzVkJSnhKYJHDK40/
BFI0vryNQKeWtmOhjUkiezv8g3HcwT/BTCPvyREyQHT3aY/8Dp083bQUD00W7gMLJ7bqjL6gjXlo
EcaL4Mat27pE+6ycozQL60sUePbNmrdhMm1pC3sFch2S8cWDOERFMG1Xhh+AvhKsRwPuwVb2+ImH
3jYEe/1o47ICSI7oAG0qMFE3P87v8fbETGzO8yuT5sQP2yD/NMVOZrMf4fDb/SFJlRp+mIXgzEgO
Pnke3U0im+dNvYDga3kHAJYRbJSihpfbj6awrgwqDQg1DTKPsR2jMYPHz1wdhWvwjMzFGklyZTHG
wJruWfIm2NaXsa+VCY7owSzbqKHTaDQbBAAXMePTptckWUxyzqMsvVlfSj3vYLakTsqiHljIUhjW
XR91nrakY2RkpGaYDVLXl8ahowVGxz6l5EnZQUnY0JQbkdZDrOqWI45mj1Ao+9baPod2rfc4gZDB
TxiE+pcr/K5D02Z+4ka/l5qGA89kFH0W6v0LQPNkgFoZ3h7pcysNRY2vAEyCfpugKo3VXJobZNl/
NSFKsUuRUwqXhVwogQsWM52mRrAdVl4Ou77q27wYofJ54l7UPg/9hr2PGDr32tJ2Ruym7YrKzbrK
AviIcTjmyuUe7QvZBugCObtAHscn+j7sw1HidCX6rnI+Bd6F1GdYoVP/rTvVkFzPl8Une+TKnMkL
nXimY0RjyCk9KnJMtJLT1OUxJtwGCH0k7DXzx1PtMsaanGUDPGZVBz5mpkkDfwq6adAsthU9dHXq
255Vm/YopgMgZGJQoX2C251OANNTS5ktPBADE85M5ytS2ab8lRPyGMdrJ5Rd2wgUf/QJJrK+sURP
WpCjhmxTuxBHTNe30OKDlWg0I6gCj4U2ndH17ULlgnWu2uRlqSUvZejMRDLkD0ME/rd22ciX8ngN
ItUBY1r5abUnJ5aiwAM+Gx3DL6gQzQVAn+0GO/kfrqzWgK0g4IRhlRm5y6nqNvuDqIhfuRIox8Fs
LhA7yT7YsAVrpNscBTW2anIwhWE6RAmONUXi2twnemXeP2YoDLprSGOkJNtP1mvOCtPcoPdN29Pz
HOPKUVY2L+SSYFfLmcJiTwePNNOgxFzx96e1JW2VgBawEENw8V26Go9vxY6cPQeg6dy/Wz+DYKYu
VgJKZhQc23sTPjmv5ZTEseDKCZevWAtuelxv2Wp9tncq9VdeemhbrCIcm4jv31i10L/uSvOBwtu8
mEf6L4FO0KrcNvEd9YrP8x+/5CaT6GVouXxxgAqjj7NHLO6nIfi/9T9mQPjrV4m+Wgff/DCtfP/S
wRRoMcQALmQoUaqpfr09m+7rX7aCeMwv4k9r4Pop3ia9iZZYBRIRBQvKl+9pui39RDJuHdOsRzx9
Sdx/LWSflScQ0/JqgPWbj8Q3K0iPDM5yrn+184gWj7RPzSfYwKGlvT4Uj2gaSbEBROqQevqKfAVP
oH94SmdfM/ptXdG5S5kWTUUvStEcEtSYOllhjDzNHAAW9PFOQCTW5hdzjDEPBXVnlf3SHvdZjfzh
NOU5Xn1YLG54dAWJBVZihAExcFzTvtEy+7s9nz97/fOtswVihUeMyffTJ4iR4Sy8BkJmOPV4IhgE
qrEto7gfNQvZwbHdcF3IRFkYi+pztpVf4ce1k+KOPqUWJecVspCGxLF9Fp18gmdH0eHHVITUgKAq
7QIvLjkQ8OK48TZCgOMnY+TclmFFqoWL7SVhylI8fhUauSiAYLkmVfTznRg56qQy0tjaiT1A85sz
VjtPiMXRoUg4k06sql6LQe7GzcbEmSnlbJC4jKAmk1dnMuzIRpneKeLuqtHjRDlvs2DMxPmZix3u
yqbH6mwkTXovlaon6sKRSmp0xrXS+pc22+59HHtQo6LnKaqbBCg6rxdP5pQEwkrvA2ffO2ub0Q1U
q6Y13VJBrC3+rtVHQ6KjYv+X/kliM54vb7pWsHBtGw9j5FIpDwsTb1ftcfqZQQV3BvOM66IFCJu2
dS3gTHxP3x0rZnzRZ704/sj7yqDI0R1/kUSBjXZuKJQT6ZnzgRGrvA475Ac98px1r7S5ojp6/n5E
1YCqz46QbEfH2kTfLyrlWRazRrTm7TMAld0yBqG34q6Sao28PT+ko8F0Wqlncm/K6OPLHYvU5hFM
i48w7ZCmgKJy8JYw3ffMRRt76IHo9r4n0e0J63nanVLfCPYaWJ0nO9wHTx77mHr/uF5Kw7YHgSwi
6u/QotQTqRGCqCMYZOIO/XIsPIYV44HNDVTjnL9mvExzEeSj9OptV7S5avevfpa1VmQhKmAail/I
j6GipFblWOg2KGKP8BXc3nqVMVc98nOqO11MLq4xu6wi6T/BKamXQG9X5KF7xWYszpbJjzGlIl3d
ywsT4PyJhg56RYN18xfGbRXmq/sW7QSF7uXU8PGn4u38OKzaR0PHS6LH4w94Hx7zEVaqYvpO1c7m
uSSxLWHjNgoJ8Ks7xfZ5+93g3on4cso262BzcOWsZQ6IbbZBstUPBmmIYTZPNu/x98BBHyTQ5jHz
x4vMuxpLaWVAPdSVPyccD/lpR7G2i2/lqV6P38r5DFkHGlrAR9Cml7zEj0dUKV8IEJavv8KScc4Z
wU3bFACcaC8j3g4iS6EkJMn1PbnJQcgLU2DxyUzuht9UC7fS+R9ZrZFW3AYCtPJU3PYQA39s3yTJ
6GJs/pEHxn7EgSdHjhqyAPLdrMGbfYIAEzjuyqlCuEt0m12+gVD84VqhcPpHwwmiG81B9b2/OwPg
d+Mm/InKTKi3SAIVTJDcZqdbD2yx6YsAgOW3m8JivViN2yGUHwbKH67DXNrZ0mhIaeWYdJtngXAP
txsss5J/KdNU/tG6jyOEIpYpaYpDGw6Vw0IkY9jfpQmQdgCzAlLKiq+FIuQ+Llq7fieXTVUwYD8Y
gvqscQJ4Voyo3v/LcV1QOQOCGHvtAOujuO9ZknFCLB50GbtDCwkldTGN8Ha/S2PVPT5x24ccj0Rw
uOcrVbZokTZtSTi5uwrBUfjR8JOcDJeJpqXrH/zYaYWwcmgP+OJlfbqDRvbNTkIRsEjJdRiNISTv
8F/AaXfGHAykDjYWq3PA5itYiIs+A5UWKWcGx2qBHRReocpKjSZ80IjKpRAyMrT6CcaqJ+PRB5pu
E14IkwJ76MpulpIzxqJZMqKjSN1JBNFc4GMG5SbOehhXJdaZFsbcEpszL2pjQzYKc0/6C0WRxoc3
MH3HDk5iTcPt9SaAgECKkQorOUCR95WJPTEmZceXdlJz0VRgZ1lwiVb9tbCxj4p5TRo79GqFiu03
QXzC5INaT4wApEUmy0Yl4sGR66f8ZUoDp9UK2ldGPCbmuCUZSzT/YERAfcrm8hArudrVzngrf2A5
mUQ00W1joMvYyPZSolYsL1RR1vwPNM/GnL3cFe2ULeBt/s57GGApYsaJPuIVMpAeGVDwLOBzr17I
4DARGbfbDLTEVj2pOtlfvbB0vGs0K9TLuW7cucPAu+iqZvjaI0RbgplBRR3T9XGN6DbU0PRYtrGI
e+msdUSEFUP9PqPzD0Z7JznI/LxfjBLLN8tE8nW6jNSdd+TnHgmK/3nHYdOz8rolzn3qynXqyS60
9A0LVFwJRPhbeYDDGd3j119PBSueZ59U4wz9bmGXXasAEOG5GMk8UbE44Z12Fl0Qv1d5X5YHWOhz
ia5j3rDeS2sCbBmL4s60jW+6/+vTdyN9V9Fa4POuWtifRNd63kcs2DW+GaG4LTbqzwiykf6pwyXF
H4BXVOUmW7yorL7zDr3680I+ltdx5sVVUTfqgwEmRvD1sO4RddLgo34wqOSvDg7FGkaUevZggHTK
HWrUvyswwHbZcq+GcVFTCLHpUreqRe8DN3gAMXf96IKdx6V3kjlvq2OBRs6W6awDI9GCCo+ITIMp
+KMy5dJggfejQw2GdjSvSX1hnwjNLdFxdHhV6G55zCHSQd9stieSMiDQaw3SU3nrX5b0Vnb4xNuI
3t/dBXkAYyVAK93e9pDkuwPv2roFBHae0B5RVPzcC7kGb/oVh36sWljKwhoNHXiNAq/l6Sg9459G
ujK2hN8ynyG/issMfdOiZI0Je711aV7omO1z8hJkNtnDfjt35fdn2qwO2CEMsQIrQgy6vjqczOIe
Qu0StqhU2tyYlHC4kIf0qMqhyE3N+t3AcHWy9lX4n1wrmpUcVWqQqgNn3c4bZHg0tjg8ZHb3uRLM
qIksjDIX80uduu4YBLrelQHC9fnc+wrS8e6USaKrjguVU9SlMBLQPYJwc+ru1qgIGXz+GWOKWMdy
x8UpZwV5pdRFL26uriKD3GCqI3+gCe+YGXQTcQ5xSTOe0TzByLwAv9mQqiuF8UU271xTEoOuIn1a
3gXKv7BBZ5CmhbrXgY6BSb9CiUUsw5/LVPW6E00h9lZBJn51XK26GOtzz1W67SgFWwzPib170CpQ
uH4eLvGrjchKZRGfRK3/pp/eLEv+FfI6D/I3XP4hvbRxqclIORqK67ElyYxEH6JFcpyNQROH/DaZ
OixFLK80+4YJQXOJ94RbpWQlOZHkFutO3A0zgxNt60kjI4d/eC/cnsftIsuJbY8VrIT4m575w4w7
kxbzwkMegGIsOutnjt9z86VDQa0TLGI+8qoGUSgS+wnsUTjwG/3IH/BwQLagjwL6iaYNpgxxovhI
G2gUM68W4cwwuKvxaXvLYFaEiQCiNkeQFBYFExXwbAQ5lwiB5FDy+F20K486Dd3hkNok4tARpN9I
1Tvn9lXnjU6cqIqGT9Vi0GacOX78iVQCmANxle6HtKxKs19CO1NMmXgEMcTysLIGy/1SLq4FNtF8
CgtJ6HyJPf15Ry6UQ0DV8VDozrLTtMR3bMEr5uPP/+X57LFl+qN6dRlCPLk9xvBUKfBbFS8vHTXA
/zAO7bwVGO4WHpjF/g2dbzsMnhBMGD/tNdWpMOpQneDlbT9163+5mWrny7RNjua3FmOZkGb0eq2H
AmNxrI9JyFP/gvXlZ7AuFOYeIc0LLvH2q5Ymce7Racqm9Ly2aHaECqbzVI34JSORjdavEmsFfmSl
7b08MvHjLS4leRTBY7VP0+yFzGJ+DGEx6MFXbBHVRugPs30Qy4Si8nI3N81nVmTTxoeveAXyOUO+
53hdG1CraJ2lV4rsPL6t2RWyU6dE2LfLESZ9ofiiQqBLu04VDq9PI57ydvO3FOFUMkMdvxUSOFWC
nPYD+osnsCraBJjSH826Or4XW8VP6NWfgtUAWOdoWlfZtIleDo8JSrBNQdtF4ng6S99ac4XPxEz6
eSzjKMQMByUHsoVMHbRpbOMM+r0jE6q9e5SH2jx9E6FSTKKnLKtGkrXjmKdbqGeF9i9QHrCnSj9L
vRM1xZSxChx3Thxxe6YnMEJr8RiVQJ1mZrYwK6tNZMfxlvnBZazydKVNdpPwJGsN4luayBaslVr0
0l5K+k2vUDwEKMUKDYRxpa2B/jvk1BqRmWOIGkyGpLp3IT0v5bae4+1QWZivhCVplbWspERSGTr1
EajIYD6IfDer7QRLk0BUyB3tNaIjzJBruTn9DRVo0jpHwU10VKDZ/iXyQ8WKab8ow5AhN1mlRUf2
pjKdUq6t/D9KFBVXy5CyUIt/pzToEUIK17sSCnx4bcgnogYQYfUNq3jcRPsY4xmjWSyDCgSIQu0T
uW2PBWRI5AroiPC6WGvC9KabnTEZ0NedvqJVAz3B6v7Dpoko/M0VFKeH9ahxXPp/ei1KJSOlp05Q
9WslnPy1YkLVv8jCMczcLXYfG2Mp3z7J7AOgPlBC4x/kPztYXHlsdKhNT92ThUFUJ7ondyPP2oIS
6GQf2wqyarXKff32dB72HdjW5mQtCBDM1a2uIiQBV58qip3os4QryCpnwodCN+/VvZQPU0iCR5O2
02WTrsNZynrSA5x+TSDlSkYbtLgAw7GtraQMSdtX681Pww9swSoxL/8ZEubd/kH2XFuIPEAe3wk9
KPcvGC7JQvGlcz1WvDu3hebTM7ejfjCZ82rtjnXAPz0OUKrP8stp8Iwkj44tNtbHMA+luxXrsGKu
fVD/CsLJwgV/VYhkvTzu/cHfB2YroWITSKNrvxYxt04IiOIUphOF5FoM/6rNVa8vNlV5E6KO5l8c
e500E9IlALEO11EV4eRgN5frp87O1ojGfF06HbV6nAiVlrkkP4L2AqtJZkwmsAOHnapDiV+xsZxS
8eX+GdearRqd7nVaxXc5fS9fbSc5X9c3WSdXOqFUYzxYxkDqstVyeU8060QI0QHq4aK0gtJpCrGB
0IiuHdulMOvzFU8ZhbmscWGEscXk7VCNVAlx9TwezDlciPzlDzlFdoELvML/QTcAd20LifyPOGFX
uPCpSIG6Mibb0fiMCtaUllIXQorIIJmETkC7u8IFexcCeddnYeURkyf69lRJLOhTRRjp1XYPckPD
3Zr6/rMCA1pCEYYzpB6gtYM39dJ+ogglG9tnXsKEz0BjfyJ4FVwqRXJa37jsfC6BomgMNpIsV8dI
M+hFgH/VRqXwHsamye4c/sO5it0p+tQWFLzpj1VZ4iMO2G6B2aC94rTlDqY5mSH//z1aopMtbcdz
PeZNJYSpgMPuysaeD4i7bzYXjVVHdsp4MHG+nHbvtY/BUUl/pQkQFMcRHqx0WPjWd+78iD5PXSQo
pG4p5SVs0kXuBOcL6Bq33XX3uVGb4q1I3sY2SwBMnTEfuiSozKImZi8dGA/AwfuRWq9XkATcs/FO
2b3m84PEWkNw3Q+a55/wUwvlUnT5PrvdRBxfF9qoAmJUcY/gm/G1aK8ISWqR008V7oUCzQiGBl5X
rK7GK3MuYCyXwRFTdeB/bYeYJ+SHDc/3Pvaqpfz0qgGcDzo4k/I0R1EfoLme7hhdL6aEvbe+tOhD
P/I8Cg+TyipdW3FS5hMNe4JzWJG+wDgfnEOckSpO/9XiLAPjZexSyXYW/MwptjGv+jDOYBbeHcsD
G1iuyZc83BCtll5vNayYT3vUWTvMoZ2vv0eYjN3DRCJ7b5bQl5mW4H9nvZspN9UNEUUTwsKW3SKf
TQIIXfxr09qJYI0jpPQZTl4zD4Zlo8zjkdrIOmr1vcJZ3oM0MUfbeBWHwuHxvdRXXNjZ16o6Qw7o
CLl1OwjL8oGQXX5DLkOG4Ppdj+LD/SMf617qZ/3WZ15sZ5UgXbdStKPPFsiwvEYcAD0BKMX1PGqX
0cZQYmgq373Z0Z+yVjvhqGOecGI1NVast9z8ZsvXpV6GOfb4coGuJg/fLcXw8sHMXYh4j30rR0bs
++QGLuUvbgBHJ9kkjzQV+0wgK8ViPURmq+o8K9G2SVrwdvmUCJhE3DhGMOzkFVageGWZITieHsS+
cJ8EYpgh0ZBWCMhg4YDkSLTbFBq3flSnklfUzmD/sjrzc7cwLfCT7qpVcDudU/GFSvU8r4A3wXfd
PyDpDIxZBlxxu5h6iZI+YBjetNEC7s2q1tcC37YfjXkCDXvHouqW4xY8iJV3UwPNifbbMNsmGGic
r7+dc2xgHD65iuHVGrJy5bW/WMCe1b/AvHLmQIOH2u+2jon4RvJ4sXUMuhvNbb8Sl0yLZ/nJ54Ol
Am58uMa57mKVbKuFxzLDx8Mw2vY2dPZVHiKkZPZns+dW6AgmtfdQFwyoTwfaer8Pa9fxr3EdPGeJ
w9SB72M2LzwPXDB3gPuenyckBPLOhTGuxGC9e2Z1whrGLugeME/ToJ4znCEcLTdE6cohTdJHL6NC
7t8oWx4Lkaj2hDFZ5HYrdnKxWjhrPMiSoUVQ1i5DczkH3cP9kAGTmhSRaStC/HMiqKzsacl1XyEz
28ajhkETVHF+LAW6WT9QQI3x32poAs7Eqp4wzNctqJxJfIr0GpNfkfkyVAuoBTAmwufclyrkQBSa
kqhxzTfvm8Ma8ARrygy4Ykm/TbY4F6GSC4xiy/o6WY+/YJiMNIXdAHc8mj4lx6WdIK7lLdbMVAXF
iEgxf7P38O//gdmpF+YPLWdskpRGFOe7lOwClgmMyZSEBV3eohhrlTomI3Sy0LSv2y6BG+ur7B5d
0EtFtGZ8SqJoRMvn8lfA4DZ3TQTGQaOh4oiQvwjGN10eHm1XFv5rtxyMO9Q8bC7RuWzS8+kQw/n8
TiSlf0a9q8aPKavmo5aD11/vheS1mBlHPyuo+q6F8CPbIlHI8QWeGss8ZvGyyyidHM1s9HZi9j1D
kENB2EotzEwnXy4WtdkgTyZRWU1599u2HVd8VL1I3+lQZsQuGriL9obpAG/5lTMZ6Gskz8pUD44p
YBeMDiLwwZLbT46jI3zqn3/rQoYpydbhy9gZP9Nehhdosn+rQel/Pw0KQ5VXtdQpHGt9MFndmMUG
PgT6WEjbkEQfWcfC8yYZyNnv9w3XQ46U021vXLiwL4oNXCnuZTjThv20QlyF+pwxnhPclXKYPLy3
GdoKgzL2+ODqvzKiAaGdQyM03j2VozRKgt3Z36ifgfrbBKl24pCQilVVkhp4QipT/B5JJvqcU9L6
FU+ddjoheFBO7SDs/puL6PiSQ5ZvSxEjR/LoqW65/hsMToJPb5OoENxsh+7Gp/WlfVnwaimesE/s
vHwib1YahNcUcJJz0smEZ08EFQEbBdS8f2SocI4EIcrWk1aZuBQnD09QRN6Ul1+wxcL4OQp2GzHt
tutuNBKgRKyh+G6nHRc6fx4arwUC4rkcKCAYWHg0jWTnW6FMKMe2SCORHj0zovW9NG7W3oyJmIfy
Ry3vbIq1O8SNZzkIvxcpDX0AuO473SMMV/MPiT85KLNRaFdCVuy9ixIb3meUAZJgQxbDxVmUnMaw
tfrQNB5iv8AMOSaIaENbFPxXE97/THXH0bkdIzDC7xEfx81SUB+MIvsazVEvvo2coYOk7m0dXKpn
OMQf/91zJ8TXRkvYjYc5vjG2Haz6GFwa5vxtJKUyqwjrt18KSnCRcHcCT67LBx7FpWGLiyJvQxHK
O2tluX9zSCmSirs4GnjYUVQdK+OkxgtGulAoeG+EyoEMnmlqvnkuTfU/MsF/stOVwTCJVXRZY/4u
tCd4VcFw+E25WDY0Hidu73kZnYzYnEjbZNuavIvs3n+sThhiOjK05kcUAXRakcnrbxVbc1ptZyUC
TvoRk1uOgAIFfVNxx1X5NAUpWKeUWEUCOMIPj3L79MDKdqjrgp1TZEgJ8p7W5SAbxgM0KCrpn2rI
5JIL8rAFcE9sy3VJPAfEIW6FB2dlG73GAhCZPvSbW48NxVW36RyYPBceYPNZB43UeFFuuS95g50O
bQHticNJPFbpHRjxX9sKKU3xhAJTsZJBbXrIAjEBXjq9WQ8tyScsaiqn8sKNE+g3cyq3pM8HkQGx
1mOVgHb24T/wJO/EQdllVLAZYWgKukRU+Uzlw7mZmVecBctLuQ/ho/15wqmHnyMYs5AOGhDLK6Ey
XPnN9z6rFSV64StQdk7HZbN1eB9wtIeO8uLY6iIpVlpSEDUKUQ6rhZOeWSKeZ0gEeQ+UzwqnlAi6
wQFLFOyHsVbr5qGgBLsuFpp2UjZRnOhmj4zMOedDcalSQ7TDh2QNM+RIVfwc1jd2wpR9bQAtd0Pt
S6rOIAiGxbyMnD6iKs0HtDz86v7/agGT62bCf3PyMRixQ22PI7OkjG4vADPdHDF5zvTqjU4UA9K6
RUpG6knfALeTn7kKWAPQvtiviYndNc/6tH7831iLTKMKPF8Q5SJXVAZZCnw4HiMH8b+/1PIwvLgC
3twFOehBM88VbHb6jvksUcMTJZQg7WPoC3kANErhceuAo56q2Fgppy5KNztsF8T1MeCGabhgtWUw
9RjFbvgsHT6PpuA5c3TyxK+Cn7B9T5wVKlI62H39Hd0U3z5UEqNLBlgIcXYgjSuhhsx5AEzjL5JJ
uizjDW4AS63z3XVMD7nwSeRGbSuVFdIlnGyXLQ0C+T8qNaP1Bq6zFgsa8IiKD6BTvCnMN0DxqHAW
IA4M+7AWEMwAgB5MZu4tyQObTG3OX0g+vmBWvTfQ9L1WP9SZ6H2NYponfthw3fj2QHlxAoOfnrzn
NqqfdLy+3DW5NQh+luh4tbiDRXtw5KCgdSvjv01LIB6a77GPHDMIRGPlY2UVzEb/64YAWrGEw+wI
ziwSor6neyskTiKxYbeiyQJKfDmCMV38jvJBtIFnsXqZWbHofvl6slcYwGQmLB2u/XJ9t7+EreFs
gZP6/T+OTYM22KjqofEekxl9fQEq7UqUr4AOJVjvdxeItMkmViuN4RTlTYjVWjjEmqqv+XxA6Qjg
/eJ23DLWN5dfeH1qvYUKIj3Eh01GBJjhkbg5G/fodvy1uMfZw6hminZ5A9QlMReMyULPhpBpsilM
jFE6k84PSHjPOqu0mTEKzJ0YAeRTJ2fcHW3xntqyb0awOTDKic72pfjWjaK+1LDyXSn1kpxQMcIP
guUcP7dECoQcAyQbf1Szpp6vjnF5jQsOOUuE//q8chUTU0NL9Ppd9V23VLV4K9ASKZNZ9mK2zVoz
mSHbdoKwnoRnJ6TnZb6fMBuE+HDPGMzDAiANbZBwao3MFbO5S5fxU4V5zTeDvExGndlGCIBP5ODG
HhlExK5XhPciT09XpM6wv6/kzXT1lm6Hnyz9eiV4oDSyl1beC2Tk0uTUbwS+Ba9w0VH95Jh4a+dz
z8OZUHW4hRo2Mtfve5AqQgz6mCmbGEzGREYPqAMlZPiqi4X2z1UsyYuhqV4BLzmo3nikV0OS01/g
mh9uS7PkK42jBxoPfI9Y3MLDEtIPoAom01MyRywYaHK4aVBracqHyCXLKLwhG8/PFGFPstc7pNbx
Pkodn5eERs0G/Kab3ReATepn4YKgD+yBRkwsF3rESiMJx864k4qWpGA5EUgV0VPC0qmZCfCXeSTw
9ZNG5CcChf0bHZxMGrSKweJaPE5+hu6R1zQBhYnSMGg7dQpQ7exo959fnDFrJO4Qe+9bEhkBjGXj
e4myKkFlzgiBhkqiwyuf23I5yk7257M48D2FRgNJd1bgFLGSl9//nHovbWwwzJ8hlBVAeV+Zy+3j
M3JEhdN3Txzv26D+2/c7S+QBV7dKaf0I0D4ewpZV3hnXebfCO+O3rJxdi8FGXYvcLHAB/8l65H57
RvLfX7PoJccZ8ZzojjapHdIDGtko7gPT6ywubtT3u4kQCRmmpnUAwbtdiJ9k9SS1YBKf0Kg4lS4a
GSixrV9/uu0gp5dUgfY716+inIs3frH1SWekJ2MeVxGU0fEYaKYU7q3DjwA0KbjpcU6JOdJXQFHE
QCQY9wi402g5vDj6r+g6BJAQXifhbCBIMtI3eK9XAlx5mfJtyPhn/8eiTqMcdh4dSbjUCgHcdg3o
cMUHv6ux9BgUbsAQw35iKecjn0g32gdUKcK4fi2aGODGc1f4B7hRpbkiWFwRUOMFb3ZtocTVpOHU
2PV4A3E+MClaryZJhc3cc1VcSI0pAShIbGQ1UyiBRgLpYqA2gYgiWkSnjmGbcTeyXbeldxexwejO
PZDhkzeBCwcQHah/8fP3AOWJuYHtCoJI0koVpeR1OThkn6ttIJI8eX77uUUeH2jdy9QO+ZJQJAET
Zt/LSyPBIjgHNq9syt06aoY+eP+nPKjPuoOxiNvWApN4ydiofrsgL5WKN9KF0GduzgJ6n1u/kZXU
LgCzP0ata7m91sTW+HSNhwa3QczI6Q6zrYZ0wa1FyIEPmmosv9ls1M5RGdkSgh51zaNxhYct2SGo
iBKA/37v61797o3974z8vHmBDwqXQnq/9Ib+MNK9mFE8jXNZp5NWAZbLNzArAaSzTxtC/LDkVbTP
uX6kS2NSurU+87e24imTVVqY0nPS/mXCx2v9pTeneS5131zIfdfyUUEgN3vczkZHZvsxcW2WyDb4
w0aQUQrxRxTAP65o5Knpzv0l9jbTKx6H02YVs52+6E+Nj/bXZFIZXIfldZV+6xFde2dvLmbfr0o3
s5+5YvQPK4ztDOssqTdeVauUBYkNlwOsfNV1MgKs89llAw1771KxJ73PtWKOxqYfmO+lxBz72TIr
WT4vaP6Sk0CjBmL1tDLN0gL3SAdDf/XH7H+6PZjw4pIMpbS1F9kNaEhHGRmKlvMxxunmVDVL6Nrv
YSRqbRv7f2wTqZJ+fbk+Ox9GJML/MWgCKmIRV9ud5fY9MovHdg50ma1Wa9AmmbW3Aupj3LLQL0Nm
Nt9C7Mq9/m9xnVdswi9rP56tCu3+BzAc+A5bdqFWMLZGZiNlZnx9Z0eV3PHFUp+kIVmOuHCBFeK7
HO4wmnhpsJT3UUn+fCm/7P5mmFAJ5PnXr+iPrTMZVe9dsuJ+jU0v2YuVMSMvFiZb5b2naQqsIlq5
9xxZ1lXkeeZ+p7HLf1EpRFwPb2rSDp3XOt7wV4doNbqNTdDJk+Bk1F1k/0h2seYK0LbV8DPfQA/T
uijmraDThH//vwzj6YhVOUMVmGPYGEdDBPNKPU5xhFDxtoapPtju+io6DFweyx/W1CiCUd72seCZ
TEU0turQ6sP4FgnquRge5bKOEOwYnbFEwX7MqgKTinMbCCm3VDJPswcSOj96nWOfGRXxxXPwmW1v
fozxjUUH4LZjiskCNkFY7YJv1/VDnnUkryR3ZyB6QD4jOxYoUdyp8R8ATqoBnc+P+7nwkYkhIMqC
vh0EJ7+nb+sQA/hvxM64ozytvcKsoBNiiD6SukXlp9QBt5R59QgN5YR2Ics79hgoblZuVrhg+5rT
NLaaa4nrzVVRE2k6Zmd4+gM8+GnKpWzpGLOJqtFWDe10QrIrJNw2YOXn4VGTxWO9jLDN7K1WNmDO
Lh5dtyeZlS+NhHNMZCLBjNlkKYkQDlPC5oC8sm0JIMtGNHKSnWdBCJsMaXHER3MNsQGmEwCYmc2N
tuUfRVazYhWPpQXl6dMdqacCGbeF4JM4UmYqd0w2m9lxQl+aGE30or3dbsn+xa7N5x/cMKj7O0+P
mxTnr37DVBlLr027HvAa1NA2xEqKIlSbS2YwnqFnoDCZ8uCWSy/LWT9KmvmcJa+/RotLkeyRMn4d
jCaBbd6Qo8TIVJYlJh+XyA0Tj49FHvaKCJDug0aoj3bOSQaTUvYlmCAJIiXJAlVyzboXEdj0LusV
AfIzDI94qK0F+NUwAyymCnamwGbOq12xxwLphZHZH4rhrd5ZEIoNXTWhmr7blOCa+MDh3+Fm67oT
3ULr0wLdYLSKA+xkiosjoA0o2tG+tdcT29OKPG2StqUKfx+cfgPbAFtHZQZOYNY/WK7QcKv5bUsO
nsED1MDbnI5Ne2UFegUbIM9f94DYTMbY+QZi+Cb4U2Q8HdsNOkfVNtq6/oO98o87oTIJEN5zWLIE
t3L3DK+XrJqKCAVIRhuoZLU/8H0WxSQ4SMwPIo837iePLQJp7fUSqpZjwLjgAko3vZnWmrv4uKYP
pKznIkQZ5LswPEnGzQ7ICmYRf+ZDelERtmpJ0wQckBUsKjIa2TrT2pxofZEGphsauFhKLcBASPhf
cVZS/9Xn9BAsHgWN+bsoIWsbOujzXOJdPAp7h+fwAUMQMHHxNs8MEhz0BfGylkuaqsYO6GLxPXGn
uxNOL6Zyivs8KYs/z9pwDrrPi17lCekfXQrnR48kJo0pJS22yTCRbqb0xHqmTNfz89zPXnWmaxdT
hDxCmKs9U/BeVClPm6ZmASYGW/voauy7BeE6UsTnbGC/lZVkWiuw/vLuhal4ZLH7RPaAAJUxnHtv
/A8BLPv2Dnne6vWtWtgY5HhRRfk+1neUstIrmhgmwF+a0GnDcAqaWq/m8yMVJCVKsNuWD8O9x7Gk
+r/sZntUmbPLEEL6kplstZNDSLZXFUZ3d1nZYeji8VNIYw6Y6M1znCytkE9mvpjleBip06THp6+y
barBKv1Xhxbc27tHWnjOpkNdEMkuZbqZ+at8Qc82rEr0uQhMUhLV/4iCtsZXo9DMX72cn48WKu28
BmJSvA9NGbt0/geM+g+LAXlDRAcjvxGpLUbAyknbzrMpN6lYWVNGabfPj+A8MKJ4RJyHXrW8Epkg
EOeslVwp1xGPDD3mqjg95lXuSELZsCTQlIqoI0IeWDp14PshPyxI0WsotUjLwRIXema6D54Fjygp
7Q3hfHyhPr5Angi1YrB23X+FbbRbbHVDZNNM5m1X5mfwry8OMyMpHIDdpZiHDi+oY305LScIvrBG
j5Wldx0LpJ7piofzaDLwDE1nbpMlRb7DtVH3eHz296jtdh/ElWVu3DYcPAUCJf4M9Pcm2TToEBYU
MHtbC65R3+BJTeLQceW2UAJYucJJM35RwhAuUPhqx3T2eIMD0PuEcnGuws0edG/4+lIcAlCXoFXW
zma9vUWZE3QSOP5GkQzxWvVWV+fSjJ0SKp6O4kSmI6st0eR8Fvc+I6UNS9SJfieO5BtPpMU4q0yI
Kkxj022BUC6fM6j70YciTUgobQw/v1n2zscj5Xz11ePUbicEiwhxBVZRI1o5axvv8rLTJ45fQv5B
XCw+hLZHIKXHmAnVJm2TB3YgJJ4qHrZcGZl/W3owHWQ8WVe+4w1WMJVdJH/DUPO4eWtYVYY/u0n/
UX1QyIRwIkls2frZNhnoSsNOTeYRrtyx+RTvI3MjU9WNBUoghx40/ScNEMaLXNbtD4wAt5v0H++/
dUNbEDmU5WwKMDOcwZRYsLHV1gz5wbfMA2mOJ4rMHWHaCyOudEnDLQD45hmvg7MhLTi5Yu1knNKv
zqs7Spy10S8gPetr2IIPa5rD/8oNTaE4kzdDY5eQEAJ71lhDrCBBGMqPFOvI5xXJcpe6Bx+bqvJY
iK9iL0luxAhAZVgvaNutmXsjQIxYxbA/K525L18vhZ7Ez5UGoViCXbNz+slT+tQ99q4XIrRHx1Ox
1ze5cPL06R0HBJsEtFsZyN9FVNvqVXyLuK7Q8yJe1aLzjGHIN+vBwoQqZbAGGHjOBfNcV6YQuxNw
GwNUdO02qVqRcQXrqNHwcE/1MCnXGgf1E23mOHw2V3AGYsP0XMZ2BUXHkWg9s/k4d4u5enqewGF5
q4qphj59r62eahQK+ppy+SGE+K52L5bZl+kSIw6iv979Fz5TOHXjU6+7lhDZ/QfMwcDxxo3tx8pP
vJH29/J8nMHkT8eeyGgcPnMlBNSRNRDaRbOsFvVKy0uw41m49xddzZuKiQ9PnmKUgxyw12N7C6dt
Cny6KZYx8tGTsNU19CycbrF+x9kByj4N1acIW/mExC4BOzvYr0tALANDSLc7SJEfhiFI1LOXy8T4
mF5JZobwaPKQe04xBhostTbb/z3mIPAL5a+VC//RfYRoeHkzguUvahVnqH8ZnaIN2eQlL/mWgaha
pOlAlEHCXNbvuMxAr+Za+8eeCoZGLuKxvvpr07QL1HNasrg3or3qrEIt6UAlSZOg1KUcKKVODmWD
Mq82ZlcCF7tehCDcb7ZrM22SwppRgOmHhL074URAnqwqynKPz61mIHIMpkFzhVlP7p0C7NQCEp4c
RPOH6tbmVew/dO9r0MHRe1s6n4t2tLrtpu3rGVwhLxjXSg7YpSmTddhIwxyNgQmAgneO+r0O07X5
bUlYXjHO87FOJXfMn2/1aI3AQp8AsWuCBoeQcWwqPMhOCmhDSRQJARNzuB/BpxMNug3lThlKfQya
FuAhc9WmswnBSUXlazhjDHXwsbJ5G+UXNArOw+0/Pc6tUlsWbF6sBeu6D4qckStr7y6zohVUrkvc
VY0NwQrFegcYvA/5TYSoYk/fDf3xyjonOMhwJhRSwcNkXH5BLAI67Cz0M5HWaI4qzL/xgjZVdr5H
MVbhrErRCmhKe0ag3vw+9l8KFt5ELkbswvrof++W4Sg7Us33DJO9Ytlwp8MseoMj26Uk4yOAiTtC
yXZb/bnuMbTFD9jDQiBVq/PKZkb6Et23942/5sys9SsateI8C7w8d34DvN8/2DCn0djSZky2dBRM
FvnuUt9336YayU83dIcVslpDiGT2opxI34XtFO9OYa1y6dMkGwikYBJjj63Y2hVajnyWW2YlrnUb
ixX2HSK54NL8Ew5SBQ2lLEM3/o9F5tlSS3OgJhxbQhv1MED8yLkx3MYo8xneqWAqkUFhMy2pyfPb
WBt3Kpitae/Mjsf88y9H04jCI49h7H+a7VfDcDkqjBVOU7MG3/AMr3rRubc4cQWcfjG21whBgVHb
s6FRKLTVBfQwkFfFpS6anW3h5E7yEJKe9km7b0MCT8p/SzF142pu9pUwEkHwSCHMLDIirLwGR01Y
b+se0JRtbR3tI+yRtAc0mTn3bWlYM1ATwWs0RFumCdA9FXYiO+Z9taumwZput5qTDjP/BpDzS7Xp
smFrmB7YhVgQMaw+ysYanK203UINO8nGMngnhSiz33UZI4DZjOh3oWx240Pb1qkishwiGPc/snDn
Mv+XupIT0slXENa0Gzxa5oB3Rl0AKw994VF3L+abAuyg63EIN3bUSl/xyuReC1dZ14x2VgroN2EG
KoIt1JtdiwQT3UOpz9feOeFZoQRAPnIRxMI1czBgE/Rpyjc8mbg6sT1Dg/DDyqZdnQEqeKLc+XuV
6Zl3HxLybsa0PF6G5kKOBjTRf/Hcz98bfNIZ1V5bCBI4Y19hDjgoOQgxcSVsEBr7zBZvXrrLwpcY
oNmY4dyKimHbki3S6eD+7yLm3PGf3dD/coSu7LcoIsaO+WfTH6NQf8Ua/GWoXhcOpUzfXYcvkm5Z
Rt8fBZkN3JufpIb1Zf4wwSwAtgYivviXIb8i5QoCS7wbdW1rwPaoIGlAjIjiW2MfZog4/dhhNK6+
NGXwS16R3HuLv/jW8VYs0jXgMWfXzqQss4OxO1i+0CR6vKmR7Bl7lVoyVEgnuKwum8XlqgvGahND
+9aYFL1hQm4e7qjD7CyfFzOWf0U+K85O+Z0+lt5l5lWxxxfr04Z32U9k8Q9HZjwY81hjNG1Td/48
Bbf53848pja628SNKXjAWWvTnPViuxs4DWWUTuzTNaKMBoi9hsk+uEs0u5E7z2w5mrhPBBhl47QJ
0LuggYcbq3Dn3D2ZAYLdBWL2AFj2PNAbUiFMIDB9315B1fosesCTJHb5/Ic1UZ+S4IF2UH7PYXi9
wtP0qRa0j7B4avniYN2h4fu17/oJfxhPKrHJBAvUrWfrdQ8k2KHJ9ASI4VYS+6kkSc8nu7tjWBYI
bLX2Gcqmw9FTexpCkW/7jLLbKt8JIlcNYDRA+q9S9EDgGh4PZ1LAcsr1lChD/7JfYroL4E/Ehxjz
iA39iqrWwfl5mLxp7avQLu9VcPaqAs9daL99CyqPNcuv6ruPzFsAGDMP/W+25md5ivPk7bcyY6kD
faKPrPAxDtD2Bp/o7Otx+wWS+cF91mllvYoAM8LkRMPfUyy36SiizN6xMNqesmrL/neRqBAaHLg9
ztCFTqIXfMQrNkN6A/ZIFU7GrgieZcOj21d6aDXJm5ayxtgA8Rp1p3Z1y82wFnSjo5e0j0OovQfd
p1FcSpnD2UJXy+fbNHZF30XG3RTFJAKScCgHs7z29Ejg2DQgQdn6sG785Avr43UrX3/++PLNmEJ5
gneQD7TXjTarDbR1VrY04N+tuBos1wyw+2zlNMtSSZT2eyXAGviLJyCE0sWV/VCoAl6ifY9FYt+q
ZDl1/EDyN6qsyuQMWl2xzCazy7kx3GBeo6SRNpemO8jgAEt08vVaqHkB06SsgQaMfurcbrsYLd5k
bwDIQlRDnkME2LODp54IrodwaTrrYdGPxTvOmsvXigz+orLkfQaBi2KQxHhgkNqfQ30LkEPYT5yb
brTOht0ePD7k9R9cWPiyl9+lkLP98R4K1QU6Z03ngwa7bJnUIIoS52q35NT6RYdjzLmz3AUzg32q
Sw1usDN7TVPI2OajqeHNKZanWycVTuDBtmhqr899Ao8CNX4ZxXtIs5OX05DWcIAC+FB/wJCAW3zS
k3upTgO0cIm1uIVYlKNCH/w4Ewk9u2DLBhToEsBJmpTfp7A5L9UbfZ38q+XdRtOE/Ih2otkIW1DF
npsUQ+l0CwqcNAoR2sTtCel988ggzF+qXxBij1/AlIrV4bxsovyvJ1LdCLo/hK1ERqpRr+lHpYrV
Wu1bBvwJqpkUlzPDhnGAsvxfkaL9KxrLx37cUkHKg5EOsOizCdSy+ZO+8GiLnke8HGi0U2S/EIdi
Nw0fSF1veZ6gqmGieg+CJYHzxJWVjdcQHbWKKJ9TmAPalykxZqLNtFzroz+VI/ARjVSZVEUu2rmS
EJwZ8SWd107JHyqW5DYoNSLVEW1oTjNqj0LVf2D1sorrRiJozTHD5i0Z77BReFn3m1mDCNAMniyB
9pZgJQOqOd2/5fndV4F1YzrKbsBgGd1umh7BGv5S+wh3DZDR6Na+gKPr6IgMa92k99XJdWGH1/73
DFosjqymxXyj0U1Ify4iyEB61nxFhHJhuFzgGMUjb6OEfzrVA0ZyR+fUN/5MrPVacs0CqmOJCck8
NpQ9vHLXceEnM0nrV7qoNfnQvTQGnezHZ+kGJY0VQjE9iwWwhtAH7C4QHQxqXKwyEG2PxBR3Rqdi
2c8mnkndzrSHFDXLN2RD30IFZyNUsx4PAS56ettPYOACr3JIeyYp6uInon9OARrnEtlSVKstW1Ya
LIhAwRw0mnLqDXgtGoOECQXt1P/w5hjurQfSTtfKDg2l1Aqq//XRR/xoKUg2xTi1Cd2F+jsf8zRl
RTAaQrHdPYrsy5wNnVhqxJtB5QrqhlSKdPegJXnuMZiJmiJmcF48Wy9mL1pmefMlkKmeFlIvlpN3
1RUCJ9/qT1Pxsjj3pTARhUuLkAr90KJ0b0QJ8LOnToLjysfGCHmh9bXzrteF9dDPsl3UZ1FDMMa1
doOskpSmw0DQeFO67OSyREeQW5aegH9DxhGNmRS1Vs0zJxzOUPNQ57G+qFPgzXZa8XFvB5y/Abd8
VTg2vNMV5WemfHPB76/xgomRVXu45S3Jakc3Yt32ZfgdUUSuboKMZXRSLyfsFu1kxqI5J2pfQjnr
UY69UtDLggu4kXfAZkEEs0w9BubjNmSIy/Fuj0WxQf5pfvqus/aww/9Lwb0nmzUTJ7Tu364bUoUj
HUXafHxYY6HTY6QnZSGYzyo/eVrvNjVsLm+N3+o+n24u55ypzpN+FAhrWFPaJlw2koTCE2zsyDvA
vDcqon22kbxGaKio9MnLKXU6fkz/x6pTATkf9kSyIDqENKPogK7RGftT40WJVife2sI0Xq8+n5A0
0tVo9oOuwLiFVCwDTEfkDRyNVWSdL/IYSFTd80ZCBgh7IwKGyMaodXvPU2ECyemLyj60gmVitiJg
ge9cYOw7p0MswqVMR8Lejaaiv/qJ6+BSJr3ghS9+WEo/UpmkjSjnheo8/Wr6ottGadlAZlhENbSY
jiD25JVjbDB8mRjSjRiyzkGOOd7yVLlxXOWbTrratdA4UvThCnY3kX9zBXu6jK8mtQbbwQuPa6Zr
BcqzRKY+FSaq3imBUNzoNSyPlgVJoYPePwMB19YBh6v/Sxa3f5QIBh31Om+YS8RssSUZVVCBmd2H
jUHxcradtJQik64NHH00ssy6soIgl8kVxaR/8LfFAYgdyb0gyp/uGYrdXwew7KhzBvItCtts62I2
dyIQS5ayl6hkQOVxPIQ/nH53SZaeZWSlesI3QYVtQ8HSyI56QEEvLsbpnREHE1nWGjl2F47+86mu
3GneEMHSYkufBggrgwuuVGfbrLz5vULkaaJdKOzquLp/hzBq9PJZn7FzmhMd0u0nm26dwEmUOei/
i17CDTQQJkRfmnr6WMMqCf7stcGQXJPfEj3G6UhSGtjm94IHfNYEi8N897ncg00Zc99eAvf3/Tr1
36XZl4bmq5nqx1OZg26x62uFwc6TcpFtbTK+h7UOm7isfGylVj9/fGpA1Berk/9SaQ7EwjvY3y1V
BgYyV57QWyBuyCdbJa+9DR/ecMnyD44bnaIaAS1IFKV7yDL9MzPRdmccPd3FX6gtHk//xT0caJIP
l4JC1Q+vkQOds9YspwA89NCNK0Z22jGrUyMNMHPyqV0MlgAxM5UAOp8IPoPo/o8fgYifGSIp/LB0
p1l4+cRVi88iKrCecFwIlBH4lv0RNI4lnSa/yMdFMwPyQrMLRTMqik1W7b9JDqfNivAd4TO8lqzK
etOgiSWwNWt3aVZILHfwiF+d65S011VreOkr7EI5UV02H7cpek6E9BKY6yWDnaK5ZGFZ6NxNHEhP
+KIEk7trDQRb0bXuwojQlF87zFz9fH6znrsgB7YVI6IDIr0yIDZ/vwSqTm6VYNTqpDKIBnQ/+mxt
AuxrxCldvJejh8Bng3TJ4ooWZUDl2e8JDGQj49Cn890ZoBdboOcFK0BE+eSqIsEB30yzgGpWGdgk
xn3uqzlZaeOWEk5Ge+HRdNcgBzq9brK9cAK2CmVAWCGT5PNqw8wVzxgm1OIQIrnow4ClFkQvrrK/
zA5tgqcHSmwnenJ7HsWfwXbLkGcfAPAt1e1WTRKwayzqiiz3Q0ObTtkb/6Ine41Jyd6pt5cJ+ffR
bli7XYIRnomL64PdbgdsThCKF7AOyS8C1itHhP7dHfh7Y62iuQKQpsYF8gT+pFpkTNaC4kTtJv+i
Dvu867CkoyDs99+X7QeU1GlaFuX3ftAwPbKaniE27y6LaE482ig38q13QrozyVPDQmPv6MLoaLCB
UtCy4z/vPaggeVmQuxLz6haH4FsPArZK5WmHhMir3IfS8dMEV2HIvrpZYFkBZVNY042wAYhmco/X
88z+I/LC4t+e7k+zDijoU+Ls4PmvJs7QDFRBSeeJWJ5RVWCNU28K7BVGRPvNpRlw8VzeqyVYFPIv
GQWt6UwwDnJC5bYwuJW7nuwu/Zc1Y91h5qJuRDctmIOdoFhSRi0mbKbfDjeMcmPfK0mbQl++qWXU
cJSX+IK/EYNk8YXO2oBu21xOD58zjEIktHmvAfHUX0unVxSJVFfUGMy6n3K4QVpqVqe5HpyERj1s
cvpHwuSvwTAL8F33UegPjZ3tYt0BMBBkcKZLuOtUD5Wq3ETtHFG0fQZzeTXyOexmc1+KseBuD3xb
jlkU5QkfXm0/QrGcMxMQOr/+BqDWNU5JJkrRSDFgGMIZ4ad1KrEMRAHpdr2j0E6E0tGl6MCXBrqz
jktC9NN1Mg4Q3/HIZZYIHyKJjmhjgDbFzpEf/l47bs9br2omgxISHLp7eu51i+F7rnRHhHAiUfql
2Aa3/ucXM/Lrncdhq/jA3FnqeefefKMdkUymMuXmBhUJ3own7DG0zYiOBMlXV2BGGmlg5N/x7zcN
+SCrXMYDU1X6KLEdsaDgyE6Am4/dmswqQbjmculMkiVVEF3lrCUd9bMtgr1a2vQeiJjtWpl0XRy8
UgsN37uR3dyLnBzIY4Y3YIj6eGlK9mduxoHWPVGbHHux31aP8kh2QdBlUoFgj8SiMmjytY/WOYc/
d2WZobO3WCKj1aqeXt6yQ7UAQjY0yuF5G4uJjulCIgSPWY4woQtNKQ4p7Vh82gLk33lksT93CkwC
7ItbXIg+ixUfB2CypxI6Qlq91ZW+uTqEabgngk7iyN/fcdoXUHoWS0yFbS4cFGXOqEyoKVod5oZT
4ApyR+TICnUudHKGtAU4rX7Vp+KBk8UJDjBvDPyI5uEjornh8j9i/X1CnCBHB52e4287gaK/5BR0
c05BRiY7QEseaLd0lO8JhtAmUST/6v0lkrFzDriV8FFBFs33z5dWEu8rnwqM8gv+8C3bJqXtify+
ghoWg0fzR8dDcTe1Z5YXcLPFTPEnP0eYa4WdtHiPadFFPX8wiVEKxQaHlxheRaZSaLhNDW4d8B08
dXujALVMYe83V6WnFbHsn1w4FN2nzir75LlS9p28nG6R/MQERRrbKld7DcNHd1C9e1x+oK+lrCJ4
XiJ50ijakrKRWThTHiiKhtgltc91EkW+VvCsgWf0cZEcZL+Ao2WQFF6JxXZVBfM9R/nxr2HBXpoQ
fRfxRCyAb1HoiPRRBdmbRMj4fervxr0HKnA5WSYqOq11eHhpAfINPi7mRpqNuOhmb3FdlRdZZPwm
gZx6a2wS3DscjqXRfNC1Qd7GW1vS4gypoSLBuG1PiXQby8ZYGATrt7DjwyU6hdGDfwVSc5vQQCUv
Jk9sAMTvAxvaA4filIkbokAmOmzYqNn05kP5a40eY0w1qaS/TeEFKfmFgjC6tu4Epz6O3RMhbBLm
kWGjN65n6u9P5RLyYqupzWv1OYOezeSEDfb0azIIu0vBWwFEOfN+Y23BzcgRpPHfj8gDsjLREwVl
uEyzulraxoO/lTEa3F/eVbRNlFZlK9lScxg10rBSZAiFywcMXbpjA1oleF0oHyShYs64nI6n6nXk
Jp3ZaBDg304A/Y/pbAzq2ESTHeD3BJD+0Bh8V8vi6+zIV6Oly1wjoa024hu7J3y91ixIEhO3vx2R
aVmgBaLNYhUs3EW+NrgiQ5UARAcE76ach+r4CxAaBEPS4ck92+BtvUepA+BIgMK6QhNCSZ+bkao9
yEiwh5eryo3omNV2hKBNI/suIZtd8f4wqniuxhZairfRGXVSRwmknUBWGEgnP6HfF7c2L6u7QNg3
aDHrK3LqI5FBLUrY/8vmfp4wogOGjNYJtjBXATTTJ3xJu4olbELetG4C6vwLl9GW1jADSc/UuTPw
MpYBkSes1MT+m0vKqVUlY3Iyers9h8nflnxQqA213qjJEzyba18hTJUY6/5bVr/Pz7IggH3v8cYc
8lW3CaBYKMS31DuCpxH+GI9tKhf7CFOhXRx+KqDbnCUkyrrb7TnwWmtq4lvuDqkd8j6yPmS6/2xD
Bp4I53dmidQ0N8S9MtUbyjk/2X54PXgu8UBskzdmwmGJ0ZLwAWd8M+wW03yhoTu8VAdErh1RKmBt
10TrYvIRlv6ZbLxI7FnUA0iWApsD3vwOUKb2/pfBMSb4vRYWiy97VlFjGAnTD1pQS2w9uCB6sV47
lhorh7Kt/CWJ341KCisEF4XxJ97Ehs5nLPW7YNodHpU2PmBQUNPzl0n9MFPd4U4CPPAPrGKGT8xy
ON/ffe3I/2IRzdIzx0iFYWVQ/Gx63h37h91YjpjL3HQH6p3DX/Tw7Xu2WtpPBp0pVGeFTIgmuRwK
SKn4f0+Z2Lxt7grzMLxS3knF0E95kHLLIZjK8PF/QI+NrL89FIxAkF6OoUxNAeTcLXKH7a+fn4Iz
ay1pA4d3IWQuNRwKRgbmefEtb0D2zSVOb6hA7gpwgFH38dxeDvi9Cw3tTSelJ8UgVvRomhX8A4Ai
K2NgA1Fcdb8eEjj2zFvU2x+WMMjij2T25CNR/PmPMdDFb0MvvN0rYl6HLK7jQLZTjNjC0SF7Oog7
TtLaeibG+NdUqjRZ4NaFYDvzQoqNBqF6NWWfIiuQxtTYfhSpk45FvjRsvTaqcPagpZEzkGc1NozQ
+z8T6qW5a8ZfaKGD6iIRg6ouvJhP5HDDYOLLcMJW1i4jA0aa/ghZ7HPeL6gl36TOMIBu5J6x9zSm
LhUyvc5UAgRsAhXDull0M7UxHVDysaIsqg/faRF0/Wmet6kYBa4VVbILXqMHyeKEmfWqDrd0yLmN
QiRLiVoGPGS+ur370rH30H+jaH/dp7B/UFKzzBxeUVYeE/pv8UmC8DUQJylH6c5Tdg3HP6TLja6P
I15ig+CDK5awVf5fCJ/xEOWEJDIyLXd1IWjseWcZyoyjyE5cOfisVPRmkHkxII8H5a7Pg2NL6BY6
m+l33oMMsJJSKvWltdCYaKBacrvwkl6JPutq1VJYYBdFUXe/GcVbCIsQmDGhMCNFJ/0NC4azfgho
TkzJU5KRV0OrubTZ/y3NK6CfZrKyP96x6Ku1ZGHRvkknwvB/T+DjM0bfWs6PoXu99iN9dWl4CfVn
pERvFGX054/Y3QKv8fo/jromqVykFyfEW7CQMcL8zVS2sQJcaXAdga/L5rm+XveVvCf0bnBEpvj0
GQI8YMhAakvSZ0unb3RmQWjYqLbztEx9fAoot6r9maRsdwotxg6t8YRwqvlDG8hhMi7fX2cucQbb
u+gEZlTej4d9VP0lsq2FRbLnvK6gfstJTTJeztR89mgDfKxOrXwEtBPTMtNNHxALXrlrT6D0l41f
nJ1gIejfd3TfraugoNKBFR2xBKUgX8i28+3bhzYOs+FQz7uHQ65iednD7qBEf7Gjtaqd6a2lt3gh
BG31G4VxAU5yalGT+uZtIo+BpSy9lWijyV0CnpaoLNh9J+tKXj0hhHgqOnLRc7FSeHhci4X28DXp
BKVyvxgBb6Y8viNGZY6Ojuo1MbkKwOM3PFnWZk/D2+KwpVev1OTpBzM5yreMxc0HDo46/SXj1An8
xOLPZXdCuMRq3GNPKgGI52/bLF3B3dDDufsAvLYobRE9m7ibNV4pigfCM0xEXZbs1VdGAm+Gr49z
2G9c9/Q/nTZv5rlL27XFM5yJ27N+VfJrWkeUUGvg/+SkmwJPuoSA1GsppTzeNWj4bKfUAp6Y5EdF
3AwEzhaow8u+KUxDqVynBTOmcU1YXJ1L9tijOf18m+3kPIKOJOdw09h6lEJhbpfimnDoD8LH12+m
BpDtT9zJUzDu7TzxMtkMJV8hVCgov3+UKQEK6cT//FH/VUArugIzMOyoflLF4MojF3wBnwLOhwGg
865dDHaUTp7Lpay24hHl8grsN2w/BwjobyRuhvyxnuOlep1FBnWL3OmXaC19fWiHQhRkPlTuvBI7
pRThoLmHyFXanX5pQqkKRkOfNkDQzRFmJQ/0byttI1AQQN+KO75xPiDwSBwcsE/ji6OECj3c07jL
hbQW8FgIJHfY85DHgnpdCequFdws6C82jag9DrSty661/KzP1g0LCp7nwq3lgqFTHRkGEBWlTmmZ
0o0b4G15gMnVqvrRZcXY/DL6xafUuETqJ532fTxaTqwN4Nc3Sy1wXK/Te3m7QHFED33tQr0/Au7S
UPa266c9TxaQ3iuJBOnka0Dk2WdGPRa605ZsVoOBwThMCF1DkxfUPOX8WnX5ayPU4ADUQcHS+7h4
7zArNEONLpvcl8DQPYVLd8SRYyU1mDCIOYdGAwXQFATlV3jzophYIVsNoVBF25eOcjI75/zvwsHk
tQN6xfn1CviKxg/i2om0x7pQ5ZMh5Y0vOLTxiLh9J9w8swJ9Hm6l/n8NR7X4zOg+Z/ZQ6VMstVjW
G2QUX50oWiZuXaR7aoZNywneeU53G+t1BmKx0uPh3tcBH4XdkKvUtjmXaeTzWpY86EbHLG7Xzyjr
0T0ezz6eFZ+4KJiK9kk0Ay3eESKa+96111LfPkBnp/bAebk6QfK/weqjMa8gzOiJLt4Ij3zZkw2J
1UCOaN4KGIzqkZknIeK5Lh3u4ytI5u4O0cn/yp5uOUY5W253LsUNWCAs23C75idE9p4z81syi2Bk
6G/C/c+D5Sn6AHSv9t000pnQLMOgsqy1jD0tT2oRKf9liRhnTgdn0IaLB+/a71HoxUGjS0xWbNTq
cxuflttPylSR+c++irBEKSFXTsgjKCi5EWHCg7Y1lIDPoRy+y4LUdLL0yCJh2z+ARfGGE6oeJH3L
rPx+kntFb+vxi1/ydDHdxDa7fPVgbgrw23OW45MHytzvW9EGHcV5+NAH+lEqUIUGci+Nxjk3bIVD
FkmcydWTQVKIZABSzITpwwB9pPzpH6LTi2oqJFXm7FCI0Ft2/jBcOhSnww3PssgDFiVJT317iWdf
n7SfAeSGOPeaemnrgk0QVq6+CCEOtIEK79mvEzR9eMXQrzi7cemGUMZAsh0BvqyzQi5rXn7qar5J
Gxq/+731f2VT5v6SAgEsg1d4pHh+/2gCLjHa+LzrpEpfsNV+PlHdROE+yhbC4BTO2z953lZXMhR0
YDoGH+ePpoEidYP5CrtOhxYDNaJootIxNuhgQlpeOORo0NjmXKTVZLvpqr8LWje33SDxxt6GVOLT
K5RFXJfukdAzaEMZHo7mjJxYuSv6IRMlup8ojEhPxzujpYbuRjywiLvGnis+qpVnSN4c6knfu+pb
ACAm6Bdx+ZGT/2YDJmCzUXkQVqgWJvIwanX/oJBrWta8KrNR2K5r5ANoEePvONROBdqo3dENxfps
Cnqx0uyJ1mke8X5tZR5GgAl4TfXdjz4naLk1CX288KH6D1pj38zHwB4IPIJ3qRxSJRJ38BBBs+vX
UeX4lUlJht+x9F3+DzQ9rJO4bxFHUN0+dhtIiLq/lx2N2bNUcBRPcYg3is+kqeSYHwl7repse50K
kqK1HD2gfYG3YOBZArYFMmbhLm/pZcKaNaj6P/u10pHS2YQcBT0Id/N9NR52sUzZjzIO8jcfy2lY
pmkxbtkptoLzwKf6FPneF/1J9RG5u6ZDfmx8SH5qc5lHazCBNan8Y12BfbMlXKAOVQWCd87O83L7
1CMueAAVqYOSTzjkJC/ZdZj8PrZxjwRxkfs8b/MECj+fZYZLT2k++i5ObUCYYCK0VDcolMwozmzu
ksyWkFlXEmehG+ZgEnUB/bGFTCoxKguflQvr4Ox2dq2upYIWdbD/2RLYCet756CCvMPOnihMAYP1
sDkQyWBZVZ73CpRZhHI66abhRqWBk1PPfXKDXARJ6/r5m75io/uC/B8BnguMKdYZhMnP44BC4EC4
btOoGha5dkL4ACbDqG3Z9vCMJCWexQNgaeyFbihIoR6V1UkIVho6TYybrzv5Y3FML8SP2oIviKpk
3UjSOmjLytgHJ/QdJsdLr1K3lX6NNLnJEZvuz3UwgTJi03POgH62/ITzKKV0pFNvRuNR9BFS51OZ
PcFTYOOT9EFYYpEy1VTvpET9ESq/6VeQ69DpHKgK6LUEQHOWwy9fnUTLviC2962r6uHwe15cV1P2
IVTyfWxT0S88o1kwF8/kd7S0ltR8Q89d5oBRhm0LVIbA6UddApFpn+i39esosn4Ld7lNZj+10IOd
68HA2zK0FE7BA9RD4ZGTN1VArjPXaNbGOZJw0DqerA9barUYrg/ZbXtK85hNkp/mixmRkY0+ROLu
zzDN+DCzqIpzP9ZcKpsFDQxrQPUirqrOJkBU2qZRO06v40hw5FXgwUosscdat1xnct5xPqG8Ywpn
2tprKXMa1UDEmFUXkFxRSJFjIOuyjQFU6HzLkizj8rsDu4rvr4+YAOjNq/+7cW8o2ZIN5kJ+gKsI
p8yW/N9jhYidNLJiMjasYm0t5gwDkXoVjdefgLOkHYANaCdJbhEA9bEUGpm5UkVSvbGgchhE1bqP
PExShy+u+Y03eq1MqMTTNUcsD23MpLz0zRmbOgUf4ujtvnyceMkO8vFkTPfftmjSpP9LN4EZSqbo
cm4ckC02pcZF3NUqpeFhKlZFRhd8yxBMSC4edtxJ7cTalnbvacS70UjNRkTHl1SDb930nX2QeLK7
kpD4NEFj+bURCF3PjaUilD9gdqVl0GZf9nkOzin5yg6UqPN44XGAnozleBq30sEaNwzSv0trXCbY
6MDhac6I2Z8WaXwrHr+OM9Bx90ljLhHq570eKUU2bHeN1ZQ0r8kAWw9DWCeyQBd/1/cpva8SaTYx
/UbmorutdqrDEZVyyDmIPoBNHqBiFsBNOdi0908e5DiuJPLaRsmBnJRyhhAT5b51SxZg2wggKYXM
kPzya6Lea7Pr5hkZzhLkpdDxPpYEpm8UUnOwOyvXOwxwL5aEUgmtNPhh+Ks7WgLa5RfJmUO0L9QB
T9Ud4zQpATctVLJLW66UOo4fim5WLhMsVrnbexm2OVWDa4t/EGDZmYHYDLQjcKMpnbd/gz2BMH8m
d4lgiqfnhSoJ1H9xtoAteLJd8UNXGClMytjLxY4r7DMuOUW1ChLZZ23M8RFRKguI7n9YzxaS8fdJ
C6OpDLo6g15kYzI9X+MoEbR1ykfIGH830d6c3wVHJYhjWmujMPJQMFa5VMQx8x4wQTROyaHDs4lo
MWoOoRiJFRtw5c3rHPOVHN4ib5FH2FqEumDxswuK0fbSwGUbfnHbksMz+T0W44IIczLtk2A00SD5
MfKfNw0NeDHLPjkuoJ4UZcyY3x256W+vFMXB7vS/owYzbuVkg3oY7dMie7yj4iT3V8czO9ipSzA9
42K4CSKbL/G73VojtE4uF1nfRXdcV4cr2XKeBblYxLsKWYpPiY45kTTtJChoV/0elGLUm7eCCWCi
v/1RD9zwmhzJLDaDJIZresUgc5tuBuDLCuGrzcGUk+88oFrh9hXF8eAvrgHXC8q58Mp9LhTSXajg
1jkz55qSXkxHCSMIM6V+8IFiiVFFlnnKyog2Jw5Y1xVPtPVlcX62bcf2ltK7F9IrecfT0T+opzq9
Ct393/8LcG5HaVq4D/9DVx3rXd+yrCiiG+bBMFTKJgz/GAi1oRSE9tmsPFoJuBVZ/Ra2yPvOMJ5m
fs6sh6apYEH2ZuBVp2w09YzJoxLmIGArShBT6ZU385R3d+h3Kp8yQBB1NU87wXoIarH99Tr6dCKQ
aI5/8SDY1bwp1QNMok3ZmnKatK9L5eQhuZuneSagJlx/jsuQud4o8jDn0/mBq6d+58WT36ep9bcQ
Dc87KTeBLsE9vf+Gf6ohYWGCJyIHRevWjq65VeDxLVw7j9Lp6iCXuhQL5ftBboWahTm4FToobolY
5hULjvRq9mSIaKTtIgufT+DvuHfBp084DO2HfM5aCDRTGgD/21O5ARJrT8fjOA9mJ71Cvzz4Jov1
jhkOj+7VQ0TxyqVjHZanB6Wces24/5SRgRmPI4palYmc0hvwnBivBfVBmn6cKQXEdBPiVhdVboH2
wqrB+EBeyMHQ+Xa9IkQHSqK9vFjmy0QcYsPCtS6jeFy0zKZ6bxkbMkMWLrbT6zEbmEIs07VYiNxW
23gTpEu6Kiw54aJCmhYsIDHZ7sdZv+t+dL7QKYqaz/ZD6EXioxwmUsFt7y0KO/ccZIR1C4tOic/q
gtyawik8eqM6xGxLfKUM8O8buCTavrkgYjV4glNxWJ0VE87VIELnWIsdeMn9hfecfhbrCUTZTsks
g0pdQjMSf7A0nWxPuQJhRSAkC5DQxKeOYfIivcIE56lUW2ietLDaLsphYViiIJdW+pkhcuPArtLD
gzhcACD1UGSLjOI6r4ijh6CKOdwg8S2xQ/rs/o5ee91M93qDV86KjQyU23geNIO4QYhPZ3s2nhbj
2AhhWosGERZ4TZJKPGn1Yf8t4dgS0UZ2jTm4A0ZOfG3nmh2U2GkSJIGYfwSVeK1hn4B6CwqTF6s1
2nEgG5PrCC144xLpQdgL5IEA5O7SWU22O/hUOy9MWSn9WDVVffBK+BZiKAUOSdG0E7o/FfFDkynN
e/8tiWLfSM6iL9o4sihx4ztBFodbYwxyuHuVAGRbts1bFbhNQt8MI0+8ClMQPtmvajFOfJ+lHhlx
7IUMS3Jkxn8bH09A2r5V/pIqRcEipppLhmfBbbukqORW36CawhZ83nqPh8Wik4iCk5ud5/3h2yCA
l0QTB+UK7hV4/ydZ1H5wiIWj2oNYvNEiGwim8mHv/5VmRNMQj4yspq6Ze6/iTFP2MZoLCk9YZzu8
yz7wsdRQaiZ2Bog+w03yDALTwms1hu2JM6lAc2nUCswWAVUXc6VYcnJU8rq6ZEqZi3+40KaceEG6
nl8RcTdRZajh0c3PZb1JE6clPBjSAX4bpm+B1qcPEivAtto5BlrbkY3vl/tipIzMQbdhLxMszBiC
s0oNk86o8Y8rj7YMT0+wQlW6aZU4hiH95ofyUJzMppd5j87DG83QtY9qA16aoKJXzehcii72y4S/
g5j9EBKZtDp5NA1IFRr617+9u8Ssu21KkPt0RR6K8q3T7ASEi1y0nT0K7fZsIPGpvn2Cb4uy8m7p
KKnd/rTJzQ5LrChmJWb1ubWCBdWaD5XQTUwY8iNjqBgaxFCNXOOf7gh3Wz53sfOFwcTzYZyD+4wf
kPToLBS0QmATJHdZUYNdthaSBIJhyVTEuXpo+LDA1xWVS7ctbjQC/qmVdYO/icgBomoL3Vnk+zsM
jGSvyBvIW4sJ17cqVOYmU1ejfZVHpvtMcW9pb+ecfjc48xCCnx6XQSoZA+LuSwjjUn3knhNxkntB
UNo1w4rwl2b8Y5kaN9opXHv91FtDXxn3y3bMWAE6XqNllkHDrjBeqCYxjX2E1X4eszdfITctEFoy
0DjTNWuTe5JHHD6ohMX8EXBQp1gQl5qKwRPPm9jtfXLirQEOC3exf2P+vuj+wNah/Xu0gxbxh3m5
yqUG8b7DokLBsk6FPnPFh8QO1TfjdlMxCBvwu/uCVYR62q00pW2p+LRwl08wibnHzuCYzPJllvHW
qZX66HN2a6sxfSrgKxbVkrKQMgzacmCT9zFec+NTSiQIOIyjNgHunMCu8skCClNJIk3dY/86Z7GD
+lyOxRnFtX3lt/Y1X6pFA8YvUS5FWOXCLm/zbtxxDj5Syv9M96aXNarjb0K1rHrBTp7b2x2/TmXX
fQk5C7E2SEKC4oduPe8VhWNsMV4mid1X1du/0q3bTDDSnCPSPF257TaHjxr3dTfYD+HDOeQxSGm1
4e7hzubFnRFZHXi5mHJjxAgQoGA50wr3bEGzwptOwC+SgKVeffdD6Q4zeArBuUDoaQFL18y5vAz/
U0rMdYsDGIUZozzkjoYVmjmdGHBAAW+ES3Ao0Rt9GiJuCC2DiYqZKxO0kGfyGiSk/ZJGeo2onuT8
HPpD9zm+ePX7vtpMjLZqHJKVI5lvxsbDXbj9KgI7RIhqduf/bZ9ML8H+CCw+ArsF8yJ6qBLAB9uM
mz4QdvKfjM3WGU5vbUpxo230Tzr/0oswo8HcF5ABzgRLC4Uc0jBi/OIpyliU4bqmkwSJS4KLDw9p
TBQzwki5FS6fo4zWTtFX77E5dliXEYWrir8gaziin/NkaQ+EO/8rFaRFSBwWwOu1q3M/eGUMRzqr
jNsC9F2I4pBww+bWyTR766VNRk1fu1I2id+Y+/HaccELJrd9Cn8G3HA4d4SCC8k44TSi3A9elXn1
wOK/WOQuekmaJvzjxNA8m00kQ8OilbmvbDMAkJNZBgES5CuFGJv42ekDE043gCbbNlMYesEgbVHt
tmDGG0jP2ieQYmAFAkJ8yfjuxT0nQ6jCJjfYAeB3cECPjxORISFfSGR7BlgKQtplrk+gVY5D6uUX
UW98wGOUUeOSLmxfF1n3nLoPV0Sgka45U9SVR1WtG7MaEEsmduhnrEWfLCpA3rL/R5X3Ix1NE0iu
SSpYc+CT2LuO++9nDvIUTqrFJJEwOstEM6UzWywyTxfCrQEkwBGkqX0IazT5JvOrXGQt6vH5SWip
fkwonlaMg93Cd1+LFrUZ18P46gs1wiTcYFcmAI8THfdm/CEGFUzyUYqYmpjAQZz3eojuFuEKf6Xx
BYkK306evbyBIAPV/3j3o87yT+PVdE24+PmH9stdabMXXq3JUqN+b4Ux7Puf46yTkSAvNF71TtWL
HpPs5liOrE5/GijiJVRxOa+gO2poHmaATbN23yg2e7iI4j5CzDlQWFfrN/D6KAWjGTnzn7Q7SPZZ
FJcBheqA5S/VH0kZGrF2lw3OKgHjXHZV2+FKZbTU237Ci8FcQMrt8jX8NPb11LoD1GDc0PVqYEko
vD+LMVpgg+x49v++TDc+huImpHuA7Aumer6SsvTiUN9ZRM5BZJNmooW4k/LlMSg7SAC0W9G/1pt2
059Aj93rprp+hFU4ZmVw7wbvoE/kLBgZ3yOAUorrgNRHlcb7wrqhFM4hrCsZy1ep6lMMuZBfWui6
5HRSlArEk9VF5LT5fSB6nKni3wtuxKbD5AgQpHY7nrOnj7dTtsbCU/8xjByVyu4y5HKaaPje6mJx
qTj+LTwiQPct1UWYhTjmvsb1H3vpeEH1GV7q0wXOrwcciSHgZDtd1Ef8fA6BuXAqojLgAdoj3Ksz
4rx5Y+VxAEM2mOgI2HQ2CuV6AaikMhOv4MyZD7Xz1gdl/1+zJxQnY6XnoL6gbgITBXupDVZpHKT/
E91x9qXwT3MaRvuBpY7qYMA2TO58JARFCF0CiK/6jxupXoxzd5c7bj+29YF4MQf8ghKC9NpeBGF9
SI/m72x4Bm//2Ck1Ntp59NF221V9zWbg5JaRDQEmBZIR9ktcxTMD14Yy+LxT3PTX2OSTB7rWR49m
6HPLZ4ZRyDTgKfHOdVs2UAxPEsRR49WlvsWZlyxv517RAfo4/krxrzQIyXLgNqZbjBEWLFrKK89K
vi+D6q7RrxQb0QJ0ne/kX5kNgB2xFLKfGY0Fw07WD8A2NUvo7ZLV0fgxcM2ajmpIC3Aj9ZOLF/9N
nl79G+sgjvEJ4lFxI/pWSqTmR8JIBPXM24w1H6kxVeVLmHo0Y2LtbZqkSGRIbobpdxpAdGKwux54
ToiPlAgoO/hN7RJ/PN3ARJAGdBUqaTsG4bXl4mXoyQ2CDDqI1RcEGq0xArbbhPiWSworX17T7YoF
Lpirb50/VRt+b9gu2O7baeUWkis4xXvZSWDF2q+qukV36YnxOhsp5nKQbJYBBxk5j/XpX0J4ZwDX
OaDx7ja1GvpBIdsQ7Qml/m15A9KwgPnc5LHaGXvyx33KilCVj9TAhZb6OJbzv072aTsFGFdWT8CL
9lBa57QBcD0DcoBg1PsR5yyUDKnIR3P0kdGF5661HpMoawA3eVSl3U/aPwMzfb8mScfNaTN/y5qk
wjKcU1QTJfNZSWKGbqGJunu/H57fOhoaH2xGMSFOw2FyeacVk3EXUILB6ucXEY1k2gmC1DXWPOfP
Tiebi4tt7PalF5H8BZ2hN1V5bRifxD8wczSDKSKXi2JGPcbOlEDxb5vHqgDcH+0xt4NrABlJp6u7
3a5lKItmedkwlvZs+gyGdclQLl0uddqFjSKcCDhOhPpu/xPZhxSZDrhbhC3AUlKEztC8+zDcvR/Y
lOOmc6wsz9KDSOpHW6zuw6RcPHKGIM9jgm9coJrAzsmH94Uq2EikBE6+34qeaOyZU+hTWBnOPaBK
WhafuAEeW3yeJLxZ8HOIrVunluU29KnBEZ9tuOoNyWuXyxEbvMQy0rdOjQkUXCu5k7F3774csUhJ
4IHgvHFEQrTSoWYfRmvLV3aZUlJV0QQDxeWV3NBDtUBm+1nzLD0d/TgIgrIv/3yj4zoJih1g5zLm
7IToZO8RyjzDjUJ1Ay3+9BNViPXozkuC4btVTZaVeGJ+DzKTS39ijVOb7j/iBP3WmEuoFsRxpg6k
cClSF0M0DZZbaGGZEpBEqFbJnsdwMCVU9MLpR0HQrEWfWaS+uwRHKmOufTyuiZlQ884xOi+ec+Vx
cZqImwxEUyzAmJoGjiU+c+DnSP457mWkBQ+FiCxMXNUl9Tqlgg9TbudLBFmLSiw5DZ83uGID7nzA
GzPsnmjIZyKwWUepXNvNn4EjVl1VHFNpMPoRct7J3GWKAhn+HfDI9S7wZd50CInxfb6wTjAOjvuM
70drb2ykXK6q3uMA9pkoZeTcomwsbA+OK3pVX/jALULluP2ss2SAkHefslimIR4ymfs8sXpTG9SU
RGSPpxVLuu96LkQ3CXuwKAn33bxkayGIaD9vMpggoT3XwTfFLd6Br9zPov26JXbYsNIEnsgWuO8g
Mo6j8u/pAc17fzb/R2VDqYLjM+nJeC8qXxH/vhWmWI3qFu74HZdAFSVqt+gEIqNkDzRCiwBNTrzI
56kbq8TaTobI+DOpz85W5k8aUWXVKE9QcduYeXedp/lNeJ2bZdv52U2Qg5Qo26p7xFNO0Bm7g89L
Ft8Z5UWtnncviH2MiDezt2vLsX0c+54i0+06eOhBWILaPqnM7zjifUAs2NUGIQHMjtFmLD8ioAOI
L8Dcq7GCqAqPVYxJtpq37gzrTdFiJT3jL37wTE/WlWLmnDMhhgUd7y+Y5TlzB/mSv0w0v/ndBvre
SkEqDblDRmw/6iym+KXPQ5cWt71jdEwJ5+mmD49ibz4z/OKviAx54T3XdeJa4ljtHxTl5tgbVk+b
6/lMJkmru6HAoCu+edxn1eBQoUQEn3YD5JTls/ajFa8OxPhnYA79/kidO+0I31jCJro776kPTrIG
2zhSKOhG3M9+4Lm6RvkgQuyQkDwh7s3ATH3t+FLBJ6clCN6q/E89WDzqngxd39D1GI5CNs+VIIT2
31A8ShYq7pq5xuz8bHp6LrKI2h2zs/hmQE1vgP+ATaoLU8GktzLH37rOzIzouu4VDVcZrNDDiqRc
Rc88ZQfyaWNwUVADQ8CX3saP2QbWPApkBMcE49HXSu6WmxMyGMSWVNDSFEXkQ3qNTC0EdTMNiU4e
Jb3mbiOXJKG1CKNnAkyWvvEYPT2p8tCaFG18gBcmagzX8pL6FzWnjEuSf52mP1RaqYv8uo0NN3PY
6PU8RzdueUc7nCmAi+neUmyRb4g/aCUj4VbrzOtc2N1NqSvm2xjDK41s5N+dbE09xuHtPD/DUZVh
DHth4ifyXj5V2GMAhwFXSqk9QQnwKVda22E+faTto51uY6FtNwaQD5o9P6WOB5KyndNGhsPrsSWl
lkmxA2PvGFUjF+ox6n4u3F2YTfzDzeocpmLb1MSptvdUeawatVE4jYqNxTNyIVqx7zcVi9Pmp/B8
RCYAOXGyIPXaLmt5ThGR5r1CMjTwR7M84pLn8nxNND5A9hBfKtj8O5+cJjPRwbEBuT+0S0MHVDes
SmkjEsXyjy1FgOto7MshpD8HR6rNnkdVzbcFHAsQrCgG/o/JFSF6Ga4/q6ifI/jagqrt/G4VxWj5
Hzh4lAy+YL8pnC2q+WZGuIiqiThdaH5/mTOUUkBV/Kllh1Op9VYzHXOfeSuFiazyPJoFnALPJXNX
6Bu3Tkynt5nnvv7OKC5RY4EjOUsSP9wS4Zv/Cmm/yWbJFpSnwwJG7HLZWFoSBx1gd87jOMlCTgsc
VkYy1HYQNDwjSqeIy0QpG/5Fy0ImPoHH5aiio3kinj1ti6ZA1bZZ1vrKtd5bLR1LHKRDJAYVAazG
U7/+J9pHb816FgGRTT2V02gp09FTV3kePMEVPS9NsIVz2HZadGRZzEhYF1cx3RaO6rRDAbNJPdur
mUqMjT1MLDyqZI8Wi6ahkIqrFj50GGPbJQ8pXSAq1oXbhVpI7Q1iTKVeouTWQ4yjmhxldRSyY+FF
cFBzaPJ60jiumEAQO9TjfkHH2awh5RWG+WwYZKKYCH4Je7NSX10dfdwwEOJ+20dW7eR4t/2n1MI7
8Rr43WU+1Kha47H5Ngj7I3GcqGvcRFzo0AVxRyRZ5mwm26exaPdu0UYVh5evTNEuDwHtMFVUujz9
nT4NxSNB7In/EJLUxfOxoeiI9N7BmbloWxIL/jgAOybkO7eesH46YXVa8KNyHcSRXMe6SJxhGdQi
hh8+s3G3C5IRZCiwdABcADpFSri0NOg2wSaJLMeyNqpilAjId129cdES/JgOcv+1Lxy0GGv3O4b1
Na7JhhPix0/yw3uyO0Kuw9b7l0f4xQ/+AgnOaQYBWxqVKY4Ju1NrvDo2miRVHWCexSflj2L8+ZM7
xwIgvVCDInd3OQz3I7tP6lrfma4BI7iLvlXXcZA3wGud71YRal3L6KAHSDg7bFtpQxrc78QmKI68
UhCWPRs2Frvani8lE4odB5NK1e7Y9Z1lwft+swYwfOdwIGjHj7b1wPOPBkMz1mXHBEj3yXxerUzO
J1IPayUw0AGZMbjetU3thL0uZbBKxriYTgIS/VMSyB5xmXIl+LGZGCxQZlVUtseTs/S+PvesdTJf
0qZnK1BQNLbnq9+s0FKaOYfbPqVHmyPuFYwnpOy7DllsxC9WRbbCrj/+DpG4mnf/tmCXK8hXT4B3
o4sac9HEBkemWPw13Lt0groN3Q6zL1OPWq9kmd755CuUOSAogpxKJzoR1ZdCtuHsX8WDUdq/PA0b
omk1huaV/6XdwVd1KH0griLcMw53PLG/VL0H23JzD+MVJsmtz+Dr2uUasOJVhSPEt40ly3nehn68
FVowDo0+d20CbmeLQ5sMc9FaNA+82tz501VWhNOOmL8sL46zPbmZoL26yp9mhwXiqiRT1ptXqpwF
x0Hs0TLUjWKI3D6Zro6N8If5b3mUlyXcudwftFKb9EyaaJx8qHJETRy6NjJDnP1Nj8HVdTzy8GMh
Zxlw2/RhuGKrbWfw93unYYi+qMshN1uE9hLgSCip2lM41jwZVFTVe6SAd8+7TFVpOE/74cA6+z0l
fIM5Im+qTCE7nJqefSd7zT7fX6M5QW3RS9ouad2FArO2U5uMe6At4jZfgy6Ih0L8P4wRWVD4e6Eh
i+tTHpMk2QYFSREcoaJjC/XjmwMEbfukY0e8HJ1l+wEfSUGOmM9jorwB30vbepIrt9dNJbNhCyON
WrByRzNZUW0xi3HCm+Na6A2G2rH3SxDbJP/O/iZAebZKd+FLC2U3Ii6oCct/Jx0QGR8DdtG1NSRx
LrYWQB7eYjbb1brEFUKMJj9Q8UwGN5ymVM6uzn14wClpkVl5v8/M1pSuAtPN+tAvFhJ9IR9NgQpZ
NvHmD2g2N/XkJ3SyHDaFM63q/nSQXUC/06HaTfWbcdjwa/6ible5UZIRb9BNYU0DkWYvly1DNBOS
GfUQNzq0ro+2jofb+PJXuyHa8IKSZFvnGEfNJX2DMQozDbDIXrpHyh2kJ8+YeQ2LtzMFGD0NrQ+g
pBAGlhyL7sJ2d534CTpCK4fL1rEdaQGgp+pqhwml1Gny+9pZibOQiqybmIs884NsrvbwpnrJthe1
5Wi+r2aWIIp2ZdfZPltFNyZN/AQBqnNLQ62n1PRQUj+qgiIpEZ7HYOsGBOs3NcxQol3OTZu+3FLY
BVUDQ26EswGWJtzcBc/gGNkn5Og+iaYvcmGtPsydBluHUICHZhSfT1RutnQCSSee6mPvOAuegp0h
PQ58rZKZKI21vzVcOnOqpYo/Sruj24qlEqWcyZBHwu6LJshgrxWmLFNfmm9dKp93Z/grSYhXmG8W
oBFK9s/3VZSx7+6YAmIw/m3umUXS+Zb3fHHQEFMnBuKCSFm0UPv761ktsprYGrGmdRcqN5Xsv2yI
BZE7T2PF1VIY6+aACr6gved3GRe3pCbDcJ/xld5j+jf3mX3800WJNIvYKSw7RdI/05XN4BLI/s/4
JNDIS8BzMQ1CchPfw4WQMIZujxI2Sd3HuhntCGvk7tONRvbdPYmCc6FAn2fw7mcQA6x9hJCqD1mk
bJiha13YZtBwwBqVGWcaLNCe5xakykTdJXBL1L4L+fKa5AcUWR7uVBjjNYZkSrV75LBSMtXVW9Yt
pNDnrtnJp9lp7u4GnvQsE2GnDClVQelhheUaSsVvr5uIgE7L7h7ClSq2SG2NfpAacWjlUiPq50qd
TtrA6N4xS5PF89pXC837JLOCv/h6RCbgaYWdyoKDuZBDx8BFGFn9tLFioYKmAcLn/Hy2OAuM4/AQ
CxgJQ0X0h4mcixuVNlmDVqPQ+8MNKfNvdKTPmwDGyOUoEVLVnubrBUgXOzktZKTCKg+/909Tw3XO
sA3y6XoXgWdt/dxEu51Mds67Pa+996MeaPrsmRcLoxbIHTo1sTK7WbEXYXfkQu8XFiJJk1SbWwfj
36OI4pYhGWXYVH9qnFAmSyNc34wTF/a18Tg2ZO6b2aZ/BLLHcyH4TrZ5Hp8jnqiR8TLKOR9/YhJL
9yuwuEEow1SbngJB/rCwz/4G1aWFYmac2twYLTN8/3v2UjqzAxYxz/iX0JbYE+83KzKn+payhXWW
G0h2EDOQRHTMR79g/myEMG/2WCCPYOgHjOk4FQcuB5T4NQWB9f9JhxQlHvXJQYQ33/UYPGkEI60E
a9syBfKAg6DR7O4OFdMwTgTk/uOe313SqTe8L9ZK2rLWQh9JUGORPmGu6jGmbJ3IndQgZ4Fd1/C+
+p0RJlMIzAAWBClu2HeMZqx3l2EJP0ZVCuYwJ43crAA7QR0I/4X58dBbrbbj8oLO87M4zeQLmieC
Ck0hNw84MXUOngU0vIlDpD1X+CvpcWUpc6v2IJGcgFM6hQ8gL1EQlx/f8VqoRjmMSI7s+urAevPe
GHcIDLnkhH8+ZN56rhk1lbmCtk2I5vtnrWmH2H/xFFcc6akHVm+KJdIYHPOdO03aI1/DqZ2qjB8B
WlJctQ/vCL+JCJTAjOVBs5RM/mDXX4zRnZQlD/qKMqTE6Fj4BJ7XNApp64xvER5E3g0o5nYV6obv
maC4FqImPQTCva3yOXi3zJuk1tOSAlTDDV0UbuTB+Aiv3s0e7V1bTmeZmXwp3rs85HWJmDdUNYy5
I3uJULEY3Rvs9H++Kx9Bd8RjyTtXUpTUpvhVaDQVmnhxG6URttHLfKlTyzt1kF4441YjG4qjyb2v
hsn1OaSX6IAU8gqSrCW9dN440ppta+Fu37fhRaYapn+rpR5nerVDGiYMw6xWk5PQK9P2JiOHQ7v1
gYYjUkpWd/NjRXi6syxWLDGcc95ZS6QZ1fZNwl+QgoKmUfoMpJyj6FZWkPbbPwTIy4oDR4lQn0bn
+pRcbYYDV6xAARlQ7CGw21prFg4Wd33wqYEpy/3618vCGkbbJx5usODGFIFdk41+Q8eQD1nsEciW
t5P0fC/cOrW7Ca6c5Cy9FTycwntc/cM89PC7bElfsfBVhvnpjgyly1R1e44HaEaSXIOdp+DR+K2k
3znXqDjvyt6E5asffyCWLKPGtSImBe8ivjepQUalx1qYYGiylacVGdxMSUl0GmkC3qsI8BdrJOXB
JIDsiNsof46e9mYSm5we7InzYVP5tBHQwz/cKAXT0ok+TqSJzByjdHoPFqwM2xunnXDpBncAenuX
m6qwQM6g9Y9DObv4PN9samCC63TYLArb018JpoAxCd80td6cRr6kRz7usflMWh3pRiYh4iaJN8LM
Eh5HqDXXPENvmwvgq86Y6kkJrrIcADicxCYxLHzrRoY7wIZKNhgrSSknRI//NZQ2tYH/g772VFE3
QpSqbH1pWMaAi3F0BvXH7BFbVKV7Qjq0LpJifPoYa77d2/gs4oZY2nJm3dojBeWOEQPeGVfCaexB
FpwZgQ/Xa8ctJ1g1hI6RvmM2oXXrr9vldgw9NBs6YlsTduo1eQ5ihP8yly7oQChkAezPdUZRJIku
xc625bAfTGjHqD09bdr3d9APN3NpjFQ7quhME/BYW6CycgzSsAr2m5zWsXj241YVAECIFsjT9x0d
W0HAJWihqZzKGtKnJKpIqO0ZgmHPgDpH8Cv5FJR51BkmGsrwYMetbl2xOTXYvC6ZT5fJiCam6WRr
UWA2+MqNdq0CacoDqqvxjM3ANL2S75hxXHfzi5vApIrifNkos7ZmFcG7viyBWCBQUuy96FvHYw+0
7FEW8qk1akZV+onprmLN56qyas0u2VjNus1cMubbvyZINhsm+TmqMQtGtlHsXjtZvzph5lxdXQkW
XdJdHMWbW5a8avR8CMzgDgeaw5XH95eoTWdK3Cjs6CIWbU+GaP6/CY2AXQwI5x8qNLAwAo0XIvJn
qm/wu/qsprN7agCcwiJPWzWuSfjBHD0G0X2OLeRj76MEo++Mj3y6Vn074E+rUuMxRABGS/bswUst
P+vm2O8jwhJ3d7teR7vElhuvoGx2BvNucFc2pisHC35BkNcqEA2ilClNGSCq5wunOzVrXKK52MV0
78/IqptDGbzYNrw7FcgXGv2/oMe65EHhQo7X1pUqwZCmMLCsVVfXJJIiHS9CFiAtK2L/BI/izL+Y
pHCYdyIcIxA0YzvMWTkuY08tbuG+RZCuQL9Y05JxwltFYxQ3lGhvachQtxPxw3zPsMjiytbRPSH/
OJVvfBgeoDHrQ6NnoFTSd6n9R0NTD237esFa5ZhcnI35qENOPeBVSPAOAFPu/IssGX4alRpe4cI6
3b2+u2zCIuy/rNG0/vGX4TF41EF32Kw52WBZwBu67QtrWiD0iLrivYV3RnN3nwMc8WgX9MBb650H
vOp75NyqvfixmTo7l+PvkcldJtBHf+AixBwR16uGPiwwYPUOOn67RKN7pqnUIpjJ/vnbGAwn/Y6C
toZYNA0eGZNd0fKvBS5JqUoX/R3V/fIHXj+g+HV7oj7/0VtP0/GW3t0cbISGigUZl4wEKmdaEQny
uRCZAOhhHCZBL3G0T1hWt/DwzPWecu/EAQeVr6kV1s+bujvXVi5OLfL9tbNJxxwMYUkArRl1ZzUo
IjFfgLofG5TAvQYA7MzUjX/ZqCZu2ntcVOFnKdWyErg5oHMWV+TzU0SKh4mH/lMFJiPoTHcWDBYi
gyMnwywMfZQy/5TLVdopBsvBuwYeteMVOulZaiuKGK2VdcrhFcbcChr3ZKJ2zK42Q3MLXK7vXTKd
lmGg0wTSlJviXAs9/nHzWR4O8fk1TclT8UZzjN/9rW3tEDa79YrZyqUfCA700XW8F1Ot3dN3/zLp
W59+gsBBA7bDEtioCR8O+4dgsOgOChqQWAv1ntOBts+v9RW6F1ffODL1lkpC4iRyz6sV7/r3K5qW
ffpc23gO4KRIydeiDp7aQlpfzXydvT6qUSM+Fj0nM7vgoFV/nEqrJzDAQVLIOXrj0MdxPVm7ehhB
bRXrUA/y3olP03SAf3YzCvc2jYuu2emfN92s/MagS7tWpnXN5kEy4aiK4kzK0zyVN1UY6KzEGnlo
S3UYUJbGYIJBWMwgwzJM/WRTxwKWg71oQvTRz/4ZXIn4AOpN424IGerpFOUlzOVrz7fJ4WRu+dGb
gSOu98EjfTn72IwWncys0tVNXPwyWBoenMb3r+h50N67Soo4x4gaDnns/3YcYzCgWwzt+vdCltQd
8OgfKl1oE9HdrnNWtKVm4N8JZv94U1kjHvsjp0PUkVvbkKpXcFU2zIliczm53qQ2W+yTMOyNU311
8hRRi+G+k7FaRXCb9B151XQk6ECeAFks/LBttgZNDnETtX5uSJ8K0floF4DD7iBpHyiXRY2BxMow
VThskkrcAuqi9LhA0GVKZaqD7w9pLXgaFRoroq/xV/IaWhwpBszHzMz+kozzvwWZrRTda/0QQhWw
yJhiIzSgCIDCouK2AoerqX7X7TRngSSte/BQDYBFT1Oog2C0RMv60yYj21zaxAsCL/rqtutNsb3W
TYxLfuvEez59ZX+t/YAFhEDAcT8Z17KfWegnjRxXWpMwV5wYBrwAxunuD4yd9uk920SYoAAtKU57
xuWpTrMzKjEpbBaKxMPkUz4CZqN7zqeGKCTk/DEzyJ00qKagf7yXq486SMbqJPBzW3xLoSLGmvvY
ls1ltlSnsE45qjUxP495yRCzYqV0EkorY9PL1OBeE0FVCnggeclrVLsFJk4Kn+h+zo0mDWIW23JH
fzVYoHnNk47lqQ47CCCJcguAZTr51tNMkJBFKg7DOZ2VaGtypJ5wi857Tg9Q7PBiBwXOyaBYOmW0
zk6eEGNYHAfb7hNpuh23XKAmqOLkWes7J5PUMj9+D9dj/GcanJL41QVMddkcU1Jf5b/YcNEkMUdU
s20NmbxqrTqs7UXcuvBUq3NoweKDPj0kvplORBDzK5I9StwcitXFneR1uNHtCZEZNlVn/A+OQXpX
IOuK2EQ2dgthQf4JxnQ2vsNBCuXM2U1lYru8ZIhlPn/qobxTbdt5MpmV/hRNtxqdV5hGf1E6Jt0B
zdZC92nScEZ0/nNxBlCZBDL4dNO5yKnSZgjGKhy8jvXKRcHZPJaiugLhkDT1VKahjTLIYCGGvU8y
hjL9YreWS2jlk5bsbD/9hq2u6B/NZ1H+dtHARSBRZ19gB3yDpwiCqSaQZfkaHy5v0/7zts9zNdlD
Xfmb81GhLKthtX4+rtGXo+B6haYNRNYiyqO3N0I0jL6KZ0krjnSUkoBlyx9AOOUABnI7dNXY/VmX
03DT3oRI+GkMRW3fQZZ4tl/rlR7Z7rkd8U79od/Wyq7qGH0tBKT0tNtHcoTItRXzM5WCd5qUmNr2
O+HcyqYBb58r4B3U18LkBSiUJi/ranEdb/In7XkJqKGgwz63RIniuXUbdT8/VXhyTmm+OGuVf6TJ
Hwkib4FGqv5eiHFAkkoBnXRj9iQl9WSHHdki8w9ixmDajYjqXjorfKxS3gtGbuwMpyqlOBuwstO7
PWeyQMJl4H2P77WoFfR3O9CFKbxPKjTiIXRFrbbC2lFYM1HRLKRYi1OKMNcf7KvZva48iYysNKmS
i9IKupvouB0RDdzR1KaAAskxqlvJQ0PT3+HGirG7xNlNrPdDs+LBCe52GrDoEeXxpZ+eTs16GfJd
EMRPgnV8Ajwm84WKvcW8u95UvoGlkjlISntF6lP73jduHBMfoLcfvBV1GZnZuDKs374sRLToU3EW
EVcUpED32CBozcbeNb4qgCJHG4moKZFPZGMlWiuKMuFVG/zIvaOcnIw++NrgkvVvEW8cQwfuCvWf
BFXpKsZVD7Tpd8S0luv6HtK/sG9Zuymz2hNRxzd8XVmue5HI/kpJwXqGwdNKO81hFn/3ufGQSTFl
tGUfjRejJ3TuPJXWTt/gQG9pa9ZCcgXeZu1D2v/xG7+1VZE/+Z7Nqzdxm6HdY/hwGPRdzXS2q9gq
N+T8MiK/o0xr88In4nbxnilPDqiY3izu6uLaZS2cwsd0gSYKRpsLc7mSRWjZh3iC5KRjq6a97cW8
7wypRGPaUpSqOqE6WEX75AbK+T1Fss5J/PVAQtsCl2x/TkLIhZKhoiyeV49TbKx2i6u+UfSxzul2
7rShChQjNBnpzRepdMjC6YnL0Wbza4ZFPFBUfW1YwGmSfNCCVsdoEoFiYVehG5gH2GJKTbTYmUBN
WNItMXj+bGph/08Jfay9GxnwNVfXqsfzUvJUPP+5qZSH9SesIq4ET3CwGW5Hl6+hJ52hPl8DRuWu
iX2/skvniFIz/q3uGpVqzrbGo8fy1wpvNqjtBxhNvu+UNRsBXiMOKQY+y22dc+DLzfg6JC823h8q
3uiS8tZSJpq6vqY5qZID0tlQUjIWid50zK6Yg24IJw3wliaC5mjr8mwSURnz3xwdJytK6E8DSSkw
qfqch570BaW1wAd7+wk83+sIx/6PhKE0pFU/AV6BJUAr4GQQoMXCTcm9H0Opy6QWbM1BbCzaaIBH
kcCmURejt32aigoTclLBhiTq0400tYj5l8MARJEG4x1Cs4sRXnmm6CADj5ZOQj5osvXjjjDtVYm2
4ANoATBBchJo7DrvEURCwySm/RvaLdJMiCmrTNqLfs3dppFJsH2iAW/JFPuNZmyBdGAjhBntRPRw
9pH9ZZED6FrqVwZNS1llBcsVWvPbC9msrFXwFDJVuqxMpsHUB/ydNho7QsL6vitcoorWQ/vxvco8
SK0Q6uG0rTZR73GWIkRZ6FcafdQ7ojqAOy94Knd/hm0g3qL5xh8JpxMiRPy0HesqK0TKlO8oQPao
1VK8LaskKYQ/fWxTjZ6Cy6iTJ3GLR8N/Rn/vQhIhzjPzGCE8Pipk2Nktm2Vz/vOQjBKDoqD73eyl
8grHJ9HXNxHfFm8pWCRockpREIQoinoOkylzlBetAdJG7Muemy69T56TTviNtFezR5q4MXJIPBCn
7qZd/n0XEw2V71PiFnVcykaTPEr4jPMsMojuiN1kTTzhud45Wi+H3ZfMdc6cTSpIHEkR1OklXT0j
C4nLhMcNlQybC/NWwLGkYPtTEfJZ2/hBGCjXCjjamPAYLjFoR/xof4+Kha+dar5E/aN2YbA0jEY1
ySRjWNxakLCBpM8yWGV73bUwbaNg5JPLsE+M6GzarpqOi8qf3SWk2hUtTsxQH9iw6eejWmTysrZJ
axXj2uJ6XW4cIXzxfVGb1gZqWCZ8Q7l8QEV6twmLO0H5sm+9kgT2Te/kNH8JVRderQuu7pKg4JUU
S5GSN0HLQb+EGlB54GObWenUHHBzJ5L7Vb9+STtqRS2gMIt+3WwoZ57MnZTrZajv7djqXSTEm7w7
k35EMVJsSiFbzqLFMcqDE3N4ZpH+kcx34EyJvIk+YPzK16w0Z+Nubfw3XtwfTs85PYIMzZnLeQc3
lX6BxS+wPwx8oxkyIiV5K3I4fDQLLfiMCjMuxS7NKFvLjv/yQryb2bzcncsw5WbbrL69TdP9GHlt
RYKL5c9pauanzTPSAQJiukHenpE0ZDhl9IwUIDA+M3nFlJkU9C3O/rUNgqjPIFPhYlR70IASiAql
VtHg1iDwarOATf2AIwZt88DOyl4B1vvGUny8mmqekothdC0sSg1WnacvM0GvWtVsGbmEtKnZ97cz
7M8SSr5ohwsLy27UnBcZh3T8bj/H/QFLBtpeKcqUto9eqISdoz9js1oJBoVHvo5wtgXYQx7LhYMn
9dliEvvVjVdXIVZc/wBa0t5Oy6kAjJBk5VAG5Hbl81djMR1N8IKQFqSPNu7rkVhoJcqwcxbsIgNq
+GBUnkv1shRzaj2dotSk1VZBXCbOZmeKOPicP2jFna28xkF/3AXBAhtsGKhlrI1cX8E6+0BQRIil
hZyoSNIgvBZesHZeYe3jrLNr+cMgmquDn/fefCjQmdPoMK2vnwajCi/RXf/clozse4g9x8JfIpa7
xEjLiT51QIBsnxXNHZO71YnIqwMQIOmc9R+FWYm73mu0rQL/9Kz45DZoCw7QLWwKEEpn6qJ2Y1pd
RQEBcSuC8TU5A2HQav2J+/k/DsrpTjMtantpxcSqVZWJJvJxjcQ/oJEorakrJlgC3IW/Xqu4KzaD
X5plFNmbgDph+7ZV4Gq/o4B5++MBbPfMghXfwjxG9IqZbtePxZGuf/pkPxJZvdGCKCkzgE51ZCRQ
OqIeos7FaEaNHNxZCMBqbwq96wmlP31luX+3AgB/khRFOeTH6y0wI2nXDa1vkLrXIxeDwZDi76SM
PcnscpdiHxdTV7ULVRDSqC3lJAldFBtOcyUZwdF1vvxeab+lkgNGZzSHlu2RG/g/xgJ3oHhr015Y
XN1S4gxqswF8Vws2XRa/cPWLi5lVLP80YFFsxku6LODfcHkJ5tRvVbZubYPkbTe7kq1PLakbp73B
ofNE0VJw0gFmkOIPUnf+lYzpYLyx6v1Wb6Rqwb5d1NFaRdO/UN9XZJ64PY52daCT6xr+t4QiDMp2
PywPf3/D1Fl/IMguYTig9Z2KlG+1nxu9WvZ2D22IfZDL9ilZ3XZtDWmra+kgTWM2z/76yRYwf+RD
8V09yzIScw2MpwcRjXV0bV812Ut/3++Q0VuPCZbJ14N8EkewP4AM9FWSaiJQgIDA4xq+Vr0mPwv1
966pCJVjjOKHJIiKPTyIhoGnxnKA/5YaLbcEZUoA8sCJVVIYVBftzo0y9sNRxgt1CKIHNacNXhFQ
R1j9GpmKW9OwaNYhZ0U5B6S1iHyaV9ggUjxwkmsWLSIl5+BBB/6lsgoK5tznInFkho1dcg7H05uE
eDMIGYp91LcI6wJbVnvXgKryxD+1zF0O3+7gTVmgwbUcqCkYR/neWEADFsTXWfJW5AvBYUfLmV4I
dj+cLo0Lz+8EdIPqa5Bb1R+xsQwY/Bnp7+ily17TTHwgYg5YxyTGCq7eeKpmkgd7CcKnct1IBp6J
DeNEKIuQvNVPr9tf5eQAqLiMkI+4HMJUbcWtHwQaASu4bbrk+X5dktO3PKvDZNpvQELosQTduoII
/HoDzCJl0o8yM/TxO0r6CcK/0x53Jhni7AEI7ulIZT+eRhKMHBbbFx20zFhnMxks+UwCSid6lFiH
fKoKYRJG2K/07VUd4gAtfR9Nd+gF7bPZncldfq3xJ6wZ8kLQVj+EI00zxeEhYA+7nEaHBwg9IFS5
W2SZsgu/23T1hkw1/Fbhak/nHRuz4n2XFRbAVlPuGB5y0+AUO5n9gyB3nCU/kT0xVqzyL9NKzZS9
TfP5Gu1YqDMZHWW8NWCcdtWqLbfjCyDfeclEFssJlyQVL7JLpaol/vW5cagtIMW3234KNE0KrzoH
N1g1uJ+K0LElFLwM84pRkUkAyqtjm8NRi5FfYmTA7UrnZtlmBl7l+bjWqi0qPpyqKr6tnd3oR837
lJ9pDLYNxx/bLPy1SKMIJ+qZ78awt9jblAJAyLdzojzo/SezC9j6tQE9QMG342DuCBbrOcD5M7pn
MTz8pbAX0L5umXWTr33mPikzseChvYPvABgbsG5uWIellpIA4sVcN3WQoCRj++FZokcs6xE6r5wt
0d+TrBYRQ4X9smG4Uwq+3hD2/C6MbWTPtdI8016Qdx1d1nz++o8IuYKZqWGTgZAE+U/W6K/NLMMn
geXaVBUXZYt/9m8Xo6+7mao5WiKEpCX1etfeDxtgWLSaLIXnb69mjAdOSY+CR6tg6AAH8XpVSvzU
48Zl94aOJaR3d6MZxZkixbu55QDR5qKKKrPqq+Roa/3DUsayv4uuv8k9djA+NckkraKkZmLLL0DC
Ct8o1b4GIWrEaaxJBywWqmJK3E7F/C5Y8/32ArvFWTC2XI/6LExCyDr7Kd42pOpvgA8faoNWUjLv
O8NUA2xkOt8yC+xkoPLYVFwo73rVoVjdnZALTXy6QoJlHE9QHXEgdVC+bypL3G5VkbZQYNTxAEFt
9tJAjIikml8itNtSbT+ZElYjorvqWVU2kBD1vhBiGsslX+D02gb1BlctZWV/M0NfJimi8zr+v5jH
lWZha8/esYw6O1JtP2IW04KrOZDEY59sg/P/g8ETADdzERixsO7geXrynX0OEwnui2r2pGAcPO/X
VYJwbahStTJu1GjIdlZyw9lygim98/3NbqWQnerdVu0gwSZlM/XtZkSvglkzGOeMmHbWr7gd32l4
yeKZSk0LDnKoQPi6wN74rfAjUBgcv4kMpOfqwWPrz27SVTYwEx7QijCRy/coz7YJOSFdjSS+/Qej
ndDYynDYLZc7DnizFfUf5XEOFbNpVxdwrzuklXq+kz+C3dxiTCs1/u9jHP7gKh5wVoYYD4CG6NPv
wXu0Gkhv7ohN/6V7VZA7ThNRoT48nyMM+99WfA6tmkSmzAgYHba0RPBRastAZuN+mme+riNh39NX
AKzfrJLbR2XqSn3agqGneyajnbgx8CYHCHhuJBvgqahfq1rNHSy0BHwWaVu6yI655R7f7EQNUJBP
YwaeLV9fSHKfF8UZU1KXWGbrGvOBAvZwGPFt41wASP9v8gWu/Zaef1AyMm3BichKwRT6t2IrRIZe
kK/7ZfPUF+XXCV4D2AnQiPdJpK4f83pH9GzAhFtDxzShcJ87m3n8XKoxhrq3nJ7ceSmb+Ywt9tlt
/WATq0tKSwiRbFoBUJgcC0xR6GbrgHD0480sA1zss+g0LKFPeGTD28DOMaqy6+eNfOzSSGMm014t
NsImiDMptJIxDYTAe9qgBksZslT4GqGYrzp8O+gaOs/12yEK+l3GJoQw5OCalnZE4Zelq7Lf3dnh
O5S2Oua6tZfT75VDCeFZsv0ADmq3g9a1++xnHl/IdPQLvewdd/txwln3jyGyQP/4GGGi5Gvi4YBr
CNKbf4svAC7BP1pzt2HNM7O6lCL6BzU9q3SjPp1ftiIO1ZeFzvO6DGtuGNUaO+ZPYR/PrUHSzowA
Z5GBOGBYjaPLWt52pWNJYfxqcX5ObGnmdJdWsNqhwb6u5GvjeAO+rMinXOKaNejwzQM79/gmVduo
eCqkf/vrQdUsUOMX/777rkfQL7Y0cvWZRQfqOD9ArQktwnsND7cwzW29FvaR1g1xQca3zMREjUWg
osJ9NQCtgMCXoDsACDHKuUashFqaE5oAs0e5RPBlXr0kfqq5LnH/DZFpptlAQT9KGTxaZYAvE2hw
826EtLTyfhc0LoUrkzOOyq+pdE7QFUVnskOsVceOtZJbOiralD103vud9yh2QWmEXBbMOM/yHd6U
656X8+LjUz3826DzlXFYCrEJf4DtkM1U+gEMXYrLbudcGf2b76Rr9mlsTXCwMrYw04xw4D3gBkRd
5QHJ8ToD/uOq5feZKHTcGIDtIW0Q0cd+v96hwAxXKjXu1U3dwEez/UvcKw9p/u2MtLPIK+WKfJdY
W4UjOabMjqz1i5nmqnkmFL/ZgKiohM6oMAjynO8uxU6h200x3acCqrtRMb+3soCEE36ncvmTB2Ci
G5D/qgtOXQfIKXGmCOd/XAqj9T7Cv8dMvT0J4wY7HTYxiqMDjfGyZppPNRl3ZVbFlPTKcREPvujO
W/XeZ6UhSSq1dm3hsCrzQaN2H7mZ5kSPI1hbn20+2OzkM0a+gqkKcWmDHbkRgK9rBzdFUzBr1U4I
M7N7iIZLTG2U4uPFMvyokczGtdcgKy9cggjT5nVhWIYH0sVoCE9L3VRNSa4gO7d5ApJxIKsaade3
8R16s1cBCOu93ruH1JyxStrNpYNbOG/BE0wzDd54DyIXKlxWeklayAtlFKt6/+h0UOadtKgDSRSL
FmB081bvk40prB0X90CyXuJixzyQcbmnBVMnnQDBz8KvBbOmM2pY8Cs/qnfbRCHMnIaMRcfgsyse
ivLaxsuu9g9bAP3kkubdKmcpoWrunZlsVgiB8Go1HIlGtKYRO9Xjvud4acfXTmfzfo5tQDDPsiGF
o/JOg6sgj3R8T7wEP80xdXCcEar76AO1j/ZzRrpY+ogJArr2vR/WcTVLNg4az1jdcFotB6owrtmZ
XFUBSwSQJ3xGO7V7fCuVC4TG7hEjYr6SlyKnWalyTX1mgk+hDRA3rg8PNt/dNv1WDlRfp181Rumu
ViR5B3a/J+YFJQ8fogs1lRh6wDtOrFaGSG1LD+DdhoLfxNe+xWzyzXajVuG6HM+5ysFDJKMtZl7N
l28Q+0mJSXr5NhtBzahfxLhPMaTg4fAmXq1+U43ezfCB2FSidTSCawAsMM/nQAjWYTX9M/z5pt1K
Uuqyzyx5b55kwU1oyCuEBH1zEnN4MxRHMbj3nJ2TUXiQuerBVw1IH6iWjYPZ0Bdos+rUMjuX1d0O
MiNHmppqtN0BxvpHo0OGkmv7PQU9K/ywqDomIozfjAi56E3mdG/ISm/ZLNf6uWN+jWHuoLEnQWHn
IQMp7ZCwwwWpL89J5Z8YbM2Hhio54gw94mBP6gW4phJfuoN/2tGclKLLPZ5Fh3B6UFgk7nk/EFeZ
72Xnkip1T+eUeN5TsDL8nE5revrZx4aj7LxXgWhI53K5o/zGyW0IrDyxe5U9t8fyHRZtNznsO+8r
Ap+6xmFf7cUgov6t7CcuXadMspe1oHJ8+hd7pT+yvJrMIHZhFfj9RD8KETBUerh5C1O7ZMqHhmYM
lI1x9XRGG+AMV0cd7bcFJGFbRuUO/DgHvktuI+TgEbPqcna8aZF1SNGKlKAkSQ6U3i71dn9z7Pzk
1VbWsdwzfxvFgQA4E0/CmuoiLs+lTzTUb6aupPtlfGOtwLB3jSkwMKvBkJ6t+Rsw+lEyA4OHU7gV
5Y7XVmBLRYXW5j3JcNJw7sG3zmQeo+pFnL7wPnrpKBRyDW3IG6eUpNG7JdbXDGZnMfzc40QSlCcD
b7jamLLykerQ2scWlpckuSjLlpo8T/lPAxvYjb9MlO1E79MFpysT+kbzUzKBJGwmopnHnbd3lcHs
GFPRsgh2Ap+3W2Q/9r3S8YcOBeHGDqTcxgpFe8OxkXwGJVSLsX8qy3QJKCOiqXqQwZ1+JT+5nHT7
jdepp24rKicjiO+78/IemBkeZ1QW2wRhFkChOOUlJrAAAu7gKrLaYggnRKRDfI8cM67qkmrbg5Zu
R2Y4iN41rL+SAsJzcWe4NuyQBUX0kiczHrJgxxf0Rv+p1PDkWYv8ZG4LxozgHzSO3OmsdK1gJ204
w5wgcejYBpgQjiW1v/9hi+hBYxm8bJzTCj89lpBtidUprQUMp5vQJDNXzn/fceWQou0LAZvD6IHm
0psK/SGHhxIq3kdh1s4RZi+K3fFnn8fxTB7g0Cg2xfrXXalKcqWhN1Nz2SajgubVXmkvo+Zywfrv
IYJNU1O0U7EVksMGVQGu6DoBvp8ztr0lMSObn1xcr+ZGJQ6ngNSMx34+h4zKqhHSNsvPwFYUqbQR
jBvcQfeeXFsH71ii09tdEpSUHTtRffAVvsd000adPcBfpPr77/NQVDOOmjugV9N0/DcSah322nfK
CnY4seGvlat2RtaJa0NofdHdHSHvUulkySnGIOjLVMoh2OTWel/uCtjrcqRgMVjJFWj8E51h/jME
kx15f3sE8MUEyE0pX3KvJML7YQHzXwIrgbcrSjI1x6vTY4HWpfoxZlAoDtqikB6pBfwKbFa24GTz
Myaea+422pMtYxN/hEmwDV6XZBI1K0bU4RTIQcjrWJTT+oXozlwMnvHp74SF13Pv+6tTamKldjnH
yGKotjUkxO6v9qHtCrhyteABT2/S8MyhuM5XZ1QyyEhHToU6vCfbtvmtCdgfM+uQ+pXuf0Nx4qqL
V8au/yB2GKbN4iZZtmqxHByrsDwhHopSdZR5ub9vLIry6B8NtDzmgAnD64LA+xbvleUK7AilVxxy
N3cCrwyo2yL5AwlM+4NPsaEaTm+4ap34sObUcOwNLZXi3ddagdcuAK8e7mrTyTCxrdY+9zvLX0wz
Sd5MNzHzYPRSksVMSVlzxveVVPBrh4kI8+WS1OTt7wwdELzitdHJMJCcMErug2hci/wRH27eJY+H
JhHtucTV1yOOZAGQYWYkqHUdzGABrY+nE2f4GnW3RED82if3ixLhNfr6N8spG5dNr2ASDI+RcGOf
7Bvl9nvrgvlTMMzifCoJ5zXAv2gXZke91rJWDOLhalFT+KPn2n26LALNWl/ll7aHAIwEPyvtYZtW
uKgPlBBXg/P6YAonpKc5LN1hibHGt4w57RcWyUP+SV2MuMN8RHb/67aSh5TppXXACbmQYQVgCtfE
b7jn0xrG8UBAdN2ER23j/umK4j65sySx6hYa0TeGW51+wlVmS9FRdQhLHgTVq/BJ+TjNaLSt+nFW
DMu9fVY4kL9vlrvPdp3HTo3z7oCZjJs8G20xhk2CR2rmJa3jX7JO2wHEFD/C9zRtRgXRaNIIhmk3
wloRsr6JYkYda/9Oxccnxmmw6I5jhuGjzeZJi+hBIkronr91/AM7nFTQBo9ZZ8NW6uvoGvAoJN6d
I5FPFV66yBidGOTjPGwyST+wVGgzS7tg38pfy8X0u/MIv7z21DHgOycaryM4PL3a4bs1f/ieAWQk
iG8+ESl5Pz1ckcCmxXgr8+hPkgU3hokN2DTBvHWyNDZ7Dq63c0FxsgrGAMwxlzWkpug6Igo9TzCe
UlLluLOD142TvGw9hnKV0jF3bWzUZNnEH2RSLRTTW+o7R0uUzjHbS4z2o5T8YAilGWByDV9ceEFA
5VLMyGWV3gkswpVwzX6GElTn6B9IeQSbns/Zpe9TVwSlB3PhuE91hNDhaTWEuhRcqZp7a3FK2/LS
SYpaV511Q5u1rKFAFBkfq+zyxQioup4HtvxUXSZQmnijB2/2Q6jSqa71Wql8ln54cVVOe5wR4fmy
j6Z3CoCJBb3hSenX8o1HaUMIh2VVfKhfolxz0MzZiHk4M/yBW7KwEcPgsXvCrc/DSNgk04NULf1w
NfgYTSEjnRyOMXtJy0wkzesWxqpRKGRYYwy/yQ6Dn01UpeIIV3lv6SEgO8pvDcdHBEz9G1ra4iGz
WBga45sMFIMwopEUi27Ih2xGJKQ89fohXfpWGRVqi87H/5ZiQw9HX2Ui3sNyiw2tgcE0hF/KqLCZ
a85OJVy80r7zPmMthF7O3s1E1vVCHDF5p7KnZeMKyZIAhFQmDf+RYDYTffdVukzeow3mrDDwNUxZ
ktyMFrBlRXcCzOkVprJ/gyGdKeRpOnhZXD5FolCjUMk3HuqLS+flUU3uEBy3D5ilC8XpUqyXdPhB
L2qsjTRAqU8ShlE3TojsOahmEWLefIQ67u7yljMLWw0jeVmdDde+gSUH+SzBGLncXlVdwW67CEJR
rhbPXNx7fc6Z2/xEJP1fxABKtdKG8YdkT0Yl3b8Fx52hD0BBP0G3heKTyRfb4Tzxf5VvjMfsfH2v
QY52WjdeDd1XoYT3Z6MWvGDaVWGdD7fpcPwKDpZ287lbayV58UxymoCpGJl0l6Ss34uHZ/46yLNM
GG+E+uL7CT1Z4/TD0Y6U1au2xcHgdtpqbqaYpLntCywQRF8MRAwaC7nxNgka8q6TWYuXKJnBuz93
r2HR2NztEnhFtDhh8gXFs4NC4MI0J6ZyJA+DjgOXJFdliveXe35cQR+14semBbsYQ//OVCL2jc12
p+5IX1VM97rtX/OEaqip7QKNrMkDXg6NZEvT7oCVd9vY6NnVS4I55hKWZcQ3HplwMJHSxmm8i760
IV8Xa6BKuKH+f3YwiHgEBiz4FLpGeMIVlY3rQF0tQQUu2h5V8JV+VZhFMWayGd6/LXo4O5TzJ5Ue
MrmVUJDPK5zS0O6m6RRxwp4toQ3oKNFfzr0WSoNgGXTpw35mpqRnxLeiBxl50+IhGuJjJj7/2qNq
mHf1FiayY1HqXbrbxxLdV2Sx+zucuTffvLXIUynLYfpe4TKINB0Eb8U7ydsqXvO6A8VNhuuHl7ft
IqC45maNn/1G6Ppq5xdeCOlR5iJENnLnFihggfnTNG1jaywVGjyk2d9a7vCsaBglj+/wWHbPAw0u
65MRVMBMZtNDLjsNreSCGglELNHtVyfD6pqHzqG/mq1uztsouvOGojqQJX05AllOJoHQl/6g+cQ6
q7D6A0Xv0uO0r1bXB/8ZusWmSBSoG+igdH0xchSDLw0kpCZOZZiMixooJSBcJ8LvNTLGVQ1FqrRo
6SmNQFsE1vEMo6bCo3xfn5sTV2BrtLOhw4bEcynnKmPtAwAYqka+1QjFTIxXtb68bTbi3k22DyeD
Mc0rq9rCMZ98xjxb9rXupts4kZZriPzKEYQolKSbCvNIGZo4RQHzlbf7VqPuOMi3ZprK4+bkrNxk
04rwJUI8cWQyHXQjZNbgHiZSLaIBKFntfPIU7367azGjGwnuSTzt8FWLc7DVJvPAwlYsthvY6NKn
dqctQnNYc7se0tOHqey7YUQyN0pOLPKcCTsa0ZyEzDvgniLhX2AfDYk7DYmncJdt8i9ZN3rGlLW5
lc7xaX0vDAL1JNo23t/EBMqf2g39U8mZOCkwBPBTXc3MRiwyxfTyEnIEXEKl92lYSWx2/Gft5yAm
sfwTgoIoXX8CVg2oE6gG7pY0mOd9xrCkvwRiMvGv8TqHswkjtxtv5kQT2jG+N8jwM+f043o1g/Cj
+yosaUXorrDmMswrem6olUGxfKZZj54z0ZKY1MO0ENh3zuVUZbtCo6p2eEsyUBYRGHmXjWnMQuPK
HmFZDsRLSjiy7MOhWNpsoigK/9sgAC3alpQplca3lECt0rA3ETIvOzO+XcIl1Wuev1rb7MW0Zktl
2dE3ru0aw3NV0e+VNCB67i8MRruoLZQA8eAq9OllkeirOKDRsMB8VT7bQvTVi8GqQDu/7RYP0T1I
tHGt+ZRAJbH84TDPYVcxxTdot8vgRJwiqrDJLBjZCW/cX6lBJemheATB/2eCwusGLoSna1I3XgSR
J8b3qZ4eXetxaPaSPqECvQKfbRMrDu6VK+ez7afF+T/q4nZry+w6YPVkQB0LnJAoqlGRmNh5gYw7
Y9lYfv/+IybLDGwVqGtouYD55wBB1dQhzeRH5zbNFRRqBD4I0wjNCTlO+sUbGqSOCLo6qGCl90Rc
HpaggZ2yjsl/NjAxl1T8/tF79j5ZMz9o8LvmxiRlK+bfRsp+Qho346XiO5QuHnqU+NYkKcfft8SR
vYePnxhol/WK61t09yY5p8AaE3OyRyTlfuRH/6iK65xl3KWkMWehs4wq4JdM1Se3Xc4n0CMNgi8D
j3jx4oazuhx4m+66gch5Ube6hnRbN5fnkMldTuXJnKBZ1WUA7bUMrQCFR65cmlPFdBSMDmvaTG+i
EUK/GUSy81Keji6XFng/vy1RTyPTNNjN0HTarZmzBhuiXcPTFsiGJAJnkVbhKzksbGRTtDAFUs5d
cb3cBRevJVYSjEP+d7i8DWekFOdTJtmE/Zqi5wPRqRmCa6m5CNN21m1T8iuXjFRxU9s3F6nlYk7c
W4TgYt+5ysAyV/VmIhBP8lLh0+Xrnmm2FK1nwgeHqh6YlAYQut7LIz5Bg4aZk34oIm/fKd8rM561
YJfgya7RZbtt2bSuorNfjluw37dzFbhMo9XjDdg32K8kiOc3vJEwwY54KFmuqkM/b5J4Pv4RXBEn
rG/xInwaV8Clp/Ko7oHnMoZPq8Mm+LXlOTTX3ekwWhJ/E7c3hPatUKj0wdviCFADQVCqAiQCbZAn
99IfVsEjy2SK5HAt3lHXlbI6a0S3UpWB/ErrjRoXIKLzNx5w/JCMHLQk+7qCFuPdUCJTyRUoOWfA
gEgIm+ev0oFkzVntTTupUdu50lNyCqFGCfeSoIok0iNm5IP/sb2dTOKZlCFja3SNP5bL0VEysd4w
0IQ0h1pFQPGmNrnhYEZcLkCUr3S0JBKOJlOZyi4wIycXwcVy/STWLmm6LD8SJQnDnUEEl7bKyCiF
CiFhHEt0i4mJhPWmWjivq3nhgF/XDwyqwvuJ9zNqjM2XNiiWYQYNHgSQIQavy/jb/BVJHefWZ3DQ
FVN8R+jgJ80HF6C4eC+OaV/PyJbm0kSbHfReqxRoO1P303XSS50dYWfnguMBlTet9fitm8vxqpmo
qL8xORt5kk8SKGrqqxJo/DY0ULf4SDr6XFo03SnaewskGC+XXXDg20nE9fUDH0E6QGUyKyoJzNAD
/nbQIbdQUOV9HuevybNXbz0ppjt/PYDs6Q6pBFEpCzif6rYZUVuWtYyChOs5WXJvyP48me4gSiay
549Pu4xDihYoXLAQi7xmdWdrAVRWU7z4asuy4JEYtT5bn3aXoiYjnwjlJ0bOMV170qK9UJfhWStp
0KvbxWIZsFKKkKqFR1Z573+hJvAeBoLCx2kidflhjKaaWFfqGihK6lW95noS9SxzRFOp15J4h5I5
osKFszzhgCG48gOUPDhQBBkl/HSa8AFEwDmI26xAnW8CgWSwILNHW6s8vZZi/5K5JPWQYEs4pCsi
n3u9Ipzn8VtyR/hb88/1RgAuCSKBxJpghcllWt6OzKIHteGQeSH0uGHJNxLf8tHhWy/FWsTkTaDu
c/2oNu4ZZiVEsyRMe43JBZh2beYCt+EiVNYMMUJzj8ismmT2qDrBe5Pq8qyZwfAv2hq2L+KV0tHo
CtD6e0UW3+7YvAp69AfexMUAUI951iJlS/r33WGWBvTyCh88FyFPW/o/tRL+BCGQB1W18ACgs/GZ
BBz8Wm6rxa04eb4Cb1PzbPXZjmBZdQjAbE/L54zXYgSfHmO1hlCgnYLE2Rp+Oe6WTW6caDub2jFI
Z5O4B1kcSyd6qGPyBbAXi3PEXijnL3jN/uhZ6Il3YM6I5jW2wl2M0nIbBRSk/K/ff+o9Q/lzYOsE
arToSbNiNRmTa5k8mmhtM7ZR4bd7BO71qjnSAaacVRjhtifdkSJ6qCosFJoY2fmxcBz69KzmzRI7
fhXC2nW8QrU0AswkheqO9+BXUMkMRtOJ4MgfWNTX4aQgYWDEkEs0Jwr+JgiwwJU8Yao9QtapcxsQ
hfCubvBzObyl1CD7s6lL4iGYLeVqcqf1GW4U4OYcryeGmoh8Gh5f8AHSklTkqUUNC6+8igIbHN25
AhIrZQL4e2Uh67ThMk/xxM2PCWy6QCF0XeJCrjl3XmcaXTetB3K+JvigtdRBZOZ2DMDuUgVCtJBf
FSXQ9GYNA3woQU53GUab6IbpKPqFMJY/AY+r3sPoFiQ2rvbKySOIymhLg2rYd0slNzG1ONjcR7ou
9dHuyZWYRi1Y7RIcfZcFe8E/0ovMXGyWWc56fwlCkSjHAtMsuKwxmtrygJ3z14nTxTozlvO4a5Tv
iVC9yuOdETlrgB+VpgzwzG1vUZItY74hzDhrur98ZrvOf5BwZwR54qxhHvhYK0lEm8Bme2NrhCZ8
Ir+Sb2QHjPLVm6BKDTQiAY/j+APdajKisxBYlLWd7bWK7r1GQbleMceSqgtLz6lnH3Xzvu8oIgs9
TSHT55PQMSASeV1i+XmffBt7rmZgbhfgQ2jQ0LSmaXwZH8ElnnBLsqYv3d9d8KyiU8WUZ1j67Mbj
V8ROHsRldhYRt3wko2XJDcg/Ymch+KNEJa0Gr/t6dVcgbm9SFAKcIh97GF9B4rX7Mo6Yb7Cmhlmw
VHDbtVjFyrA76RAE2sz0ScMzeI6EbpCBuGOPCkATA641lSrG/yAjgrftsWMOPfSvVdLpJLEDndC4
sxp4fCqD4dDL+9FKJWFXHXwu3E6bsdeDJ0dk4HE4xrQSl7MmhP0ZeSsOQ4NBdHHbOToQQ5UdsRzZ
nNmSkVv+1y8gjzHhQBeeVrkOl2CCDJ1x88pw84LKmjgcfOZujRWzmDNtJNLg8qLRcVs1E9PSVXV6
C/8/TVD3pF+Wj4Wp6VByGI6c/p3ufq4ydd92fM84R/6B9p1KHKoicuPMT4W82ZIa0Gf2hnOpJesF
dlw6ty+VOvDo67OqRzPRtiFNNOuuwdWUnSpajychr4i8wifPKk/3nMMRP2JKrDfpr51AHckKYYCP
+AQJFx9KnUxl7pPzRCZuUv/gIGScCFwawFCKEXhYhLPh/vdv/VQN94cAiPAxMCUtHhYEPZozDL8s
3ve2KfiX2uW7mLOkTL5xdXgEpTPbXX35dvZsObXJfUd/2s5Z7pqx/yecfgMJfzdrbhMUTAq6Rmpw
oiipMcLArCRNSJhY81Fwml5Oqpazi9BkUZQ3AWOa3KW3NREGRUcC5hU9RtOKGx3XgOb9VWNKezjd
/yqH7tYLxivsgbn/zfeXdgSAeaIX2mw7FBdOXfK/2ESicuLa6MWkeh5qYboSVd0RYwhWlgPGe+RN
/8R7ud/aeOeP0/M8oYSXg5QXVDnvClF+tzDQxlucGttIm1GOzVFvSbjEwXT81Bv5sE33SmABlq4l
SHpMIUaxmpEo7HbMJ6GPubGD6Dj52EPwC90XRC4DrcGsQPEwIbdsrPGtHWtlr6CMPu2tUOyVaj7X
dZwC1P4UlLMdGjoNFFajNQrElFjkAQ4ZwiPVjNREOWHw6rtC0vt0m8FTq0C1tMBFGxdMbZSug69w
Ov09C+6+hZ9JzoUI8MYRYt0k2OE9YYMIWiuknZwwqgwOI5zgdgvyWq6VdhdqJ33FYwrpwBHWrGiM
AKXEijkAQwbM/L7qaG+5iv9YPAotw5Yd6rVvEW7xvEbajcGBiVVcMN6GY6Yj1XbneUna2ER0sR9V
RKuWNZLG3oTqezedexw27KkoXW+ikX/mOZpzUcoOofEhm0pEVXb4THJz/hdyYNyDRnnKvi9OEeih
fOGyWvx0LkctG9g1pZMW8uNLRy+VEyZfXcY03InUa4MMzNhI5OH5iYNjE5do1dA0ke6uY43Sau+B
p2wVuS2kweHn5Foytrt5Vsfa8U55CkjPwxWk29H3Cstf+t6b20O228Ph6pcPTs7UMxOHNNmKMij9
HsOoV4vO6ZERGFT6aevWzn5jDPxRR3zlTt4WpRKLvRrVhzlGQHfnF9M/C7mfbOwb4PpLA9lK3O0g
SaoyXF6rd+UhFiMkIZ85EzUmPXvj4owh+ldAzO3ovc4r012tUL96zqn99bxVyRzaI9ujRjwBjFEA
yUD52dO4g/vYLAmitH0DtfNya6gX1trOmKpYg0yIxUdWFe+VFqKqc36hrKqzxn90vQX2MdZdt/0Q
W6N4SpwvdSxJF1Ho5zsrgsv2GwLClHpAB+Ag3ACWozW8yKfuSNoKe+BHV6rfr5dy1dFv1w4EhJ90
TMiRVsLi+0VGc8CswMzsOeY2SAjPrT6pzNrvUhNpG1ajzjs5ERbYjd8kNIE49F2YRpKdaQ9888/Q
fzSk+2t0EtS1q61FYcWI2vorHJ9DTb3J+tPQmkOfXUny5RwE88Z78oyyPbebkeSbIBVPiHuJedHf
Cv4lUgeYB2qr8XduNWUbItCuWWbY5lwuEDJq2eSUDEc2RhNMQ8Tpf76nL9tzN71ysWMatTZuZFDr
8DiWOLguD/R8czQrcjXjHAagKeJuCHo2KuHVWGZFjfoF6Tb9KfVrm7jJMg+bWQZCxEzhj/zOvbnL
PpJiIE5clBD+4hAXfa9tLtjGox4DEYnX2BIiG+DWXLVJHtnKgQshndwdosLeFrBOhHBzTYqCqDeT
T1ra7CWdBcEQiaY6FFIy8n9JgtTKkT8TXNDqzCbKVaNDMI9tVmUU1AjyKtf3ZABl4pGUJ8lEedLu
Nd8VX49E/kGQbjVSaH7dq51fe0XZgVrssQTeWE7QrYMQEGUzI3wzOt4AZIjYjqmjQ6qUEyacEdrL
Oyylp4wZGGbjU0P1qkIiz8hF05MimDpBl86oictMbWarePSJSyu8MA+h44UeleiNc7v+mT81LL4v
n6HcPCkqnjr2ha7LkTCyhPxMTXgRRJD2pCtaYT6n9woE33We0IDn0sRBBYskmRD6W9fE22xAbv/E
2CDe3Fzu4WRLyAMA2++C6snxWqfvaEWKzkgyMfkMA6tI+/76JWXeBefTrTeS5OaxGpHv0gacwtss
1Ek8pR5I+1vVvAblt649NhW+Tt4KfLD7UQqnIZKuPG1TrwzqzJtmZbqjH/IYR5AOpwjv1D4o3qrY
7vu6FK/17hE8H8rNGAaug2PudXphjJDQGHFLxdg63nLYGmJVZX5Qq5h2BQCu5zJbV2A5nBJOKVZ2
kqZ4SliLKHQ3xgeNIbldjEw1bWXs9+XbQ5jFn7ERDh6U9pFU5ZaBqD0RwtmfDkalm0NyP77mcjZ6
M7aEP9lNm06RzGACttfUmuMYP1uTxvog+Gcxy3kTOcS5ULiR6nyIowyIwK6QvA1fZlhoriqDS8Wq
IGxSQkY3hflMIwpvoNlifDAPEQqqCGk+XT72MKmXgV91Tvh49UKaMe4xjPWf32N6Bs1R/AIBTkfK
cg8R3ooD/ItDCu4NYBbibv+e/vzT0iqXg9YdPUuXG0x/N5VQl+PWkkkl8DUjGP2yN2sCmpUWY+47
khN2TSj5z8+Qc7pvN5YsZrITWIunn47Tm7UrIaPleGLXS5jqGnyZdCOlgxlHxt+9umwFJPGZTlHd
LP7IrDFApZMDYEtYECJcjnvJXzNgYjeKg9j3qmiVcGx3tVDbIGhOszXsQwz59P2IfSz+Ffo4qrc+
dPZ03osUi+xmWd98LoQ0ezzv5zT7qRWk7vcRqeIfKyBtxHbsqS4jTId/Athyxf0nBV6GJ3aPEKnC
E6DNIkrf6wN5VkMc/4zg78LGg1Ol9NO07pnnOucDkqXTOJgBkIWLWeHntwOMWnUC2jVfSgSaOhc5
QyGWVM4GYMJz211AyGNrSvg3InTaJM/mU2b6Rej52clUgrLAL11VXd436dwLpO1wxA4RE1CvatWl
TcZobmZQt4M+hKuuIQGsXv0bLj6dliudXKc9hDiuN1hHg3RAwV9Hjk0VQCaZAUwa2uPkVRJgJfTd
VFDN735dxiJgtuAc9jHjywmHspoxIfmXJm/0LucDXuFfUdJm1kzRoYvqas/N/AF62nOTlackO6EU
mY4+awlZ/dktcgrPt6eN9RYRRn5BqIxIhzqVoVd0jRvvvxHzZylaOMy2jzlz6+cEj441HCXmksJ/
nxwiwk2xwe5u7DdidLIfOicN+Jta3sWG2Zf/P/MQGwGa9FKxKyGyoBmuqhgD4LeNXpsA9K8GQTq3
KLhmEpzL0mej7BUPj7NKKRszqyGN0qyQLvR7w9R2FSAqXsHLxjF3WP2Mu+Z3Ro+Bq1uKsROEUPM/
6Cq56WY/PI/C7DObW1yyikx4OqektRIkqxBLRfcIV7YDTXZeoPSlp3ERTT+GQE4ZojInfiYL8CTl
ysZbw43R642t9wL/FprxzvTcHEFvlk7U7onlM/sr6rIcmL73/M1I/QZEnMjNgupNXNMPYfDDrArn
/P4Ltc+wpJ/w8xmCPT1TNrFo5bnQ1O4Ph16YbNJ4NbxaiMyOHTaLdzADLwuU+a7vRrqMuB25bhNp
oG5w3YoEas8a8dKHUWDWrtFAJn/xvM2TlcL3EKCs1UxVhCSW3bD28N1coTDcBRdgHTv6m1L21SKT
tCeDriOctx6yJq/iFiLbAOvqvebkJJAN6F8jXu8CpRXTpqQN7GFpL9r3lH9V5EdKCtjO/QlqznZp
FcDkvNFN3DFSbo3MxAW+3A6WKEhewpGwhezDY3Mzu4ClZbZFq59/oFfJrBQaRTiGu2577MXHuaiI
XSCXtV7CSyiY7mjIiVn8dNZpC/miqZd1UqgCHJVyHd6sFVzYI0Joifu2FcNYhjgk+n2FNHJROGwT
ZShDogGp34Ig6UfHK5M+5TvM+W3DqODxcJEAeq9xHNzLPp9nSEkCofoQC7EkiyloH30ZEj1nrv5C
DC1iXDmEQAJtAZcoe3Fu1HVp5mvXIfckxm68pDrggewPPLA5dBHoKGkXGmOLgg7yqiPNUiv2L4g2
VxxwerQ8vYbzHKNyehzNkSHpQei9MVrhJJ+QDGcTRsvk8eJs/T5RD2EU6VbSmdB1RwFCu/LRqlvq
3Dpfayjm9KpP57fLJJiDcoGvPd1BwVJkuAU8Cv28XCfAzAHKzEkl06dnlY56GxOP5Crcv50alI4J
HL3FN0ir0xJXoTGlVZKjWXdk/mReEoSTGrmKMwbHEhkmVaiFgOLVKR5rAQZGJDC3XltDCu8YdH5I
YCbDC7B4U9pf/mzfSPTgmhJu6cYHm4AFXeAkeI4bKSfzcg8eSguZceK44cb8WorKbhVhBaqZyftW
G6MMZ0NfLvb8Ikh2svDjy0H6EsaSo/gqoMkQtcT3wCWido5VnAM2wQ/QtTdcFvx3650qO8iJicUf
m4z6vt0q5RuQ+TmmhzGs0u5Wk3zgpHo5J9pLjBseMYQtqXhQ0KgS0qxSeAFuHtYqoKGRpIY+hNNC
OonZ2fyQcw6g4p6EeQwo60kodEMG3V6Ea0RcW6gWVHU2z6+GNsKtrWm0Fv2Nv6jc4YqG4qzLl9CK
tuW79w3wnYSqso2YN6vjiSiOb/KD1i6zYjKy4jE2Wlgx4WoevP2LZ8HtEWMwgB3OP0TDG2WPfH+u
d8BWRL3ykO0qv0t4mAwxfWEMXjwo0v4MjcCkYSc6fuS3f8/RqfJfaZ0EurZ9Ny3Kxb9NY4o6B5sl
wZhb+ySwga0g0oryIBB8pHqpPEqYlRLIRJLvRMx9Qx2sYwvBRHERcG4IiMOiX9A7K5Wc3jI1EMLr
7dxhSg8oi1UrZW5jQv7zj5elGQ/rB7DFjqu15dLNeRof1ORn8LQMxUcI9SloouOhlb83aUedhqgm
g8Tg9MeonzasHucqcYknVuH0Pclvm2JAo65DHyogvxGLW4l1fBHl89eA1AuOZuLH5mzaCjiZ4GqD
Pu4AV844IvzQl4xQZwWQbzpZQ11WkfONxzpCCQ1ZckjRRObvBHt5m+lbDMgXOYX0Y4d1kYp4Euah
5UG1i+lbW3VzYqy1tny7Oa6VU1I+8eAvTVG7VWbiYyhGuwtPgGx2595GQVd78yKG9KauE1f3vlil
jEIcElVJD3c9RrTGw25zke6N2alg84nZr4C2rUKpuWhe0r4Sju8oHjjZrw//pMjiHRUKUAuAM5TK
KLQSgEaXyZvK8lcb6kRdv88s+NXFQP74A5oZM05w6kzwZEGLDXc1qYaDea9bKUTHEzuEIVHw3fWa
rJVwBHp0yd2filQ7bQaGYaDrTw4TKOTwmvZc8uZXvjRHaWMZklv1MaSiWsRL5UuEjUrFDZAt7Gh/
uCsOXK/UfHcEvJgsquwI2BO8cQF8Af4PE8O8L/u+BrG7k48kkaP0IhIq2JDrUpj9aA59VUIYgIRg
kPlUPuCnlMI6O8ZmU7BgdGOcgIYpezVmF8tw5Qsdg6WjA5WeY5HATmv2m42TMnlDXNRVq7j9ncOU
e29aQfZY/dHq7T2a9BmtaMgdZUYiR2KYsB6zj6uN075QrNeUVfa9ta1XcBnQ7iXpnIRXYOW2eldL
XvfXbBdd9k5GcpWn1qpe5yhxgCVy5q1Mc+EeCpoh3CMNvN1VEHXbTqS5nfloxhl7X5LEJGUuQWAE
sQo/QBcTrKG+Z7noG/tRYAh6qpH1l6nuV5GX/JI3KSrmoCvf8BQx+aPaKqI3jYG8eYLn48CN2dNJ
S2GRrOkKgD/cNh+rnCVCRlHhj2c2Pl3KXXIPjUA2CCmpF+WhfNw3/rnQqnNByiX5E6Co15u2RW3m
nhfdIvaZG88cOU7FVGnmvOrosErCqWpnwc6oF8R1+Mnq5HYe1/YkbazDwQAyP13OMGL9a4FYtzXV
lWbdMAtXmCSIfn+anw1HMHGO2Cok4YRfDW6Dc5dQxAaebYWfR0hFzjRuqA+G3pMW5tQIPaIHrdIB
8zmgYZuLUq1/y0JNb8ub8Hc9CL5KmVpCxD4MGGNAfbAx3tLdUISxNZvCvAxknNNE4J/L2XCXUlwl
BZ1DnGmLt69WSbno4Z1L2+yJwaxm0mybA0l/UXsb/TdtcdNbLCjjHhnRq/tKbZMNrDF68/ZIUdvO
RzQ8jb5I2SezQyEA+nPhOnf/3bhxBVtPud52KZgYxRbBHWyG3oTJoR4AaOM88KCEv3huVa0I3jXB
hKN8ltvqrrRSGaOv138OqKK75eFWwZLZX2X74Wc1Jt1awYTKmvfYfiYyhI/YTj+kQjJpXjF8Ub9w
rUdbYxz6sG9M+/PgAs9tM9/jM7WyWE8lDa/fjA4aXJBYMsKoVxH5Pi5UY7TNinVpzhVOeEhXH/Lt
z5doOR2Pgih6Yto4WyxGVRPX6nBt07riVjWskTxhGiDut14s/CHUGCvms3aoXHKNdinPxm8ilrK2
ZZebUeA0IZr+dIjkQ0OnU7AWpz5cvsNAnfKUkgftVz6xxptXe+K5USeCioxgFd1ZgEOeIPXeVRH1
/GvYD2tzTpodo0M2om52GU28h/ILCJsR/0vZQX3jg5IarvdbDFJbcfw+A5x+pZRBP38WmAvPw07b
WvUXGpOPjz4hOmTb8Ye2XkFPMzyCj7d7YR7pCZVKW0xZZrjj2KA2iNIRhMvR4DNsYtMbrelV9NBd
0K6oFTH1hmoNRVNBKFmMpHx9fFDCp90lrbUPR51A9dsX/uM1MRUG/qGSKb51C2xY6ig0P9f3kc7k
XMa9qPvPi3Aheto4Mo8nVEEJUTI/UiUsGEVKQvZHw7vHfoeCLgOTuAIiL8k1/xKwvvbimg+Hxdh/
uqO0uT1yzpBSrj4RZiUla08zXw3OdV/hqHKXWyhtnN2IWAji1TFTew9lsi2dwiC/8kWHPcv1McU7
OnHVTQJYmV+icqM1oqmrXs5/eWNeM12kDPTgYvqddgGfOwiCp3t14IxFq2SzQ8m6RF/kopYlGu3j
N/Z6BqV5428m24iN4tcwN5YAno2cfm4FX4p/2kzfrEfH9DYN8/mCDzUNjLCUQm+4rLu0KqCSrDTB
rCmkHlNNw2nq40VB9mAtny4KlUrR4xlEVKF3RVTkRjAmbdvr3EQnTIVG5D+MqSCkVfcaSV7H+sGT
VGb4I6DOGn1nNTfVGx8MbQ7welteV203D/9hhMk5LK919al2fL3MLqjPCmOh8I91eHCuVDWtIMDD
S6CPotNgO222w/ez2ZAlT2L1bW8KOMPW2GyPw6uocpa341dWo543IErEqoJ0ZbqhpGKq17upo7sh
jv5T0ur5Us3AVQSjVyQmvvzlYVk4CtHgsdorT9wPH+x4nsf9Vk/4x0vppowPF7RBShANA7KjDxWx
b6YE4yAnVzfN95WbFHtltQPaqSLJHOy2EVjWitwPJlVc8ZkBU6ELdOQPjqaaFOEw1S4QKCy36X+g
JrBic3CyVpgF1hq/gPO6yQKpsbUC5goapfaUV1C73I/27gbYDaS3oOT/jbdhf56DxUJ85fzsXdU8
YCZHOjfMlyaqMZi5s3TkJz9D9mBuk+43RPnOpwJV9lgI+5z6YL9DoqvyEoDRcevIhEpU9Ytkf/4R
asGk/lDTjgI3GyCmXLHR2RNWfLx22mvrBYrUII7/6DwEP7dOxVKRz1nxONOnsguED0r0KujJi6wW
K8gZc7u9K8dA9LbS2i1rRFk4lPlk3XAEWAof9a+uaeC7HcjTD0QtVMcWeGWPGj8OMm5kZ9i4wesI
cpSrMo0JmauSSQxsxvh9Ysfn91ztNWikM8NKGyZSmkGB4kaXm0JHtG3VS5SKSw00vxnJpUksDUYe
+Qv3FMWVHXiuXI34wUBxVK2aiLsxi+LwMSnbmdm3qxktDOcPgHQrhTMoGkzm+FrXJryKVA750dwQ
Vgioj1ODt8jr3cyOtxjFP8hNloeEfEYuvWfLQ8OLLkC1A5Sc1R75NGs6F+Cijq5as6oUxqb6VTiI
f91OKoqYJJGMyaD8rbHHP2Rj9o9ESunQM5GkpHU3SqdCi/8opJBWX+ACSFfX6xEuSJDNp7UMsjtm
uGMrQaAV/WPD1QaS9I9ggvHRKvWPKH9U6N6fwF10o3Vh+7rBQdas/vFWHDWu3MVX1oEmRu5P/qK9
uT29egUoxNipnhR8NR52YIwzfZLGAZcAHJafGk6wJN6+QfbCbxO+C684XRXO13wUpLTFRWBVzyo1
OWW8/sUupxrQWtNg0MwH/Jrof+/EPWZIZnyc8+7pxjBjkdIxkx0+iSlaLTduq6UJZPQhVgL3URzZ
mAOiwOVGKvfQHpH5rs+i21XE6USkjfTHTFsZpx/lMhV4e7pEei/s2t4a2KHWJhogmY5AETgAEEav
86/tmrcoU5uNdurWba3meCjq4FMSXA2bbfjgTiSXlIEtHxj1i0wn3a+0u2ABFyeNR66TanPa2Sy3
fGRsjn701b2oQwyCSKUOhPh/msO/8bdrodKZU0ngOcfkhl+r2oxtU+OznQTYlRGJV1OykF0+thFC
0Mfm6BH5rYEdLOVrmVftTjpq9iuv5ewy+OwJlXz0XCEyVew23ZkvSO2MsiwYWW9OTXmUm9m8xbDZ
XLiHgD5scWt47h5MB8IehCB9unp/QAEfGWLockMVvI9UMRUEivW/AyUN2nfeC+jMBrtWU9rVLVrk
Z7z5gfuJsykruGOM86XX3Wd30B6c2fAGxNIIxUfShexikTaiXBDw7Gifx0DgesZiPJ9h6Tjid0bP
oF7JhKMVgrFjZcTsx6yi63sWQaCfOUqq7zHuMFr5yY2ZP6LRg2qDmJYaX2fQGthSCvHTw2PHu3/I
3i/O96Irt8OOvHb9ADbxTSAfx7FkG2biAcSDwKm/1cc2hhagaJShocNpcYk3mAbttYYljZzKFO/3
tcmNmPfKMFjv2PNMKq4V6oBl+D4jm/Ts50fEZH1mGQDGdEBJ9U3nGqYNJ3pfFHKxELgvyc8PpINZ
vQ6M90ybtMpsrj5RRdhDLWlrd6xyt0AkMmxk+u7Uhh4/ISdejZAnQgpOzB7CznHj9vGTstXttIm1
PqPpVMF/ZuvPNYSSGgSplz/leL0fp9yuvbfY1oPCHBhM+UPuhy6GxkaRlzk0ef6TvVHysLqnPEI3
8EG8f2V74W/hfsicb2kMaMl8IY69srmTciwhztqGKU0Y9rvzPuqlCBdkmNI8rINRMNSHXxNu3s28
RPQTZWRB9QOKHa3i5eO7X7kldpLaDqwQn97F1s6jyqIrqfD+3H25s1apH4VMoWzCvnuw6r3LKHVf
vK87TpyVXuKhuc3qDzAxyceDjlWctWuQo5zupbIUkFXSlqBZ445Gjdzlp1dVG30k9oaL0kUAY2oD
E3r3YOTn7RWqfnvdMU3gu8xZni/0Uek+WdND9bd+H5CCc/L+tVkvpueW1EoEzhbWz2lI9BhvM5ip
jFa/7gag6y1Oy2lmABHjsOYrc7fHqaL8+I71+U+siwz6VBdIGmOueGgPnlR4Q69PCU98yXYiIRI+
VY/xzJQrADd9R0FTSq9KjfvYzDdhx5nFjvYuCxxDKTsjwILrszC9oQRz6XYqoaw3E1FEpKJ5q4Ku
NZxZdrQFJ+wPEIHRTGk/MKkSbm2+wfYw8PExH5hMcCj+fImcZFSt7tqq5mrGPUL0bjduIjS2qY5N
e6iQNdyATigeIKkWqFRS8ypMByNsPiro7MOvHrReS9JttQek+4i/uyVPJKpjAQVMh1en8ayV5nHn
6NoFexYiYnzWcPKa8bavFrkpo84RMdgp4bnC+MmLdJLOzS1unJvI+KyiOtvnr+PXjmXLj6AlgZhB
LjXSlisr60dSDxsFdYgMDxkmEMavkeQw1IA+lKWH/MfyLG14C/SDrLw8CaDKXjgNz7GhJN4b16YA
4FqV+3StwCAhGHanjYFVnfKnX/1T3ZT0PnnSTgphsXI/i+ItOxQxDMy7F8q6pExEWWYRTj8i7CPx
4hNMP+jjWgOBdY+Ox8JHCc5zW/i0d15vfWxBCFhxtxYu1TWvVWypmXeyXg2jv4jDVJ1f6OljexcC
asPvYLt3WBbQ1AVbu1bkCPH3H8jWg5aNQxjmujMS+LJIjIKY/bjgvRUFGq0y/EfYdkXLqHTrk+rx
kDlaAS9r1h86IxFqgS/NHK+OZusCgS40kerK0uiysOOFgACxccckBuhikXQo5qibUztGVuXtz7Q2
huD2ZFLtTAqydx0awdk7cxTEUT1pwiF+mXRz0pAUcDVKLLJeNzgIFxlgFvr0CxdwbBAwGITcErl1
397fTRadAtywR5ns1wQ7WZqHTcpY/iy2uoY50At9EOhK/i3SrOUfelkpqCPW3Gae6jtnii4BCJXc
ny/lXEhj1WLhGc0SwOsjhVBdLPD5crs1+cjAuPZYcVCDFWOwNhAg69hcW6AbQzVwGImfHDSEEG2W
sVIpPxlFLdU8JQRqhJkd/Jz/m9DhcmHJM3Vass5PFjCuhhQ3exoQbqWqw4lugvaRqzP/RaA1X1QN
Tjsa7BCcQVUtK9mKgsr6nRZc406TPnBHzdDUJ3P/rlXlMfV2UpZeNmKTS4LbMoV9XlahQ3A7SmnK
jOb9X2idBr5Vd6I3K3uuRr5yLYSWZrx//xUy7YUBtIgUVU/JrQjg+Fta1isUaY3rP3HZy1PBgmRW
fmuPixnJMimzhK//OgAgqrWRxUSloSrOT82s04Khwhbf/q2sE6RUfzcI3k48xeDQVED1EU7BYVq0
jMMskF18U13nSRqI+2D815XET0mOCoLIZDT+g7PZPT/KZ0QTeSRT9e2GVnBhtgHCBIrQ1xxuwb+7
tiZPWWRy2j33jpjZ+WKdklmXinh+3xDd4O+GutNI41uBBb6oyRYx64pNeYnFV1UbXKKytgcAhmex
Jbg1lAYm/gL86sxcYMCjTu38Bb4NSbLSS0NlM+yXnmln5lD3m69cXFG5EHszWvLaLg8b/09JhkpC
+0GJxN0KuMbcDQ+SAvJLN8ZLyHqmJsIxNzclWHQ8ER/VFNrFJ0hlgi5758g3JzX2g9MY5uzaWNUV
0rvo9OC46p1E9OwzGTc4FaVMaIij9TPn6d/ebbtodNohANUP84LA7K75EWH7Kk/RwARDlT9mPTch
cA+k0xSsLbjBXlWov7GBw+cPa7t99BsborJi873EZ8TZAVd+8i4/idJKDVX01H7kp0lEDqIQko5f
m9siBSEeh4ZV+/PeSs1+8rZ+iGcQ/aynHTpdVnjP2glmU5PfyJJlPkLJvjQEjP//gXVQ4uOJF0Vt
0lm7o8NnC4lmZg5zAxNhEnzEY4oeSL/Zp/wvpzAnwokgqzW8h3eEI51tDeK5o1t+XanJcomQCJAr
VUfYaaR53zJiUc57F6O5F0ziq3Mhm4gxFc1952vUGzyNDwDqApL5S4IPwgOUUyise3cW6wru+i9k
Xxtr0JxWIvXar16DorWRtvCSl09oTcICTQGsGTYkzPg4cjYL5l2z65tRrcbTfbNqGX9/epuz08C5
0Vv6FMvtYXZhfLZ8lbJdJVcOg8zDPiPh3HEQ4TnvpCxNd+tmBK6H/2pCAF66tETlXwsJOn/u1nk4
XdiJtzlMfLEjjpWL9fn7H8R2QkAFVQ4RyDH/jW4sf8wCY9IGLDn3XlvKtJsJwCJpKoWYROeZbAm3
dcEYqe7GhQQjuIvN7CLSSvFjjp5Lu3dOTCIFm6N2LVrgzANcGQ58bEzrOIlh1xOaiuEJYQ5Q542u
eCe+JPz4HE7siaJB3/YFEh8NXhISjW6ww5yWx32ZWyr4cMGig/7HC5gxKRoyySQ1nHDBTu3bsXG2
nXpAcaWny+AxxxoO4FywbIXaOwJtt7vvuH3jTx6mbezK0lEMJSI2TypKX2grLmYR0qQ9tSOWZ11/
nyLgqfmVrOPcBJsaEfdm5VYc7P+ptysgqxSM7fFRGNGfQILf65n5f+sfOvENcFdFd81+LV4ePAkr
AMDWBgxyBoCVZKoavfWo8xv6nakBY2lxQ2GLac548lh/uiUhfz1I6O559csOyyDYj2KodRG9R+tC
7RfbYq3uDRNpYaSUXrPpZYCtd7Duqw7hHyAIDKbsHCJvG6edt+sMierpNJlOQ+Rp0rrMsIywoXVa
2ALq9walpNuCW9DkATJfI3LLPc0MVj2IiLcpQfE60cpZC0ffV3VPA3D19Tr5OKdZw/FGhSfnA2gq
1yw5YsE1vdRs02NRPqppieyfcu+Ew6Pb8EE0xXrUTTuz5RZjx5tMP94HF724hIvreNllhwJLm205
04GD2e3sjXY/TvYqsuYope8Q7ww59grnYgfBtX6eLKmtuAMphwSgaXIhzjz5wtnZS+GBcqrMTGlW
ThNknWdlkymnu78oVyoYDeKKxCl7V6s3NFSRTXx2D9/6rGWMYZficT8DL5oqtZl+QIMcLS44qjFB
RpkWVKs447IrxKFAW4R2VmGzRau9ElW7PoZG98oN4C0frMGFQcx3mYSXaCUWK20Ef73TNMtUH0TE
kV1BldQpT+tP5kcyQ2+y5PqomAeO68MvD/Po2uHdlAT0glgPtxBfZJmiNGHJfUn9TfUip/DHIuYU
FdcSeVgWaVD6vst6focotop5MCIAo1HIVWZSrZDG3bOApZsJr7lJXOi3AJLehohW1qNHSq7bSNmc
leMs/a9vTRrXjUw6QPg58STX+1wwO+9wcLHrsQkaaX+w/g0uGB91ypiX4s0GLzC9OxnB74PrDk51
sMRGqTrEWE94rahtzsbm6ZgArW6D13ZOo1zXeKLKKvJpJaGVHqjq4HDBE/lgrL8x9yVG3nRWM6Kd
IoEQIea2yxwjEM5HbDjgA4o7X0aeHCTvITYy9d9zKkvLKNghzh9ZMaMK9z7GDbfIqeZHbVr4nVPV
eDwTdfR1DMLmGCZzsWtz9YSHcT/IqX2XE+FLw3N1oCT1jEOSq/KlISf9i4o39WYtleKHIw4JMKhD
3yKBDqDT1rplR5wq8ckbieK6GjRfPc9ep5GMC5B7+6Xp45Ho1H2IP14qxKWbgdNLNMbpY/A1LE/8
vqy+UTRaRzIAZgGTkrzL8Vsfu6355BqpkVwtUFR/KhgAqpOuX3WQ2xYaVdkMmYtsXDDVpihAHywe
Cy4Jj9+07dIO4bvOcDMvPEN9VAdxng5I8rYVzsQKmYdT3QYtjLjrRtaUG8nNuZ/vPb49wukYLhcE
wfSGpxUGBPk3dx2BC2crLBgG8ttdKQ+3rdoWvZVZn6TDQ30I2dMc78QvmXJRa0slcs9XdNhQOTMl
D8T1RqpACQ7WFmHN7ZH5snHAnO7dwU8W9p3kpWogffP/iddUHE8YACAsBKuDY8QQZLp9QUQ727hY
7+Q0yhk4GGqIgT5m/SUyPqzh3ywbMfLAnSSQ6MKwK2+tOzLnkkEsw4xcFNU9XZ3WzMh+q/5Oj3Zf
kB9JSOmbDKYEzNYZf+vdEgEmaSzu+PZ/hAux8u6Uot91PKm7AVPBQDaYQK6x2BYqegUbWxAded0v
epvPIfiEi0G11uKVKDl6DoRAADgjWDA5aONaAzLb0HmayDqsjltSRUUsiRcWnxZv/qQzu2CaLqAw
41uajnEVZ40PWdyj3MZS/cexwJuBnKcko/5NLD4K2SftpS2OZ6TyJ92k9nmQG8T5iDqQB6KTNl9F
ve1xhwv4O/d5AxqDRjy/Lfs1aaKMemuERxI+0EHdLXWF2NUA7Bua+L87pPgajGjCkmE2+YviKCfo
NzOVe58yTXGPZjjCH3iDy/I/EB5bXNY1kwWqMpKiL9ltsbLyQnZ22MURu8QTojInzuD4ZihyFAwW
rou8KpB3zkTGUW8B0Gvxzd+tNhp9aWS5vvMNKrNMPA+qhNynrehGvnQtJaLNXsSI+w97QOA9ajsp
YrSQNKc5Cs0H5JVwdugwW6tIwT51ggAFJ64vMvs3jhqd0VkA8ythkqPnaTc9+s5BsyizxN7PGzfD
HCG4I520mSZHqYdx4qZTGkwOUciTLbjpDQ+0+MZw7U6qttJ/y2un4MPliox6UNbB6LM91umrBy+A
dz4dnkIwZ78H9qoa80c6noJXBJ4ozaDf6Iw492US9cOSXoVZCWKrkq3GpRH8zQmvHtpyvpxRHbmB
FUwVYoLTougLEsj9pCaSIbNYDFo5chGvh5UmXzy5QzYA/9phY5UYgIyZauNhnjf7fZv2v6eN0Cs2
3hX4DyEFHW7Lh93w1QfPqhFDhvaZnKcKHkejPhgBgYwhWmBOdue8v1qrxhSq2GUdBFLTI18VCZFs
exZHPCBHVzw3D65/XA8JQR2Sv8tEq+QvVt1OanDi00g5ha8UY5lDQIQcI0Iql1SRj9FLA9ml+ERh
LzjAWLlQz/UlSRkf1b5wuS7MMMg+Q5pQbXnKSfNZZsj5DYqkibSsdfLmzUjvpN/OTbR88q0OFQ6c
C2y8mwRMv+JS7Q5sVHJhDAAMyMdn6/FwvWQru6cqlT/3nXUgITzv0gLHLeJmChqA+2/Vr5DOIt/3
Jg8tR0YH3HyxL9BgLEjbOtk7/O4D7akAl1ntHw7PFGT8faLU57xKE2WSKIrT4XsZ+gn6yBycpc8G
YHrfv906Nz+LQr55UhNLes8tdXT30GwVJmdJ1+Xp3i6fzGbyYoYF1mONIt4JRTA4OIkWs1aIT4gU
ry+jAuslturEhEN6duqseP8Njtz9QQO7XSGm5LH4K3JXiRLFJcy+Ho785fE1zs/IsGLZ72rjJ3YN
IW+PV6lyk/o6XbA+WSl6+s6Ll9cGbV/8IQY9Vfijckwh+sNSEriDn1rfSLryvrvahPIfN7m6OLzY
WRz7ecnsEdejsPjz+H59blzImbnsEnkVHdBktzVJL+EilIG5wXXhEn5JRJaH9EpyQahWybLHSNX9
M2qAiRJh9kc6KFaEmfeTW0K1/zvHyx0vwLiClG3IGrZGmS9h4mbzxuSxS9s+aw8cAcHrSuQH36mH
g0Q3gACZO34NS5DI/matCLzNrKopNdKj/R2wiS3+W8fUR3UgDc5RbnU7TgVDVeElzq2S/wg2pW6r
Hvc2OO1c5iH2sPRc+AFf45+yVUQEioqGewDp9OLLtNCanGVQhx6r39WBCZ0ZLC8vystFf7Ssoymj
Ulxejxene32o0fPPtLc0AxGTsMf/He0aQrlAbXfCwHrRpbmqpRQmbW7O30VdFPr4P0GLhXx6PgMC
xkdlcgX3QUIquyMdqlI7lhAlMwL0kBiAj1Yh0a/KRRiVrewWlEObi4N2l7f/SjPOmrOu6ytQOkVt
OC9J8N2S/ydpEb0de5tLYTcbIk94KV5gQs9FVkajhIeTJT0mVmZJIADoSUobWwx11ToNWfv/aevk
39Dp0WMc6Xq++BeXoCzKnbSj7IfSoiZuYS/Xr78d0mYiJwNiP+Ju3AFQNEIzqGBsAK+89J6b+mz6
ATIkkt7KfhMmOPJEOrbOrIuh2hQXPxGZWvXxRrvs/kAxr55+0zYCSjUBAXq/zfgcvpI6ORoBSzuu
xMzUrAJveOddjmvLwvkpWv2Duq+Kk8gwoLaVXWuDRyvwOR8lq0mS+VN1hxuHd6u8nwokm/h8FAaW
gydnnZVcSwo0BiI8kP8RXe58cTsxWzd+v4WXK9Y00yV0MoylPJDf6+YlTN9yuzsigjBxB4s9jguA
6Mku/TtUqD13jwWzJbccNTTBwHfauu6Yczg3mIOkUP87dDaIVrZISyeO/X3irZdbAH+dcRA8xqBT
JOlf6nJHZ818RpfxVuwyLMd5TLZfsptgHUCAzdJWKoQpna3SA279geSBgR4u5knNm8aOrWyv3gR4
u6q+ryi55FnrMsVFV/Kvm07PIxfaqOn5j6YKmO3tz0tT5t5+NmTxSbhLGJ7Yuvh8z88baEQ1BUVG
vvQXSzak7v3eLbkdQulxllQqGN364okAQ4Ekeit7WSsuVaAIPEUGCvw2avS/n1Jjc/yegJzSc44g
Bt+RuZFfybRgoXcv3E3lZj8SfKipsC5D9fDkNBr0V6IbBtDeu4ReAPN6u2Kun0ZWXM8E1EWI/5ku
TI6mBvWr7bzmotEp756SSn8G0ApcGCH2QtAkX3xC5PZbvVC0Z7JVxKtTZSeX6FM+IL7oHaZ/ImGZ
oEew1RVrqPEf2qjzXNv4J+1wiOlMPr6ABowNqrqyFelb3O+R/xihjo+yLNZ9BEz+/oLltZEShdHr
IqUFOqpWAhC7JSX/+FjSo59DHMxZSMfgL5MjJqYlG6GP67U2MfPg1C/bwfZi/99tVZWVd6K44jaW
/u2oKVA0Z0LIwrhvDH88PONYf8r1eqEGJ23ggH5uV8PYnHj1rzTcvyldlBGVnpSmjPDJpbakzwCL
m5qXlNdJgq8+7508HiRegBqpntWUTFdp7v+RLXJp4v3BJZIuK+emmHJLU2f+ij387g/YQj+YGXFf
vVNkY+Ss5JbhADx5SOmxzkt+GLzLwaKSHUKfUAhT4Su6GI/LVmQkuIRYrClzyTqCRVNK71vK8a+m
s4CLqDcfm29ywhmaJSng5Xq4o+5Cw36UGtHaXOkDbKeHkA+oCP0QQbLh1pgFqe3h4RiL6ka2JwN/
HtF4tmIfpZDnP66cTLBoYcvHWpyFZs+aUIeDIjIVjubVABmPfEFi3H479nSIKIh575U/kkAT5QHV
8pEBH5QSh6gsrNonl53ZBfR3iDUClg0dgVIIo1KGHEU6KFUokt6N/N4DAPLTQ/qJ30PjQ49Tp+ST
QkNRBPMhLesegeMrj6P2nAS3IcBK1jEobYc+6XK1zG7Ofchm36rG726ouWYMK9onXMBkAc6GdmZJ
biQY8vHIpfHYao1FP2HFZ7JBSgNCEZAHlAYqv0tXpoQ+uEPeIak9+FZ9dAfK2AS+97lDYRUPnr6e
lU6iv3AWYO5e3HtjARs8S3IGFCjYQgTk8sRR8LkPolKdR22Yiqn1o40uYnMZec3ZHxztJRMg+Llz
ohytdlpSk5P/hGkd3UhiD02wW8AZkIOTTf+KfvVNtEqjOq1I18AX96yoeMCA0Yt+rWJ+ArBXYK4T
7jeS7lUKnQ0dyC8n9oLpKJ/Y3vm5PLIrmzKP13EwVKVSxq2NmrntdKsDJWxr64r7+5IKX3mdbDhH
S+QXQ/lIukicmzf29rt2SVZ9c68cg/h2gNrCE+006nDerRoMEeWjYTFX2m3kNP75pASotHXWqTZA
UQeksM6CSVHyG3msVLGbzumkW2deJKxljzCpD+5b8w2HCw63Vhn4wHoSe4lpBrH3EvrDBE74uSeQ
XV33KOYCwU3KVYwD3++8QnMau4cL+WR3c5l69MSpIVgm5B+ngvkeV3N+x7ZGy4r2L8CxROjuJVw1
WYJSkl8XXoWRQfwUffTxdqLSPRz1yr+uHVyX7+r+Detyzg7HaqZBPtn3VwaNN6sLhTiYBJhWEAfC
f6XkfOCXsNySPVBoeo9ejh1faD00iEreg6wWtLxt/g2T8xwRgG9Xcnc/KloqB/1BcdyUWb8ta6RR
6fk/mHmZqwSJlGkY/haHUXQYOHFmhupg3iWLo698JqS5bMaqzTOrIFsEC+p/a+Z4//hzwiAZ6Zvl
kFpskVwDhlLeXluXXR5pCipAEz5aeDkpGSVTZzBsX9LYbecy8Dk+9WpOPyA+UrtT4z5oD/suh9Mn
PuEcnbrveUlsPo4F951WMcIuwg45+bk67b2Der1VO3j38BpLqPrTttXpTjdDTr98B86/u40/4SVr
ImSdHlyrSjdDcyUDZuRuDPAfn+jBXARNYMHKDx/Hs0l5jBjs0hkArVX27iYQXEyOLefw/xTwZyJC
UQy0zPQsb/gRa5EVZONgcZd+jZnhnQZYm3yHme04Iwin1nGNV8T/4arhTNufy0ldnu19h4QMSqyQ
sMWz5/LmLMz/PjzNp2DqSSXuUVf+FPJIdfgsQiReNrEYnyl+4mES8VB9m8Hill+gjsoAX3Ory3sz
7O0C0s8aEX4zma1V5kX9gAYOgVoCf0GfkYjhJg9YMv4a7kBWpJE9hsuhDtvPQuQAimSgJdq+5AYR
5tzF1TgjGXLdGtInBEHCqx4yvpTtlneemBT4cBeFtdk6WwkTqYfQqmO7o4smm6x/iL8PRlCEULTN
d8q1lf0HtoX9o02tWKq0B7QBtO7yEK7BBlXiz3w8o45fj6iY5wlPBHOQhsmzupETJAejq2gXRMPp
C+RPww/M6BwZKDQuDDL6BC3ZRhRmZTJsbjg4NY6a7xC/saG9PRBzrT0+TIKvdJSQEQ0yAxbrBrOm
OHWeRMj1cDqdK51eLK0EQnCwaLLYnS/YUiCSrzazK9yWpQBYb8gQo8jn+expicypFb13Z8/B/Yeq
9EYjXezl+pg9EblyUBzhp4jcSlGLPeBDhg8INduq4LjgcRneh5xSmaTbkg6/iaPkzTAhXWHepOoN
Bl8fX6WfFnRBeB0UDe4386xvgYGduVEbmuw+/ycVOKHbzOIKGcfAvV51y4C0VySMJdMrmCEsJV6O
ZBpCau+N2D+sWkZmzDBbuAMHQQfvW/ZPwYzPMOgaVDslr25bjC1f0NxViIsx28ZxlVrvTBBfrH0i
gyVBtGLuyGnh7f9qaDvD+DdPDe+kDKWuy4PE7QMmvVwsKtgcNZg3GEjXfMRnfzAcbR8+OUWiSpD6
jQ2CG8PbSvqR6fOmsevRMooolQF10I5s9Uh9kdYlcPIEeBYNpyiVrRzW8kD4+ujCmwZLYNdhnLRn
OxgIaAgtXqPGuV6EkrJbvFatwZpdg4tzRatEkD+thrbMUDGQ38T964sQKtKkvmjXhA4eAlD0HFkp
jNl/AZWoJVGXtcBy548qxh6iWCqEkUx0ncXljKGV1iaMEEYfUG2r4ClTgFUpjn61FXjB1fLsXXu6
i57aJYic3EmOLJqPXFvQaLuCEp4Womael1RD1WZ/JaKZyQn67NYYysUPxClcAbc7SJ4KUUQndk6n
KPlaWR9C1BZyWNqZW2TE/732yMaAsHt9TvyXQZmB+FKmtlZSyqC7GRvmNgbhSbixjYBV3aiqNGSc
lmQgl0XnZWPitMBVgqTlJoDSqqLS+C+I+u+XG5TTx/sJdJKXhegkOGCoi6BdhNfqZtFYPZl2fEBp
QSvTvcQwTN6BUfFlR7V7Gi47cy8tpUMNOIceEK+Fhv4ur3fzUG470RfTcoiILxYwrW+w17DkaI8A
MPlyP7cHalc9RCBamuPlWWQyhJ9mCsHoFPMN7QYM/BH2Mpc4jZISRF6gVaoZzffEAO5HjYznkWnD
8CoHfHkHeDmIrMIssGQCNfrN92tRsK7B/d5crl/2JMucr9SKx8KFIMtfCQN7XC1ev8/tzh5Q+zip
5QmvzqSx7rq4G6oJ+ePXVbf5RtoLhlrxKekndEtuPB8K4HOhbsdNucApnFVGcein2o+5iuL/sEW/
eb6WhgZKrAyGUnO4IMMgd3JZ/XAOHhfqnFSYgxbAOd292YyegfhJxGA/6nlGVUdEUqoIh3W96bZa
6RECb5rmoPn0kV+uvRNX/uyPw+9x6jra81KTRISbOH5JfRNuzVmDfp08ohr9MaN1cT38joMZKAFA
NdqoQ2846ucXhZBY4DRsNHX8EldDZyW7ckPUsmebE4vXvWfLgyzjPx4M70axrNwCBEWvnWNA3W8M
TwHkzDVX5pboL0efsxtF/CfKaMEKvRlf+2LT1w2RNe89seovq48fxNrUxC1192NX3AzYu8EVazcX
LKknGx9urOwW32uYf92ffLki4S9VZHbueI91AfOO5dJZmGmtfgjE4ibO3nT1t9t5hr3UvtWOkXP3
n7Y/DuESiYZM9jejostocZThRF2WNlZN4PZX2je0QqhmhaAmTEad1nVhLS0idhmOqyTVoxDzrI/2
Cym/OI4WxJD47Qa7iISNQBltKG8WlwLfPW6PAtbdKyfljwVwSvcyfaqB7ffnS8jTud6bncU5f0Bm
h/TjVfIEQoHwaNsd9EMmwlySwQsZI01MwFRyNrD9Vbw+VL4Hha9YQ8+7vPELF20pJBD2G+rz576f
5K43XZkG6IVNuo1VA26CYiEqFXM+R5yHyF3em990zrpIxAxX42cYmSX/yNSD0jgYxOBu+ITCu0Tj
nw5H4U1M3yDLm6ZGCpZsZ3IEqYv6xNKSLaW38kTKeW6Gy38RHK+DbUtMZtMZfvmm/27k4W2eZnUi
99HHtw4yNbk6lvUl7L/qDvcwy0WxNOANOZZKxdguM6DkcftKbC5aq1tDCSV5y29brlgMVdxBgkXG
Z+6EobdDM9eWJkN2az2hxkci7Yn3W43A6pPblDo4hsiSZaqRthgtWx3aAwCvha13mojgDQUJhht5
ctak0QaSnaUd48Q5LrgmZ9Ct8y/c2rA++4rOIjvHYEkTJjQgX5SoDCkZTTDQ9lUDIFU6iBr5LHah
3Z9QNqQvm56Lf7RVqvVvqkMZ69yH39TICzIGjlXXdGehoV/s/doRuJpcbCnseIcdkYaDUk5GFUAR
FnN4t+zUDQmt0td4bqRIXWM7jsGeIoZEFacTNYJEAyAy2ouoGaSiFzhm2xemC3MhWh41Y6H1Vpcn
wU5ec0mOXNgipMtXatDCS0kiwsDuG7bkuHqoQHygcG5dpxM4BrFqlDIY1YKnR8i6N3F/FpzypNW0
mIbioQ7QZT+z26xPPHm3OX0N55kK9uyjRVIaeTP9/b2eJkmtYAABhw4vsTnSZdhgS47YTPXQEZz1
yQdX2CSmGvDN7AWlCGd0a36AfWtYlNTz7oEt9iokC3Pck1Pn/F3feoQwTjc1Qij7inwLILrri8y0
5GRmiRXDK7EKh5NQwDmbmBFPxgx3MqaD2ozrfMPe2mh7LrshAH8vArJmEZWOjXDjGknPvA3wW0om
Fbx7NW0OFuswYgAO53HTdQCOHZ1dzlz5FIqRsQNxgla17W855XaHPTsbpdM55SQfOcrXqJTabwkt
b66z9bKsTvA8T1h+2soDkbKEwesa1M1cCqch6qqHM2A8eHQ1FtRf3euXbTzpdegZzZBA0ECy22ir
9XU8soa995Liodw7/N7LsP/AkCDSIKkRXiW3ToABIG85UF+88RF14H5Fj02GN7yb/ZsbUqZRSSaf
bpXCGVs1pmAxqcOQa32zXq6ffPV759k1uuSo/yO7XuVji2Tj/seRqfwxZFPM2Vm42nmfsQ8CRHbZ
7Z95BB6n94/aFkxhrtyApTYvVQ5ZCCbOJGDV0hzjBm0LxzurOZGFEZ0eOsmkOB2yG1z/1sb8lOXp
knHnDkDFEXW3NQR/V2uan/bRqTbQm95+qohiXsTTtQL5fHuaSb6w98GqKMcKpK19H+5qzVS58JaP
dk7ZVR2I3oWM8+Cd3zYOy7wu996pxAYSE0box0syEQQvFEpcc2tWluAGp+IsI7WKN2LOUKhQIVrC
VIRjJ13Q3jXT6TPuv3FwfcLRVfqMBPBab9qJ2/VnjHkRyvTK5Sx293pn2mk8lZaCYoFDQfphpHrQ
F7z7QBu/4W5IDVPo+NabeeBc22VyZTTHtK/PPBfXs9tHoOGc05/1653mpFnndmol+W/lu98O9h+o
MVSypm6wJjH6DaysFXwlxga/P3iQ9PmK5r39HFK0l1NmEW80lVFOWXrPlj34uQTaiuKKdD3VZsd3
kHeCkZ+kYJw0iZdGP0nedYuxBrBzAwbeVC1+1NzYXuazlST2kHeiFEf2tzuQ0GgsC3Pu6jXvnpFP
RFuESya1/YBO9zUsA1UIzbhxwhPTfAdn+bJPoF22y05Z8r1N2b8QsL60JDPDsykIbn+0O+ffe3wv
1EkiS8Az5V0pH0X/EEZhHcjbzJ4SgmNqZ6KWiznSGwGAwzLpCRBQESkCAMTUSyayPL/8uJ9nKSNR
EEveWMYeGM/P6L3iVe+5M2pxpRL81QMEB93GkV7FjG9e1m+XeaWARaWcDwPFb2GjPmCNEJZZz+fz
cmJhB7gcV1jE2SDMXQCSIakTxSvE1C5miYoAKiL2ySbzYpebuEiN4P/1F3EuDWT0YP+MddjezaoS
4IJ6KOE1HqYHFebeTMVRfCIshNyxDv4txL8PoUHAJpjEJ+4z59chVAcYLxxbyj6DL34ELXUzA811
c9xqrh9MC9bcZh3FpFYX68oRTPacB13h1dcyAivjDXxu2raUUpueUsG5RPxK9revcoAaUmG5+W0V
xuGZuO/B1LOXBL2313G5Srm/5uqqyk0iy78xHHwJpB1fx/d62zQ+lIZztkAHay+CkEhv4G0cBLc2
jRvrDTY1b39hyS3aDH5DzeLa+6W5j51mcmXPYUzExyM+h2Jb5xUVkMRCOdGj6Ww/CuxjFvXeKpQb
Mtp/9zo8rfV+iNhjU/GtzAexutbWjuvOZ8MZnRuCJp9qAJkWnU4W4NqPCbwL00Jhes18fDKe3mDJ
ZUmxeWdtWQhIJ2K6XOhcBWP128dbaMc+sSVKAfei1gT2+WpFtZGwMV2wrqzArX4sIikXItXLAU5V
YktIKIy7EUo+rPvoT86Cn3Lble8clTbMeDkbh9kqiWTsldvwMwKCXu9Y+bd/1meuBkt5wZehtfu9
qci1TulOKiTsKn9anzuEyZXJDJgxxocUNjKKN+j1dGs7kt+RjwkplHF85304cYsXsuIpA9I9v1tW
TG1/dPvD8lXDrPFYEFPFdMvsQ10qIK3ki9ddhlpX62VNNJo84mpOLULx6tZKJBhOTO9NduE+iBvJ
wmfGtZ3+ea7TSfH4tvqXaD38sEPhwGLVOiVIqiD5HEjETW/DAHBn6rKPSnnnvGSex5OtGpnm878n
uOw0s6dhmz7ORUmxD+6BKPW8mONwCjfjX3nC+SQG95w7LjLXtdpqOyTQoCVSPKwCu7XNSWBVjFuQ
I39Jw7r3E6Lld9ejDCWlbYlD8SWl6OR3eBwzVu/IRfXcRkRDlw5IbmZ72VtcUti1so6771JfxX4q
2PYNQtA6/8wRMBs1aiGIZAbZcyiRpIxZ+CPlEBq0XMgxOwYM27KlTbZgDwvwcEpLuUppdQv2BBIK
osVhDp86q6QRUiLragUg0xmCzUcSMkLWEoRAJNa8nK/taGKASiuZlRIV1KxRf/ZgdHGvIWjiSDS6
gcFmdT4Dgpp9qbnygAOpABit4dZnHFROetcNl14EQ+kq9GbjbTm56Qa1u/K4sOxRE19PlZaPTAqA
42/BqZCVoB0EHHpZJZf8Yo9qoVDgDLs5s8ABOBsXxZJT+UMCi5X4mIEk+3VMIHgz3v4e+D+pgttm
DLRWZl8zhBzCbq9APsB2vSORRyZ+tiF0ts2r5MyVwb+oMvwXqQ09xrogXyy5b3LqW+0zZhFEyRyT
hdS5Ol2wVqt9VBHspvxdW91KpHvF7c9rKve6WCexyl/3Rcd5H+R84ix4U41iOYbpFufQo0+GDlAR
LxG4X9tw5NwUaADuoU+YuLx9RSxyE1Q5IqqnGCBJhz8UIdwc6r+fMhZsaCJGpuntrp7wLY94ogbC
j7g9R8gE3EetKalgX+QS+KhFuB+Na2ErU8sc4oM1XTbiLjSbI6xm3Zb1s5fk49va/vVcaXpckcCr
7A2a/HBbApbVuhUM9SDq99qTWREdyOlAAzJKXfa1NYrLY4b2vZ3fbB+qNF2HtNStNNv3nWlO/Bpb
2yCd1tz9csltmmkGge6wm4q3nQK/MMd0byGLdyKx+9RQQGejjx9HkVto4RRRC0DgwoOnsCtrG2NG
Vqp3x1zmf76bwjSmFoAwRPheryb4iEoIoXb29StynWtz37u08lNbxmZJRY3+tQ/0ezCrmQozKjup
Kle6AGDfMH4Wekls1WQPdoItAoL09eONZQRbFo5KEqRHoehsiyfu1z/lSLE2uDm0tgOr6mBrs+Ss
E2tx5opnKiS7Cc7HM2FW4+1wPCHgcd/8zp7Ox3cA3m/7XXd3sz1FaGvD1bkQL30oeoUML0S+NBS1
eojmFNZtW7PeVFqCqpouRG8dzVWDoq1KMi+1ltoBzeVGhgXDBPTruGO5iJr8fuYf59LuLo8yJRZl
4sxhqfUHQ5PSayiLmIBlrMG/xBdOqxaFQKwaejTl6pAR+p1ZzWLeFLNVsn4hr5mTl/E6W+HrmH3L
pbQ3dCoARAtrJfWBM9stkbgBE+XXXt3C3Jkv53aA9T25NcrWezu4kiWU4oDGJqcv1Wgcgm31MkfF
E0SxejeVhGKuTN0Wrtf+7Fx2sbA2xvyg8OLme02N6PffCkq1lCY1NBFSThBTI94/M9JdeboZeqHf
OsnVq0swu3MDzJW4RXYztAiMzuuRgr3T4KJFGw8K9KgVV1yLiEiEJoAkEisclG2ifzqyco7j9Fi/
9vseAb7GdaUexHvhTTAYqIhuoTrQi5LVhY4XtyTVOpy4GjZyde8WZIxcosPkRzs6FUKgSTcZgSIZ
MYS6NQSFrNy4daApSkHFiZR5WeRcJQOryzyvwUr75phlqzYCW9xSJsxLDApyLTktkhH4pIbYkfHa
sx47WixepymrTT6ybajdTNeo4jJ9rZ8Z/SJUWVRvG6rXc7wUwVio+1sENA/R0DLGFQTi0FkPT1FU
iqT9QyY1igHCBJ4tHdOukpB7n5d2ipLp9rWPC0MZC6Fy508p9tj200VdorcLyEt6KJ/1yOVWvj+V
jqI/L62BPhJ125A0Ox/ZhrNjIJfmNPmM13yYm0SmYVjMCdZ4p2qfloPe41/1hTRW63P6fH+A3l8l
AewvCZ6r+a1Re0Tn4dMtOaOLdiO5KH5UvwPCx+JRIb3g/VWbmz43++T88fxOaOSynxHQU7Nu02a2
vM1itDzuO+aOX/gJZkXhyeajKxn+EhbKtP19EeD1LMNV+iDVE2mlWX41TNorBLSYlw4uKu8Ne95E
bbWqoSNeiofR6VcRVxL8OllQ78rzTZRgWvWGbsJrzwzlDOlAG3EH+sjJvqcbXhE/1OJIoD1i5b/5
ySk6mu6dN1AS33RjoVrlu78ugOtoZhZdL6XNKoFKW6NaAI3NBjnyjGPHV8Eq8TKZ8IIMFZsRD/xL
6xtlhL7xbVZzoUO/xph+jrZL0P48BLpmtDijO87BEJ0w+TLS2QISeQYXrmYz88BNW3bWT4IsaN11
atejh026Ko76Xvf+FUcoiFNHdr0rs9JRZrNd4JUS32C0SDZll330fjkLMo6k6xdQvjnVxceKxscJ
3KZDz0lkjx43Fry6x5yx/lqdEzpzkiEQDmbJucfv/j1hpy+osit/YseN6syGU1a/OFXlluXAG6CK
T7+31UAeZu6biU8NLKdF8LaXn18O/m1M9Q7kKhN+KL3nubQNqFY3T1tmmI7C/CwdFu/jsKhL2KO3
m0zdiPn2oklbzLW4rcqelJN3IOXVY/j6eyuT2uDBzvCxTvh/zL4/5YG4zqZYnXLwAwMa0lVPshMR
+a0o4rmejFJOUn50TUfix7Ac3tsLonscJA+0H+dCvzTCr06HIlWRZTQjltplzr5tIAsj0zz4fEM9
9/ncggzh8uwXhkgyFhfiyx11EI6d0sutq6MjrXqGyLdw3mXBYAihEKcKwmMo5F14Ul4GF5C41gu0
wCFQDQIT8c1bAa/NFh9+K51XBwplnbuS3f/FLarlaD6wvWWumHU648PFZw4Pr1/dSnr6IsfAGtu5
ruiV6Lyx7NZX1A9waqaHdqlX1xEgXJQVV2WlNmxOx4yFyS5pORL1M5cDJl+3KPQtnbkI5INuMcXz
HIZGdYGTWDiJJk0wGfN/AGg5jp2bADCh8vw9zaVoC0CQzCO0TPQy3jULm7ljlFhRZkNh19vbDll5
0HzyTWfsKJDeNkOYai0P1FYJJwWW9ubdzM9tIrhms9BM7GkiplzIxVw9JlxhKTJ/LVElD91sP1Hj
p97nVvQPryvOLb6y77kGHWFyOmt1fkj5n8ND28TfExCAJUqCxoSGGFby28Wq1jCuWkwJM/woctP9
pgdSA8U4X3M8w+iTiEhbjyXakoGLwHt0QsOvDbMWOrbcm+sVNWpB4BL5E5YLxIa69sEnw2H7RHkc
0s9GnzoqBqHC6KVhasNcYcv3OSS6mnc4sTxH2q6taSDRqZtXUogCkWE7dGjCRKtuFUucHzfX4cqI
wDcWhksr1uFrGqgLgadbqnHd1y+MM0/vlXOkzrsXnw+wJx/Vt0F7Z1MrQxBN0undDhexpWK4lbYT
g+yhQkJcBzK5X2MzEuCwLQLqhYlipW4XgFwOE5PBILjfU0uNELFBL235PRFgMjI2hmFBQbXCKAKI
gvs+ow/h4FlixhUSNZw/PBud7wbopy9GvF0mGUxLPjMvjtcyB1zSskYSeLktqxN8JVeT6rw7DWef
4t0l+lxRAcy1PW+Y0El7T7OHg4WaS0x84ufQwjZ/5ReO81GN/4LnO38X7mBkghVLF3ChTr5UYaAj
NURd7XrRx4y1TAmrcPA5UWna5AirFOv58r7Z/8XSP0IRdMEt58C9Xs04YDJ6n48G1yRW4jEZWtSP
TSvGLlh21oOvl8TfXR3nTe7bqcz7EUXYrBrGMcuC8tqEeCNY84hf3xuhz2b402eXB0sO4LFp09MY
EpYNaqi1Pv8uLSbujUQxYsNWRhunqwAiqJA8v+RnamZfl+rObxRKJBcdKbGNFwM5JIevuNzd7oFn
hKzWnEy9AqTq/FJGwAQHLIOpcxyMZWUmJGIg52qGN8HOMbVOTZgz77KLyyLNx4gGwRs1wHMzzIiC
v6SEtvdeDxaby75kcC4uSSzumGuMCG67AzeI+PSaNikFdItEJsDiBoltReSmQgmCNyiUzrjtHnc7
BoxhTm1UPdT/GGBXvPeN1cSJxu0Zu2OgcqdefBsE+Vfls0udn9FSr6tM9/sv1CZEfahMtoDimV/D
gAiyagr2RHv3+8F9LZc1bfnJ+IRq8qi/L5X0OT8jukKluTa8oTRNwLbD0DNxtAtv6HVY/O3EpU3X
+c91UIumEFx1neBktFS3kMGnBC9U3GgmSXY1hfTYDtrL1YWs+cYNjYvrPK6fZGb0U3FPgPgxeQmG
1xGU53T10saOWLJ/jasL4bikaTbwgoyDHLINbLqgDuOHgBU9sr7rVTcQDT5buIJn5jTVNZDS+oLM
CYa9CJGaGotVsjttzVS2axPCW3ZvdXw2nNyXNqqBXGIe/8bDoJ3B44GVfaBzTjd4eSsUiRz+6B8k
omL84D8PWcLLMJCuQh7QL+syo/P5IrbJazuFkjUiAQt+3sjatQO717Wwo9ntq7UVRpt+Vi2ZepnN
kttrpaIsEXxa0s93B2U+siH5g0qqg8wPZZugi6K7oIiye/0iPrtQ8IqDSQY5rED/fB2jbiVyMC5u
0gsYkokO8ZEsc73TwAxeivLoi8nXcC6Zrh2nWk/kgP5DaVoU2bdTn3aVeQ3pf74QckvK6mRWGAx9
k2cq245194Y+NJptT4epQJUpgw+zZJ/klMak+Obj5oqvxOsJjtGau7ZAP3Mtw604EllY1++vX7iK
5WZhXiq6TXnpcDLjQ5yjYP8ygsv1XSlvewng1A9fygX/KgZ1rCuER5d5Wu9BjKKvb2krAV1zTf7j
p8TPbFY8SapJN73eRjsAa4o29lA+pYXhglGonQ8+siQM8PRafK+CjCoeEeEWrB+M8MxyViIQkJKp
U/QxMOQJhcCqMoPAajtoKl2fHfuqaqhKRsNYiyGIfCjKarQGVD3szrZ/XaDktIoIPWJJE5MEXT0F
coIfiJxnB3OfwFymp+cJhWeeotAWHJxe62nZZyXGX6kVb+Is3KqMnGK3C3lIEMH+Dxtu2M8UqA6e
qdt/NiCkqgsWIPUMruja6epiBjxMTy0uVzolvT7pDXSF1X/SYB23SLa83NjJbTu+4vlHHrZVD2WU
1vwvYcwbHctZkHAVdCe7INN6q/W6CMlPhrgQ2VvO58yBw0lfj5Y+1EkeTro3uqRlV5Y4E9bSS7c6
1yiITNnzswo1BgWdlHj3wHnTF9baNnD2xDTncifA7dkKZLp/lnA+8qpwbhzt+LtSFbZslNRxoKkX
Nb7s/4TbOj+AjIZKOaRNpkXcYjSGOQGimrScetrQUXXCuC4H9aEPQrVVIzMqR2AmX8nkFuZKKsZa
YnvPvMh8gyZOY5Ix0xhYdOzEzQ8n+O7+BE6s/TY/xz3aPOwl0YgIjusa1Ek/ls9rzaenupyO5Yrv
/qsc7OhXux2fC6QQm21X8XeHtveIsX9QOmNIljEDYSY2Jpr9lA07jHdHpN8FkuzpQbNPuytE+clv
LyZ10VUdK/A65JViXXN/XUjRI00zoLq7dt1anQa8rmRIZsr4yyUnuqPOw96A603XDxO1K9S1GUwD
Sn2DbjCmyYeEzFxOzWZTNiuZSLx7tVJ21fbFs8e2rLIrGKaUhDoGkMfdHYOEoZwOwAmH9gvqTNfk
IGQnQcgJ8dbZ/REi4HpwH9iUtK2SBEdZXhDe9D2pLCn/Z4Hdp5qsjF5TjaQ/dhGwUJhn0WQQ39Lj
lQCJ5PQTftBesCGm6dI1utmoDPBGfynwMYIL3lLlvhHv5q2gHTlELgU4/eGZoVOqDKk7/y4/Rh/n
rsdyxnB8Ah52lGyfk/Ex+dCJZNcS/B0Im7Je3+SXPDca196QdM0ayY8uVUcpY8kIQuSrnnYJuail
Mg7Zw43466jQgjHGUGM9fdyqErQyhon+MeWtqXUr5EKI3PmHOpevxdwr9xK6/5Jw3952w3pMl1aZ
WYLw+1SvU+MuwwJ2GowFbh7zk75EjYsi2SoyM6iv8dCZfe3KTxef+6ad4+y8bym8ghUCWjB+nS4G
P6zJ2nL/06A4tRRs+Kbefvx8h0c09Jw3JipBU5GbAESHkvLSdxIxBwhUbXb39gFJS2VkgNjB0WZD
5nzHjf4k9mzf0Ke5fR5G86kGhG8o5Z3HxgO6znylXq3vJiBzAugWv87Hf3fgck+x03cQEahor/sG
Cyjf+L7zbnG0A+nadPyEqi+bKMe9NkcL1KmYOT2o4vtN/i64Rdy5+M2CEIAwifK1zUjdjayC2pVq
3vYV3G3ngwKdNQELryHue5GZFzcB2aKNhQA2mW1l8mh/QXHZs8FM5qggCwdnExg5BH3OHPXBijg6
NNlHF8CXM+qZy8zHsjzcWyNSMSb7ZTd1PF/WBRBrYTt8WM0UrGNLAL65UgMPns9hU/AmgZWklc77
hkgog9LoXixUs091wMJyE4djTPGQxMO7ItynK3F6sKVqYHtW9bPzg7IXn0BLpIjexS8fc7afra/+
B2HaPeC6HzZVcn5BU4iAZPq+N/rYNipXVpqY0ZyIl1VrZld9tKv7drs6eZWToWa8p6CPm/CEtToT
ah+9mishT76Up/laTA/qz4vWI4eIfIkRmzcK105CViq8QgoHnL8Mf5sWFfxhWXpfuRAPeKb5XL+n
cjd/jSYLPhgQ8B8C6iYIn5ixGPP36lLIy9DuMD2ki8vBfPMduvLRR/y8S2dC1ynPPY6tGRbkv8Qz
g4gCTK+FIT/E7UGMtPR30edlpy8WrSJqdIY8/fVhAF1SP724YSFcjDlq8Oy5+Pi8oH9T5xM3fZPz
NZGMafnzaoMkIyB9PTZPwuHSqP+0ksoGa3KaXAvAspZrb3DhZ3wO6aFaxTkU8XCI3CI8Hn9PLU4y
WFE1B5a0hVOnhqWbthPn6MhPU5QZDoYGSD6VA6NpTRU6pWw8YyGs7ik38yhsq+eH5T4yLwkHh3kq
GY5fM14gcwnH5h71NvPwH9v9iDiRg5f+OCmboVy96+Eio1AoJMD75sNxd0JCLX3ND/nnIX7KFX0g
NoZI12OgoCudrW9fVgN3lNYak4lZLLy7wT/mnur6SrkfRVXXls4QWvymeMzfaebugYB9cndJvldA
xsIXtq1ANcldTy8rz1zchBoECt54nt43OB02bhKB2o2yEvu/laQFW0DxZCWBQI2B1XUHV11kngwp
lDo1EWyZTc/iFY6DeAs+ZcyT7CL4zwrFzgWabEKEDKs7n30BgF0+2rKP+Qo7LBetzmJmumF+9jSz
yPDPenE70Z/46qioQpplCrzJKK2yOSPTDfKPvTqpaiv2IWEj+8dUFjQx9fPi4hOlhvPEgg23qFcM
ti8BauzACDIFf5DrmBdZ2OUUbwaKocArJhO7Tuc3RKy63YCyY6MKgbEsKVoUsyM0c2JX1t5uD8mp
ECXNy7q4fI3ETm7CrSq3V/Qbmypwp0WH/hzLuTHregNwxI4fk38worg7eGeO3JY/ghKBohLInzer
c2TYxSJNGFFA2KRmThIvzwUanqpnFLcSnaIh8G4BWQJBI9MWZPqxdA1OLwmvwVjqiUNATZ6dIoCs
1/sooiZKfUlSHtGz7JF4JW2hqioAnJAs4YMEoHe+ck9O8OIolSOc0iSHmViJl2/N01gMTA6JEH9C
7qXw9wg0FJUqi5aZPZ5Vam2LMRFC0S28gc5Id3ujKXT2mh19ilH5u+eAZ+369wLCfIWV9sQKdsil
EgcscRs1sWK8cJxfSKcKRspgQitao0pG9ksR1MrfjqwBMKcfdERyrDC95NXkKiIRhGvE1kM4t81e
y11uNC8AgiYe/5qO4YS7Tml2/pFNhZ7g7Yk/AC2lgBzrN0hTLigyH8RzkY/rHaJyA4ua0I092971
9OsXC2TE/9BEmhX9kBcftfBtXgq981rl1mW8FYUjN2Z6EdSfko/V/DcebczuwuhdIGa4AHEOMsV6
SomTbm15FGQOvv0SFteRW31pCKFqUl3eGaKDUhaLFXPQBlmfOkH//pRwefcnyCuHxg17Vn3drIqO
2/vhbkSurlpwM4ZvRXA9xmHjFEp7AW0j+KmYMBaG4vVQ2UCH8nwZB49bLdi/gN7YBlQUsSJUWGt1
HXzgPB/j302TPIOzOBO+80hc7sXKe76pHOFwL40NHvLZD9gQ4kYAYZ5AxSpPvZcrJND+kSWPM6s8
9V1fbOQ4Gj0HX2GJdO6/eIGztiNZu6MxkY5Bn0STqrggVxr9SGgpx83i8H0MqZYtPN36C618/KTb
wCvjdBZfRlEBC4WLs4o/2qRF+5UoWLDcCHYvhhv0HesDVyIIKVKH2xCyRK6qcfL9nRMCyNUqb2oB
Z2mxYgZsqZUCOijJEARGHZWbwryDNEJaObQZ7ApAgkquwdq6zIgBh/5A0kvAsiLsoWHgbGEpWHul
3OvuxorJKBZ+0rrg/2qGXUFGV11DRx6xGUkMnHj6lHZhMZ4nyR9pDZeL4w+mfGomH3Ly8NVfQMry
wEZs21JgGq5jvdKAaD//j4WDtJflDlnK0hath5mfZpLgYr5NtVrY1H22mGXleKT5dBGnZisQ96FE
E3nQR9Enlo4o7uKJd0GnRFnVWpinev17M7ZTlcNdqIZznIleGJoCWfUNlBQQrssZMSlYHjrtrmAI
7uHe3fzYtenIQFlIUcl98j2eMW3uMF+G0iWMSwT7Qgp12pHmQaqcWXfbaG4CGoxO0Djkt33aF2N6
vqfrM7PTLAhQwUvFPsOXa4U+JTz7egtskgIrQMUPciZIarfmTNpgSGTe5/4DZfzrd9eWcK45kjRe
c0QkjdIdJM8nG3V6h0KTfbPvVSdiwBEJ3mpIMp1l/yHB9PR5VhKfwHRMVyKsi2ycly87dyoXRsEI
C1no3dz9lrU9TRdsQPm8dHHJhXyqhXcxiiIqGX+sAvmBhOLwtsxq/jQJaJE4h0pZlHrc5YtGkwB5
mLnwLvJMTlvtmqLSXyXkt69eh7FamNMzOc4fGiPE07GH5lIPvW0OpsWzi2B33pekY0GEkiTQDnOR
cLNFEvD+p4NJct1DLx9tajGqbIgwKGV8p1THENlDXGJbuGg8hPn91SDgx043xbapevK5Y+cYHIC5
wJYp4VTp1dBQVBm/6vbhUYbjg+msxEM5f41lwm4yqb79NuiAQ1QEJEVacJDM88MldFZ3Mzaat/9/
927Rz1cQR4CVxTcC3Dy9K5Xd3aPjmTD1vIoERSaUXPji9KkoIAy8tVlbFYSTXrQIEmXnm6YR6tPp
Ye40j+7x3ENo7eXz3SEaZv4SjN5bTKnnULQtS+arDUxB2JQ21OxcyjekpvD2xZO0EQaJ+Ls/VF8k
GKZIkq4OPmWi66yjYTJfii9Zj747Pk1f5Yc7t5G+T6hTrpFl5jkNeNJB4gY7JMa5CZ1Li9Hq6cVY
/xlLXKEV3sA2nS4tbRwg6eGSOn7cF0SsRvu8yVfTQ+woOE/meEMh0CBkw7BGgUju5XAdmPEYxJEF
vWX5EAXdejo1dKckg1ctLb2rKrJovEcGx9/UynWKWmRXrcequkphiHlb27/yBDjiWiQk5ZT/2cc2
tNVLnEUOdcTWXb+cadJvaU0QKEPJDqW1j0LGVrfK0zCH3NO7DW5PosbaBetCnGyC2lcgG634pt/Z
SnQr12SKSERcxJLI7fEpPkXi/ttk2Ph1cFVicp/WMc7AuLUlHJ4wV7+QhD5B1PajeuYB0jqwf00R
PshAvY4ZIqk+jjxw14/67yBdhWZIaXE3DvU6qyNEHVx7ovl6YPHA28RMZfz9Tjmp5chEtzSCgDP6
Sp9Huy70pnOgNWC8BzFeXiMRVr3DEX7rSvVi/ajPxVxb08OLY4SK/WUo8E/LktUEEtpHq0T992g0
ZNFmvHViVccbm0Se//OnIJdC3m83S5xFOTmQ1cOGtAk/5oGH7/8HQFhHnRh1u7D1/R8yiOvjxGkI
WyLJi32K0UrD45Vsx7AbJriIVkjXTwJkDzUmRAt6WCCv9u1hMVromA7eh5Z2Y2MKzD7uYfHbEfMC
FXiwkrneG+EEcW4rk9Y/E17yXiCbRDJogpO4B23O9yXkPXuFOIcTV6zAN0r7IYzYVC8nzJSNfCqz
b+RwixxhyFbMxsls8BrGgUwEq+c51InO8abuplnpZBgDJDqluIh2G/4Mg1AWp1g4jZKHy8Sr0bZV
IzMaOWrWQWb0Y8NYXx3XcagbURvPk686HdOvwsOVFQJSOUskvJbYAIWdq+Kj0ep4avM7RmSwX/ig
GY9zOmfBq85UcwUwwYmFX2QKsVqlN5ZeaNWnieOU7jGTdKjKTWL3cjDr3pckcd+AaPtjZIuDrtWS
92nP6gCF4a6M0JzTP1JNIl732uBqHV43eyzWxkZiJjkuyLj9bP9GGc7TJ7/tZRp3k2v80E6RnaDF
ED0E5+ERTcJoMqkUp2Ojlmm4n1cGGG2OB4at+OFXf3SsuBtZPVEXN3QxqkjPbdqK3stY+jXcjUfa
h8Bvoz4f+rc/6DojDn6lPaPqyrvlN7i+V27pC2orQ8dxNNZ/HiKCPPmQZVdWK4jPyngOpLWjkjIG
daeBMhQa4dNhzGTgj5whG59xamo2H5nUgMGDkJVf6FDoOLpYGPyqeqitePeMc00pzFEQKcM7djfP
bDl3VA2srWJFd+W+o7SrXD2J/NkwGLkuw9uYnNUQTpq0mfWjHgi8+fHisFRfNBFC6+m95P4vEBy/
LdwMZwlwjN3pJXy6BRhdSVSi78FSSyDo+jzgbNRwaChtjG89Ck4gDk30r9q76dUe3QbsD/1gmOqW
5h7RApJ4b90hSYgcnzYucmKF07Z4C2KCuT0NAaHIqKguuIDySKvCIQXd5Cy2OQ/TdVv0n4ZyDLrI
ZLeUpfokLVeRjdyKpFHEFcMpdcETRy4HVvJLEfF64nBg+UfNN+gif2XxTYRO6/ir74uYCgWS68St
RPmLnnueB14E/inG0z5MNZ3FkV/hktFpZWl9SzQmKpZAeFRjU26HVB8yX3FeGcWhb9Jz5hz8lVVZ
TuZRLotDg8rQrz5i7ScXoie07fWnkOIvZOULrdQVM2iHv36BEih4MsHcGJQxUn1LqeKbILSaxaYD
FRb+R99Hd7dEZiw1r1NQ5GIFnoKYs3Leg1BUwab//uJ27fp0vj5ZAGrDA9WpdyY1Q5yuQph8V56G
G1Od5vYLpZtyCQHsa5J0ICF1FArWgrYRpHuNNqzZ30k1/OIr8nQUJp8edQAbYo/LHC4X3y7m6eKe
785dX1ome2ag5iovuwEarYpESwalH9ZuY+ld2pbsmfZanwKFtZJvuJ1dksepp00v0tweXiUk+c5g
fGX6oppQICg+nMtapxOXbQCLwh0pIgB6da1fO1vW7CVQ0aANt7KYs7i5dmDWHt2ytE/jwdH6tXlV
3VMVpAa6F0BmFyJpdWeF/ULKI7ltx8DSv1WdQdfM45M+u5BzKGv1A3lF1ryDL+6vqB3ArLVzz1aq
QQ25OrMRp769gQNSuoL93kJ0qg/JVR2Q34gCWBj9KAJYGi+ObHkh5u/+/ZFW+pc8m5n82ouQ9kVg
Czk1qzpGSYUZGJ6i+rhOAkkDbQo8MyP8+NQnbBjXbmLu1HYfGoFDa/ttqOG26RaXpR4Bf8g93Uo2
82TclWMzMtDjq2vnlJXSa8bturkQSSbHZVR72d0Uy3Oco4+R1F+Mu9kA+ITFI7BORfK3XdPZD/Yj
UM6ixL6KnFyN/TkN5Nb4TQ3fZB/za2P/8dddivjOntdvUzjkcNf5a1uipf1wmvIC8CIqEL2leG4A
m+UGBuCYrtywOVCp5hCANbpFt+/739zsZeaLIDJEmAFUXtpSUsgt0c/s2NKzVgywu56oXuYV4AN1
TP5A+UwWl60KdVxgqhiE85c4YDM1xvueMIjvw2838AmOwgacThM06+RbC1AXHL+PVjV4xwv3YsSl
MSdiQuaQWGQDzGV/usdI4UetPTYswYGWPlsc0fk9FJwMWhdHMWrMjjgJ5G/L9zUJ/Zhp8zD4tAS3
sXMyyz0nm8OW6ldIJViF11Ppvtb2Kde8Zy4JEq2hGZkUq6r5pAMZ9lN0UiJcsRW4Wb9Bgf3IJ7iB
OdKa4ttgUW251wOOyAIFhsXyduhYxVZRc6uVvbjGKkePKoau+s1dzq//cCuI7UIGV0ny9of6V7Xp
59+Z9f/ySqImxkLZgVtWr9DoNKiQL9E2XAIW/2BZzz9xIyriEwmDBczTj/pP/CbG1luZKCFZsIuz
1GI0lpogCMMi3kBO5E556Ab9QOc3I96FpRkY1L07CUDjFuWjKhkuT2mnbKsxOxO5yxIZSvZtsQ0y
AvHlkuHyTH/GA71fqyxXpaHHIrBtwiJ9se+2SNZi3g/R4aTwRuM9Jb+LRbUGou2ODQB9gsBlEdmj
rU/QBsQdS7FQ9vIM4w2nifyIbRw9nnSSDN7mo1JGhfqFuy87Gr+IjR1bDR7VIU9JV9p1WxxY5XaN
v0KD8mjtUrnsgs5oh1FZMn/H031gLxyCs1aRgSCp7TO0CopfRYvXnzb6E8noleAxgkfKa7ndesIv
sFy4wOo7cTiY2b4C+N6VDWOiq1mYDjcoX/fw5QU5BkOapXxAwn5Upz7Zi4t/zK7RsnpQaKwkBHoH
XZvb97Vj6nZ0fZliGZqjq0rnnPibm++DGIX9BLyXvenUiAG1ZStvfdWyoPrUp2eSh2RkVsSI+V7H
/qLXr9cqtS1ImVGk9SRb20Tr+9WfecJwNFTtisYdgaYtz00u8LXigeXT0J2RZ/Li5FpNbV46Onvw
EfarBeJEMRrnQ9DnlzwFwUsGR/gUClwGf63mjKEEjrAf9RQulK/nDNe2d9kfumfiguDrCMVyVeuf
xwQb+IY5s2igYhvSCMwcIIwxXmeqd1NkCEV/He2T5xA+lpQbK5BDlWOGB7mrLPXYb9o/fFlxSC3K
EFddmGkgigLRqvL7sHDqVCo/wNtmYYhJNDgP+nIUpgS7ljdUxeN8Ri0azrwMxtMvjAHh3hav1tzo
DlENuyT9UrOF3heEw+gZ2UT59VFTKSmot7OlA5h9FfZOsdn4vdyZL5XZ/p3MIGvBS1Ne2E0kcPCD
AJoQYahthrAfZKuKIFb0ngK/reMttxQ9vbNfsjuOMlJhP00XLgc8Q9vEH9JgDQvA611qvaUeOfV/
IxElz2sjoQfEeeRlQB1LkUL9URUU4Lzbfx+bmkeL0ZCx7GjBOgAmKOM6agJKda/Yh6qzd7ZQGwGx
mov8Z9UBvEG9AgcHCE0yLynaC1/xHXWecSBOOhWJ/KLTzmioPBqtnw7cp8pJA0WGUO9+dI+A/zYc
tfvJoasCG9b/lrLDgsv0a8+sZJIvC6sKCDsgCMGiQAP4ObtSjfOwUeGQy5M0Nkm1mvRPGvhCZofC
4057PlwXtNKjJZvxaRMGX+DrEi6t2W/Dl0ev8Pmrn1Bellz/hzN+0TswO46jqMGCMFjodnyrOKgt
YdY2bhLezEcRDM+z8hyMneeDxeiTM2zWV2FnrHB31V5VZp1d2WVXTZf43fk2OyEoXHOSqszz1XbQ
S29Q9b0wMJFvNPm96SMNrHNrInYOFPheui/xZVTJ7qTFQ9Zmkpr+dEnHgc0C+ysxwPRCADTv8IBH
Lf0MDNNCx6rMIIdU0z2e9eiF/1xqTxSd1pR0adUoAnrjNKc6EFK4vvSSTd9p473J5sS+ENBZTqHy
P59HHRm3fmXJqP8wvhjHDyCWXw8W04ekVAUldaZf9jlYf5fnvc6s7qpscpqFyngu+Eq72YXRYuNY
mhtxrMKd2DGMPFxJK6QkaXCYaTC7RAsFE/lBKtoMDz8KcnKZJd0Z/qFu6HEKzRr6vo1UG184J8m8
osKX6Bxv9hJUxOi6zqssy5utO6LazYBfv1nhZm2mUmNE8Bxfczoll2vgyR5qBAaU/nLmhuO363/T
OqqlBx24O5tvYVAgWf68pMCFCgb42HUrYQaZ4aUR7/loqdk50K1qhysyB5nm96/jaXDXNbXu5Aue
4Lkphe7en0LLDqM5ZvYIXHrGwHN37vvJ7DI0I9x3Ki8KLrieIWchm0MAVb7dc3he7FcA1/tDkwMA
/5IyQ2r56mSJ4IGapK9VE0RPGFMrtvLNEucwgSpHFa3I3zNANGX6iaAAZcEWM76HY+EmC2Uwd0Z3
E/K/MvzEOQFGjDsHtNbiDmFTRunw/ikTerQkD+fWX3MOYzsMkDr7vHhaiPFKe79CT6UntZxzUt6a
C6YlDNWszuZIMgPGJLsc5k8dPANubTKH5M1SPA+YoeZbveWZEmV3AEPVsa6bIV7otHzt21PC3QnB
a9uLWxs6o4IwZEktBiwed29bpMNMxW8uoUrCGBiysgAmrUSnSbc+KgG6Jsaf105SBnQWPZvCds1g
mUbROMDUlAoM1Gi8ESK4EvagPaN8rhfq31u4D50/AelnUU4mv02tet0LDdm1jU4FTq78eTjm2Jwj
B+J2UifsC3I1lPiZpQWylkUeC37XrBC/ObMNsU86ryLK9aE8dOqZOl+zQdm62iHyoxa5FMXlO1fz
pmVztbCPgVm+ElF6yhpqj/1O9NOXvs67q6L1rYLQJ7+OIxPjzxExFK2h7Fb7S+bFQf16GnBIUD4q
aP7ijNySd7L+r2OZGIM06t3+9hWpoht85fky+wESG7ZIK9y9oF+9CO4Ni8cJ1CjTeEg/RNR2KYTb
ahnKHbw89AJ2ZCe5EO+7GmiosPc466eH6uWqTTMM+Ss7YqNDo2B1/RDhN2BLoWCqJL/0mDVJQ6JR
RE3+wWUbKgEd20YfdFmECdG//EIjsJiMWr/IO2XTjJMG7TfcYmnu6hxFwU0a9DO8n4YVn6Zk9mPK
OmYeFi6vfLL/FsX0lBQU3rbvGC+4109HVQkuVZjIsUiR/XItffYo3es8qm54KYs1EQQL9bbBewI1
moNIxJi4mAJel/vWs0cSLY4qDmIEyoNZQ5Ka63HyrG1Xdncjc/4VIT4m1qvTYRvVhDjaVnNbvrx3
yuktzXqaz2SPxPsyV5UykBIsv9J9u/TNnOVOw9l5MeFZSqvUj+O73ldt9Erds2tKnqFp1DAs7+Sk
tgjs9WvFwC3B3sqa07o//AQTkQFhWiRR7NT4+4UuFUYOGNzlKZRUZXEPu+5imTHaZgerXbBuVOVO
V58OsCBbtiUn51JqKaUBtaVP70suCeg/Gspe+ley8tnLFlTx04rl2iGfsNDUKqC12ectXsmxGHTU
wnbiU/aJncsfpXoqTfjFRlhOFvml9vHivM/vXVvaKpMm0xu6OERLXRNNS1l4alw8pLaR0cjY9z0Q
L7P4hoPPBNXB2oC0Rb0bqPPpf3gC/3dyUrGtzEjrlemUDEsQZHK1bYkMwwl7+SAlJ0a1NGK6LlY1
m057PE3LvpWWYMESUV+ocJl03EElOptPLIWlkEGlm8lQcBfa9v9PVbPQWwu2GZWU8KKOtyzIm3+K
Wn4aAMrvp0DfSvWWeZCzgE2Jm/krXyWqcHgFXiR7WjeHBPQ/+D0cpB2P8TpbGa+GufH2OadkDeOc
Pzg/tZIGa1WvLbk9JjohBT1b3eDlzNcqSjGYRrzQkYd8bqr7g8BhKeDef9fUN0Hd+sF+I3rIbpdM
mKWOKqADDfzkVO7pkXoemDElE0RtnFakRkzbPwSjb5VLMp1UVJlW+gKhdVTAL7AGhtZlOow6WBIn
BSaN/xdeglwirGRAsGO7i0yrL1IZKMxWjonhIBSgJCqLEewcmUKv1I78yNpG9sE5ELFez/+W4AWQ
rwbGA2S4kDZp39Lzoqh3a2kbkl+slyjZ+vo+Qdvwsm534zR4zr44rRWltFVY7R0jHOyY4QL1SqWo
72Dn51JWGobJxhvcwl1cdpi1VsnlW2WmjBuv6y7frjBk1D6tiroy7GSAWxV7rf36Z8gAGCOV6ZDw
oX6c/wtsTsEp56qvwaKSzhMYrhF0paP5vOAGoJKHCx3vvLX4RHq1WZiQkgxB6CqZsmABKaiykZey
XarrbPNAG1gU/TJddFSFFpRDo4VA9OtM3h60PQVOjzFz5xxyORLffpceizBfV61ZTWnPIlcief6O
0jVPSRz+pMqbz043bfeEMRej5kA1/OB/GALVQ+MeGC0f5vRRh/ykH7QdDQ9JPUcebJqg8RCPVGYR
I3aZbBc27glxpcoCxuuXuEKK+tiVCFFs1tTZUA5cIwlUGWNLp62LzrwB4rbGXFT0n/Qg/kdoTTSG
k68MSeCDfZ6QBX6jR8V2TOZCDdr3wD/awFNkW3UMND8dLU6TVdy0y9kzx/QKxT47+TqINb9kDKCT
PCIyTdHGOP6Okrr3OiFcwBgJG4bu1bSPpTYc+ws6xMwPupQEEsmCf/2ROF0FC66zYKA3eVBgU8/H
fFHHoVOdTPfLYmIArzly3pF4+ympxMRtxmp621Dp30tEa9V/lx94eQd5U7IYkCj8zsfyC5fY8olk
6Wn5y9F+7Il8Mb9BCoPqD6fKPGvu7A6DyFsA7MLvM9dr91WEPeNC7Ft+OJBBH7Rzw1AWdYvrb306
ZVLpwCbvTxv+cswOjCdjPJIP2R6JGRycyDZyP0BNZMEeVfu9YsFr3kLpvRizjhXQefBDVddv4Acj
b12JRV2RXgN6TnUXCIW13fkj7u53Ag925Hmhj+op+NgmzwrGgQoSxgieIPQcuk4CxlZWxK7Xalgw
TZ1aq8LjJUUYiSaXsmnhWYpSxryPehHTVxzPjoI3p2keO28i6HZ6bFhjn9GoHmkG+CLGrjBDG0Vm
n2QZLNJIwyDy2LClSEX0HWvtcmIUTuiiQ/Pu7auRSwL0U0ECqzc3L82ODf0t93zXQDlr0goPc7Ar
M2rRFSwHSuh6Zj3mUCOHuvgAjC3fbwRoSdTTJYc2tPEsJmdi9gVigGw+xAOi6gPL5dW8KEYLKq25
naO1xAGvW3A9O8dR1cYF2EDgax8qIC+/xkVN76mysRbkph2H9k2aC+Xf63GLCCiyF6ey6EuBH8hX
UZPs1Kvt4unC8MSz8mt9P6KKd333fuhLoKfULW/EixaMosdo/whRyn+B7zIt+k1BVmfVNhrh5XQE
pBLW5rEEg+wUkCHAY2hdCEbQ1iLI8hxhmRmtmsRjSHgKErWnoUMIu9zz39r2vZwgwjPYZb6zfm6l
nTJG0aJtuDbn4VI2/EUusd5ftocStTqvw5O7pstpBHxxsYNO1X8YaTETFCwyGr9lgtRQfAfn9ZYl
5BNGjDRjOMFQL42oAmL8Hj11K2/9wCvabwAzReoZ1mDcpV0qSESIZ7xCVpNJypClL0xsi8Hbjd7C
8efCLqg1kcDTQxsh038w7J4SkyXvsKHnq3O1glpiSGYcLYIlHOa3pdmlFSz4gfYTFWTAPRN+RW+M
xMTX0gLb/PtyAuCodz4F/K1C0dZjiZY0effuKZgAvDcmSfxPDOsVbZI7VT9ZIzoQGcXLY+Hjy+nw
/uj/caEttX0QqXCgeRtNdQjo1FcQLFS79I5HB1t1wm6Yp9lF5uKz2bgVD24edqoIIzIYkH5B7TZ/
nykMCcI54sJN1+dkoruRuuoN9L2oBHPIdD0cnvv1MXrHCPeMZvPR+FMpvNdEvO8NwQ7B2im+xcA5
yNcfPAOEO7sOFVrHalg0L/crKYfRCFyhHIXKNPCAxsJbhqN3AnOd4SjsA80HYp8taFgCkNIidq4O
HGcYhaG/xfFSKmybHA3OTyDLKdcg/rTDGMHA+WuJshtpHgmlXP/WO8dx77p6wsfHTgUbPp1Q6egQ
Ne5Imp1oDyIlJGhEUT8V+rAzTO1ftxeOLRZMTi1XWImkVmPQ4TBfkDvaeAn0YMoUxh3i390/WBMP
4DQEpXe4Wbd4u5HQWkpac8lQvCynnVm7DQl0PpMl/5SqDkqbFxhJm8ttIhInVJM8OCCR0FeS4UjA
Vnj3k3Etv9GSQrF+iel+8pMvKhJyOXVvTx7mau+CU6RDWLSGf51bp8q+QQsPp0VxfleQ9fJ5LdEf
fqT3We7t/ysQEeQqxKtKxeXcrf8HEXmey58P4D/l7DRA1gOIP5/QauXa+DvY/lZ++8aX7RnUPxbC
9St9HxW3Q8FmHg2kyQR25isfUE197D2vns+HFZngn7v7TmdphMenfiLd2vvIZphmegZGsqqE10fd
dOM1mVCFfoixXUdmSWQNKoLf0bDo9i/oXB/bkwHew0eZas9iwnNRh7S2dnRNQk2l3eAKxzBKz5np
baVgngZzed7xOnhH0Yp6pknOBEklvHRuCnJtc5Lvc4XECHWMxSvGLVrUGFKwkxE2NiHiwShTmGv7
pBHe39EyTND9xALALeiZ7JbJ0zYXVzsSw7ExVeT7sI0u9OC3rDoxhqjUPn/NA9Vr5675ZyD+o8Ot
wXjaLxNtzHPjf+8AcumPKYeaC7/mqbUxmVt8L2L5d7kSW6hYyJRe61QlZyMtBOA02+v/wss/rIP8
rIl1AmWuj0AQn0652ZUCPs3iHuH3NpLq6KQLfwNtXaq3qazFCLMSVQ9cNprwo/kNMoOLDRJcYdY6
hcPMeLSYRfvceROmxbPNOdJSTJwe920SjkzZp/QtKZ2Mm1iAm28jjdZCVY89hLpEC/m9Ijj9YE5X
iXH3c2FdSeDHpTdi5IJMyEsu0XcGXIymMxa9f6fgubxDx+RweLZ+wXyeWYT4pzhJcfC3M2NoTQJ9
6i3kXwU6Wn17Yjkcu9qAti7oxKOLdIhYrPG+9d3bha5Q1otgeofccDCfAhA3uzzDzEg0Y80WC0AZ
G4Zc0OKrVtc6hjZ7v5Kww7YQnD9igqy+rYqns39F9y3KQIdk2Ih0HKdGJdMq5IxBcC504cFEyFQg
ZFq+2r7JhUaRQVAfCddZzAeC7IKGA7yMyndYy2JyDPB4538gtIxku6jb/2m5HGEHupjUfZ9LZc1f
5xt8BmBAKeUftKwi2AExMxK+RmXlw/+KXcRUjH0+JcD1knqrvqenclym5J/UTBbsXkew1pov5bAV
fgbkP89QCcwKxPIR87e3wC2G6yR/4l0ldLA7TdenzXUOkZW7kxm4TPqB0lZd4k53/IX3PAAWR18E
iDZTq1dZA8GuuzPgZnF5leujvqnT2LCYTAdicbe1rXCG+S84YPgOZDsN7vQ6DtuM8gYRMTGv1LEE
SxD9S6VjKtf8IbdAmUMjc7lrO39rclnB23Hznuq29PjWRbdn7Zs9nz1terrHTcln1IEREx2hvUjC
d9Rww530sLJpY/9njbe7Nt5GhWU5lGt9Pn+nxazeTTRKbXrOiOAi1hhjuY47oCWnZK+favzTK8Mg
ViM8fjsomanCiEfwDAQ5LcPJhxjLWQgDyTKyu10Cu6rp8BnoUTJf2QXwuYdYHL2LTTi8ju9fM+h0
Fw/PDrDQA+pcheJgouGdce6JN7Yu5nuftLjrerwl0nZ+S/NK4hPM/jSTnucTSQvT3TyQ7yPTNbQi
tTlfhK/fZbK7oK+bPmYEkHLtCK+f67KFPLGeVpvg/M2I//4ltr4tmXlSkhfIfgkKfy7BY8P2uDQH
qg92Wh3sA+93d7VFqAeGHlDJZJbUKn5cRh1d2CzBin/Cv4xZUpvEn43XnCmPuX9LUSw54NA6knG1
zkE0Pu+a4NY9+R8RkYjuK3boufZXpV+3nJSBrvJkK+Uco37DNjokmV8CbL/SYT80y7o3ySHpTdNJ
w8BREktqYYjLed6F+5dwYGSaIEMgxlXcWOni0LogWkhWt+1lkh67GMUJOpSJ2yAeDAHVtaspKDw0
PTArW95FmqoqhuPyLx4OOYBrF2qmve8fmln6H+ZbVdKU7nLrRVP0cWtVmd9/h/2tjoK5bb5aFMx3
oujlXDC0p9cOLP0/hSRNbVW71Hsm/ad7Gd01p2xIASd0tf1fUNIUtjmbJgCT5rNIvxwWKQMfls11
rIUCWp9mlttIYwjjTKfUKj/gN742CevUeGZWtovAzOsACkRpLL9VwgkDCAKbHWz/3tLGg5Xoq9tN
8LUCNgTsUpLEOUUiizeijszpak9GI/fuxO4zaVAoSCD7yOjpkVtA9vaadBd1CJ47EX7gzX2lMbaD
IjaLtLxNvMj+zS053Hb8lxCig3pSL4eNULZHMrLWZ6qBXOp6pCdNHylWldUoejcXR8HiaYyzhT7z
YA0cJ3WnbOswpgNg8BoyjYUkH3B1avdC4KbhqP20DRqKujeaXDyo2z380cTyxZ9iGUVev31aHUsh
Hep6wGd+O+LPBpklZVJv2GXHkmKVVAP8/dCbDj2sNUd2UyCPxf6toQUdLktRNxE58nObHEkWQM2R
TeTBbk+nTHPk+Ww0KQI3oVXvbZXx7tPupOdg7aoAZGbxhxP8RafZ7NDnsYOc1pYlaw9iNhr34nSB
QD9LXp1HkK1dFa6HlLa0QpHc6w0bB7CexbBHWQj5LWkKpVMIgbZ7l980AtiAhk64tqYbF7mayxiW
96LfxybTF376bISqxGgNInPC4Xqn1Jt1y502CR49JrVjeGHb/+ibHnuF6B6tLYxLer61Ba1T1KQ8
U+K4cQPhBN9ar2KCeWKfSF7usnz26owptgYj+qlSCjyw+/qNWtgvS64so83PYrJkr79HtcImWVGf
xxDwjWRmgFtayAb00jV0/RiyRF2zIUOja4+AIXwAnBPjaXcHWYMfk1OgWcFR8zw8IGHQSz154msf
Da3OeKazegUp0Cud0u937jEMDAF+6kB0HysRL46UxAP7fw5kHxjvyyPtGRDiYlgpJNZjYh01mxXS
Ww80NYXcpivGZYWKUdtOCykyy2CJsO2nDkioXb7V2ZjIRs6yvgA4ayGn1/Z1JIJLZtrJ1vyKWOBY
V39OYX2gvQySD0PeFu1+ZC1YohRcALi78htVPU5j/dFvQCTribuz/2PjKsz7RaAPlcy1gJUAqRTJ
BFGxRunN6/kmvalqoMAPcllLZtqKLxvuaDMk7eT8s2YNl8J1G4cg1U8PRZWfr6uT3vR9Z3csA71x
jAzYZtOM/NREUXorY3VM3lR+MxjHHgIcBzq14QbvbrMnOfHpU1ashMDf1odMqrvtULfRvpqCyHZi
Dfu7Cn3sbycuajsRwGDl7kUGrZwhT5DiSYbXR26y/21jd6fnsSYW3SCWnDi8JySneZ9ySAdQ3tD6
HFX3eb6Z7RFmgPNCU4irCgjj2ox70l0OMyWM+dkmggsN/jbNU/fuAOMAe2fbpY+iJG8vkDBvZC9Z
wBdSN7bgmrSoFGQ1h5CmVqYQt7rBsQ8teBhTVsZrOJ0nWaTtv7ZWlXKm6E7gsvmewjQZZbbF/SWL
T26q8jEo3T7Qjm6pZ+9bmBi0uKmL/oKy7ggii+v/sBf20rJHR6dl4FDIneym+nVJXfRJHIPuCQf8
hW5fl2fkZyxkRUdAm/PjrcxusFPTmKa4Wh5GeMoS/IChqrMrHOjF52Zu19DxOOf/JEK8Xd6ZMmLd
Aoe0VG6uhMux8OOuYu0e1nmdmM0Pg8doAyO1KHAMiEjv3UwmxjpneUIWfOrpT/H+DJ7xbrnBtQPO
9cYWsp+y32EdcFYrGlovaD/bSne6BgYM0ARKLEwg3Cd6Y3oT41Q6k7VqUsuTLTAPHgfnzJdaHtmE
c5cF4jvmhIfiWI6Ou76mZOZ2aGYtOdbq7vnbGBKycyYWpAiFhBGpoSROdxt3tSRiEOpra9aSgdO3
sLdLXvi2dG3ovkHkl1SXut5rMMf/mgeoy2OM2gD7+ceCi1KQkf4PLV0omnDTOL5Tk0jEza5xaeRM
jrwimKbSgxcM9i8TOlSmXdZ7k99BXNfDKslvGVZ7zsK/zkQeJ3HYtOy0F+gl3jh+JAAtes8L7eOI
RL4M7Xnd89B1fxC9xtJaYMeAybK+IcJyBSa8aPWbai9FOhYKYcSXio6N2NLq4fuWhndIEOUee78O
Pu0cRThVceuHBk//e3CugRFHi3Uh0eY09dhZwv9QAspAeABm36krlR7YDPRphyYiq56rpkbC2Jn2
X0q0K71kWWiHFGUfnhNINdV7nNQRFj+F4EfHL6bsUjHp2Kr1+++ss1/JD1I8IRYd89q3jOwlMn/r
v/YOMbC3GyP2lMLy6C+fET+T2H3oIJoPrMnEkTslrwesdytn5pqkJ61hsB1iEXm+PsZVYW00zbDu
Es+EUUQanxpAcMDejaS+hZ3TMZvr5bWTIIwno3I3QZy+qAgAb3DO9HaiXp4E0bXkCfslhmwifHIV
mPwbhAwjeaV9pR3AmJBaYw/QEzwsdM19r+6FPqiJzl0jBkPemNhcfTb59gP0KQ1Xi4CXEfThPirk
7DKq1auwvfXRugDQ0yeRjYouBYAFOF9CuYXuWObQTSZTAd449lFze+X+GNFZzcUP09Cs4uG1FcyP
ta21jZXL0QzgSTGnHd901bawF021O1P5MZrm9NKihzVINXABc1OidxZSYOePayALRUajNhk/9nJ1
KYXlohp3yxIC5G87B9JVt9mcjwW8tm0QNn4e/D+1IE0hiIUi6HLiZDE3Ftur6vGvywrdiRk8jCYX
ahXJ0+HVVCkxf0k7wvGzeQ+ituKhv3uEO7P7xYS9/fxuBsiJTVbJNQzJSYfvTX8ZNVojqM4B9A7Z
EE/INVVSwPGY9Wh3dRERhjaQUS8nTrtP6ryxxyEnWznFdiJZlLkYkZNcU1n96fK/td2hcCrebX9g
bPWHlCPkmkMmPH6qydq8yZpZfWztSFebWMmQgQwn4eQ90Qwj6pe2A4lU+8Gy1wFE79/5V6UdX959
6eC9S5JLBHJBEU5sSPX2tsOOLErxywDU7O2KOI5RjXUwO/hdO9nnvESXS6c8/9ImHK4wiRCKweZ7
JhIQGT5dZR2mA+a5YlvMWX/7b6kGEbwfeET6NpzMnm4C9g0Rm3m9uc3341T7tyDJiyxcoliqLjat
7AunwVk2ofog1ETR19omjy02EE8pXa5IQ85IREIZV3ZF/U2viLEIkgKmFf7FhhdjawfZ+qCaWEUz
HTtRiug5mmooLkI9gur7L+E3iSEtlC9zWHDEdSHv40c/TTgibGH3lDX15cm7ypecJ3MTURlllTpX
J5rL34AU1gY+XQGshhkC5mXuX93HGB8yrLcBg6sULguMb51p/2+XnC76mAZkI3P/S4gAjCkMv1kq
hU7uaKDolmmbWYYDiuTNQ1iD681b1RQxoU4PfRHmwDI96h3dmcIV7KgJmURt+Q/xQbY6oo2KckkO
0nAuKPuAFlKGsoi6ociJVAlfntFoqZIuXThaTDlv+UNeJ2MB9D3tOqGw+mENtutPDAJO9Dm+0YWK
n1zv3A7P0HwETJx3KbOgTxf58FIDd2VNtEg4wbJDh7LXDfvKAlXXojosZ9c3dbtjLSu+JgsULmmJ
Ilc+kfXn2zgevdAkDRaDMXIXbEab2iyVTDT5EaQf8AnpgRtr8WKShwQJc0MphakOiAimtsqYfzz+
yKAfC5Tu8rZDIOYoiKzrF/NHWxjEJQf4tH2l/I8fKXP4ooR/ENzdWcGf0l2hydpiS+DflrM8msj4
ploIGnk9kRld0ycbdkgC5c/R7Dr9Q+DrbeWTL+2hSumvgVaTqiZQ+qsAa3Lf/rx76/uBGCHSUt98
qGm9FaaJQCuFMxNbOzITSC769sBjHtglLZSbfAmbbWOxf4tLeOv/PnUDC9LYafuPiQEp+rfi8t0Y
+axJkmRAql03Yx36zw6hy3OUDyMiDJB8QySSLXsSc7IypSCNZLif/4Brlm4c22nAr2oZV4J6qfu3
OezoHsfKgW9pqDNda7rFCVIsrYwj6Ss4A8qGUi6xVIrxThNEjmn1DnEbEOpDBSAhDoB71RvYPd4S
L89MoR2rKV2JNJnGn/nZbt5wZu08ffYhHffzNfV9uNIsGtBi3yYLvvbpkU19d9GavfC2xujFrNze
kDtnPiAhrbi1aatoNGIOvq8YORensixR2ZOLCDir/G7BKlv0GLEDDvHJne45aSz7KcVYYVkzmx4+
veidgAPAAUzv1g6Nk/XpBO58iM4cDHcKev8uPjRH0edEP1Yi2UIYrgNY3/Kx5lrHtHXe0r2Q01+A
srAs3L6KOSFE6K+I43TUIoG7t58YE/OOa12+l/nJnRG8sH5x4UzogklgAG3MyoyDEgMjHL2NJYUU
pjuahpJFkAAWF6ynyz7CGu0lh4n5kOA2rAzo7uwHKaRRHkLXOUkmLuYXou2nVjeUwQIz9UoSnKF1
67a99wVfIxT6SIn8dP+bwEF9/oypCZiyc2oBpe4V/uRAAjlxq2P8k4s3UoEPuxRUmgSOpJcvnSpB
vtA345Ny1m8fzjMhoxRTP2Chx3FNAaMCrxCMSu/E4nKlofj9aMDaH5BZ6r0eYIiephGG0i67zBQC
U6Q/lXIR5/NHE67d0tYuFYDhtHUal9KiLD0yvX0+Qg35UqIqIVfcjAPgKT0utnBBPTArLHs10Cow
C16CAbXYFU8+wDdfOkVJ33Gfipg+dsjG9NIMteZwzHngSFsWC1AxQt+nIl28l2U/uvv/N02h7tu5
GT5sI3LbLV++n+5xy3C30anOte/ezLN8fjrYRhNUbGCIHHql8n0wLhIsMym1p61W49Yz4JwHtwwd
yyfWzUjwyPfTA0G5reRIHr5he7101CFTTF4D3/oi6Qp8LlOzJvJbul1WHzkxIayqVo50xQbuZ5T/
Zngl7g3oaaMhInheR6ronneE6R5NmpTiohpEU4Qwx18/9QfOFNoy14qAI0u/5nr/UpqAG8+K/myr
voE/g6aHNNV6VNOPq0duElKilz7DidUckriulgfhTSY9kXMHED/8f4rqUH2ETCRcXDMJNPK7yEoz
91xzaX2GRFJKo9rXWr/I/CT0DHkiOo1bFWe3WaQZvlzBZOvC/igZTXdnQIaUgPod4MCCc0Iipl2A
mlxY68E5eqjSWCk4AEJy0ffrPI5r67TZHw+wubZvx7/ta2JAsWq/ggPJght2cZOvMIaX3dWRixcd
OS825HiJwkxEYewy7yCVGNm8RkRShrtC0bSaUXiYuT8gxWFNtsLzfXLfL5SJqxQlg1Ja1Px8h4Mm
hc1fK1++NF7IMzSSb3vDQSvnmaa4zvY0STMa8JNR0bx5b2r2/Jf7RoBSRvAjjtJLdAsLkuYtE7WP
0wb6KWu8t/oGprBNK2XlFAsqfguS0KNKzxmoPSMSv7jnY8MvR9j2MHy8FTI+oCBWZq4pDeZKf5B6
X1fUNwEdMab8OsQHLHfy6eSTwPDATmWdjtlN1wftM5pgUQ8KtvZhC5DgGJx3YKlItiFdkai7xioq
93v94Z2ydOuNdunRk1JeG3iQyKAP4Fheca7x9jb61s2IfX1jPEbIqMqHnkncECRInWHGGSNjHYNZ
KiaIMTAwdjL20/DAJeyqXM22JPF/efVp6tM9dJbh9DF6CLWGUnU9i4bgxsyR5AUGb1UXqmVq2cIk
7ool2flkwRlCmcPeREQGofDa4A4eBqCEsX1+L6mymlwesw5KjqwlmXD8KdLyBfNNun5fM71q6B6G
uaSX64bESPJO1cwaba13sjiYoZszVD9qDTmkVi5qifewmjomFC3XxePT6vwF3K5ktj1khrXfLFBh
7W9og9R18J0kx6g4MENMvFOMjkNp4LqEkYTFz6XTEB5Ri8+Wv2MoWsEAv/iaRoOQmEs4OJaDkdj5
gfOpyS+zgsJE2OvC/HiYu3Q29OddWtuM+X5pAIciDT0snrlrtpZCzvionFAbsTiUrhe9vsC91ppI
FZ2LDveGm0lOCkNhnh3fmty93JKS7ylLq0vRqGLu/lnNO0v2XeHNZJwYmIcwMt59JFaJObab+ip/
c6VHOINfTFiOQDA1oiurYJqJet9qHIk6qHPzphjkoDW20RHRbVdKqIUAzz7sfeSjBFuzvJEsvWAh
DfnW6Fm+9akJTqGJfL2YB67pEorhHnahi0TOQcFV5alwFg868I4K6iDktTGc4a3NSl76sQPYkj7+
uaZtF6ukx9iPZDszVoPXnIVjcPlMvRBPHalmuzBm7WMZ6cPlORXI/tM16MWdWn9oJ6XJulv0aUDC
E2OGiT06E915fLjl5lDCOCKAS9Vt0hXtEhP0GwCdmBygBkorG29aEmlWeJItJGen2RGlEjY/qABR
o6ym8OMjtijjWyCgPzMVKTEZV7A9Ftj87d6mDhzD+V+bf0pnqlM00Jb3nVSs2V0mBX7k00GXurw8
B7BBzHHrFrEN8dlOx98yHgPNei0S/9mN182ho1mDbF2+VypoDz7Xfb6RO3sTdc/KiwzAY2NoiQk4
SPCCvaMWsfaZKZeJGsWwkAAIJ4dVz8ZcW2A82Pc+5+l3egf1lcujEWQRLoWmpdOujsMeuv0xyQxr
CKuMuL6+W05md/vfw2Bl49MRh1I2ASb26UZKAERZIQVPWE2ChhneRBqtAuJ6TI1Lg1i78d37iKoi
YEAXsDXmBRmS/32rn65ot1fl9KIgaDeFB8hWlC6dr5peDjalVrpH5czdTy3jiDWV7Fn1e/iOOHaJ
TNUEYxpQdeJJatCY7r9qD7gfCcdFiDY8T4eq33oNJb4lHdEJWFQ7bhOF0Vm88r6/sczOwNZkp+X2
0O3Ht4aKadU7IHPIGaZx1YPM1RIhS//F4u7PrpNRE2nJv4gByjgnYizDtpVzjpglGyvaGaWV9i9g
Er5hkn0FNEpTLmIojieMOJS27QAIXQ/dmG1nj6iJxUBQaUbh3jOTutXiYUhJIKSfJb+pmPwZ+Mbe
waZtmSLANfp7eAaVpnNixRT2Dz5YRl7A4h5XDwItm7Fjec+NFKbfhWEmn/mnprKv4ev8ZltfAXlT
/iBPRXWWm8RKUnv8mLTW1euRnOk67UkOPfAw7RU9+RDP1sOM2uooqg0awkDVXAouuQZwI16LQNe/
5WZyZUxqnJbaO97ppqJXcBBnxaRfUJ3aiKSuOTzxE/1aipLVET8c4BXkxNcXNZAonlx6tchxIBv1
nfy6Q+9WHG8lu8gcaowD/6hktRafxu0t0JNVbiC7rbUESQFqqzletOW7qxclu0VhkyOlbaWASMWR
Bgb/tOQTxS4uWzRx+pNhXyOY4Eos7blioVuVokoOEnMracXYUBEW9rWMEZ3tQU05sMvbZ5+8epTR
h2UtRdFQbhUit5Z98/nwLK874NDBtpBT/re7m/YZhYQqawJoPLzwKfFlUJIH3d4tyED2e1DRI4Ko
S7fDuqfdP6nORsRyT2+Gfir4hglPtCD7iS/k+K8EsUfLOKdUnZ3YH+HSyrw9bsa8Cn/I10Q+F4Ey
UKurdwBWUspwAXhAi7oD0Ol75sg1qQqoPoInFQdIG8+hPMvVsnMxj7h5ulIbNITpMV4VybPYJEAk
k+ERViT5tnq47IxawZDTBvXwVuxmCSjQGT21uP9EEIMA5UeKbOazXwQVkFnonJWg1VF4YOX8Xpl2
YS1WBVrbxBesxp37xJaGdjlRI+dy4YhxhDplrOo19np9Azr/VcBT5R8SmA2WHPbdYwi0Hjj+QUTy
2whvSLZRn31iVQzXqul6XYyuRNfW2RgRJnwE+feRmw+7ei3Ws03WLAH6prmlUj2lKqeZ1oZcY8rs
hHMcGG+Ac0QsmJNVYOl3GmxShTNoIBIlNFYwUMLwiIMIFaPwALuUMtnk26W8NHyAjN22FNVZEP7m
hGTz5DLgfgyj8/PpImR0OcOI+UeAjXEzNWZAU9V03Y7M9xzJTS0Dn3pAJo31Z3/Uuymld+lnvhs4
hJlmqtgWsI3bl8X4eJzG/pBtYva/BDBL7guB7WCAf3ewkkzQ10WTTlgFpDilwN43w6l/2RmnkVgR
uXf65cT0I4MQretpdV5NABvgw51WNVUz8LE/OSLZz6z5CRnRT5NwD0OvjGW85Z8IfmeJwrpOKOaI
tozWB/eREiG7xc/UqzQmhYF9rczGlKYmy+bSR6NVhaU4N2OZ2sstZRfxRLrKuxalQx93BhbDGlBU
57q5sNdeYPjrWv3aDfHS5E0jaMoY18Zzp6Hm/t0/PCrKLh81c6BNi6uVgU9wZEEU/DDS80VTbwBl
4UWSkpe00qWnptEykKU4cJRFOSdEF37UofXpzAAVqk5FJGEirVOAJhrYja9/oj/CtrjDjXkZ9Jg9
ST6Z83VxR4XmPNjwBTwTh2lXGjkGhnuUYdIiim3D2KGpMCuxEmj9Sywel7I4l5Vq4aNlp2u4cXQ8
Dr3YMb6lCNp6g+koG21HYTROOLyHSBQRULC2xzHjQ9JRLIxymSmnTJTTPPZh/I0TpnyduvjJDRXO
py/SWK8qSrw9qAIMluMko/0U/ja0enccqsGhcgWVVdp2DUzBgjl9SdoT3F3N1KMFZvN1CauESkwq
05VbmTkBXbVStQPRAH5zfoPkXipEEStsiC37kOeKbj5PGlKc54AsRY1yGpfsbo2nsR4V20WOpRL6
ndIv7IqbI3qPNuMvGT/8PyLjbabOYofv8KgPgnsmJ0tKTANV+SOt9bPRk2MUcgLnGLy/PDJiyMXR
XB77HipnNGcef/k9hQwpLKjXy1XlYamf7Z9IN15EAzgjN4m+9PKFB68LBgDd2801N2aqtMrpE+8U
PQ+IuJoalwPLHUiRdXKAUuhRF4QNToN8lk9ODx7RHjvrDMt6lvo4JQ0Elg6gSqIeFhW3GKL3nQS3
CM+SkXdsb1fcUcqpUCn7WqMJdcmV2czcRguR8VV4n+3fJZTH3ESMyePefm7BwmPoGtKUitM+fRxC
FWSdYFPlAlkiAmfWBOg3D01xdB3QRSKXCRCPUTJS+BFlYEPGdtPxYMMKQPQTu+jv7xqxQDKldMR0
4EMv1woOjqX4WH881bqpGZkmgVEOs/FVOdFc+61375Rm5HCeWf7JqlhEgQQOpKeDADr601KPN4qg
c4d60dC9+yMBL4fqInO4qZCzkPh5kzMwSJyWCXAvJkiiNU9ZonG2qwM/ReBPZgSwY5xL+RVkF6BJ
JIT0PetJpm0qLjtQe3Y7Q7QeRtSHhmzGMy/2xUC+hyA+8fEJYyko4rObwa7Sy5ogvHdcuNXSyJcJ
vwArgIZ8+rMKlwQn/3RnxWi9c0jYmyW50hhoweG8R21gh+9sDCWKRBM8P1e581E05QHFwJCwy09D
MXBtNwFxfyB+Q4XswgjxhxsbBnGvLKPHbKf4/EHFRhP211rXkTd/8Uptu0O4boSnFz7eeaUwD48E
85e0et29tLjbDt+pb3nTQ42IYux0QDF4vzrLnWLMSUiLvjaDQZRCcCZq80Rq7iGB4aahW7mEVHij
PWSmCC0mbulaA5HVMlENoYYVTfFjdyaV+GiGz3AvqCngz3UabDhkabPnq2jcN1wKUVv1WFYUGeFf
KoaeDIUaHqXcaCMuyEfgUMUW9Z4EVhM4jDcr9RRoKAtsPuytka5PCgSeojzTosm3S6BSfzvDOblq
wYX2oGg51KYhXGLZNQZrWh5d5Oj3uRR0GN/a8zOhZGkD/JHxwrOYShrTlijkVNAq5z4yA5cq2VCi
XrvbZXYD2Ku8Y3QPYoEcr3PWSmv+vW0gpzr2YqRFD93ZEdUTkrx4aSHK7JI/TCMuuumAOBCMycyK
SGUefqSrARp4k9QhE1ymNgQIw0CDHaefB8oN8vatv//rOK2EDISBflHV/sM7hNaIn+Yb6LJHs28x
k+oalka92WqdFFImRlcykb5ex9zIwRedlo9pm+6lQwqaVZUKnlJz12cGQ3mpQspgaAfJNripeXXc
gt9v/WpaHJR/tRRYuAvVtQMY5R/JT29qe0/FjVd7hrfUQDyKs7p6degWPL69yGoFdVI5Rysw4Hdj
uS9qyvO0bZ3BK89+nCPPqjokGHZpLa74UANwn1IEY8ZBGRj7eb5YEpbYHF2HoiNGQ4Ke+r4wU1wC
HeEgkrtVH84nOtbioapSrXz3u2g0baJ6m8dZsFKoonxrpgM2Z+ejyjvxtJrVLllpEL9g8FojWb5m
QyG5yFh/DwkgSvC7GWBXNCrULTmPsbNWha/kQPloclcPSYZfZ5755PATeZWyBRoDu2m95pmiQzlo
/d6zOLu94+cCDD8SeM+ejd62oNcxuZH1pC6ADz0snR80NOM2A7lGzpDdUXPArFBfLPG7kzm46ET7
rTpwoA8EN0bZdFTfOfRJ9TJeSiLMsmTqN1bwpN/VJru59QLYVTQutEwCgPlgyrYwtCXhxr8NJyUI
cptuzC31kmTLT/GCS+EKZSZ7oYdEitLFcCk7HIBmAHchRl+iC/jbJD4ZtufQamM3BJHI77jIDosU
//3ZOG3GuGkxkdfWovC/zt+SA4v5Sb1zKfwCKssXqJqOV9AxoHAd0XWRy2mwK0Jn4kMgfc4+Qi/e
VjAE7GIPKoyGYaiMMeCMXe9y6VboVcg5VWk0UFYNUqBZQ8F5VpTgdepbUoDrpIcxAfwG+RxQrMBQ
9HJX+5RLZq4SgQS7r09VckIWhEYIVrhzjIvnUW4HMHHQekNvFHia5GftlBweAuqvS2p2woPOu1+i
u3QOaJuopMxfe6/APgLD1+P0E5oT9kVxaReklDQGcBjvY2000kTyAV4almpTrQWmdr0AnudE3n8E
Jbq8F0iuow4ivR5jIaupJ/PzV1cPxSgj2ecaIJL0yhN6idhRRNAUgpuDi6dwvvnbANN0xCOw0bLX
79ry3bf9sFK5hTX2yBR37OPUpozMb3Xw8MzhgsJu9Tmd8o4Yp814snpZDMSE+JekEXgCvnZM6Mno
9+3xbkPX2D4Q6sR41tmfWyZF/czjNvkV3QVQQNFI9c6hRIxnAmOnRQSUpUkKctBiTO283dXOX1y2
PKn2dmvpvIPtrwxDzjrMBiVH4bb/ByEHKo8I045+6pBw+ElDEKKkSn2FUKBT7q5hDOmZM4vS/xfx
VwoSw4HgJ6fgpNTpeAOutrhMoVvOJ7yuEWaRpyEYUpmUMilscndTqBQR5BmP+y2YUbT5iz7AuiDA
TRcyq7KWo1Pd+5YRIibbwTuGKl/UIiCiwtn3Ry4wehrUptrJOCjHibd8qn4PlZQlmHR3RXeHp6EC
O5rfFRrxiNMZQrv2VZZtlDElPRIDiu1shHZvPs3tnK87yqw/usESNiPGs69jc5/vi8frB+bC2ney
Fmkow3Gb7wCkOlxVJflzhPGG/kmYuqFpaRkiIuRRuvZUgHtOvz9ADyGaSZ0tclDuR9GcrH/1RjKs
fXtCKtFbDjicNbDQTkKWopVZDfRQa0KxH4/ww/FOKK76+kcP6wU0jYl06OYVcfyWBSQHUGcWr+EK
955pU/CymhU8Ewhgntn8E1Y9eVYKptMUN3j2y+ToQS5gXUUlxfVrJC7TA1lDD94TVyWGazx0ZoK/
Tlzy8TY0b3XBlGZwF/gS8Zk1Sdi7SHyO2WKJjtTMLhP+BV+5KL4CjyH5LbAWsQvxZA2KUhOdL+4K
mjPi58aCNkjLuHfNQzXp7SMxgaCwBnhfHvgWTmi/OZmqflEk8HNjI3knahWXyOdxi+SwDKDKpD4F
lj0AZczTv+ckxiTRb/eLtAmtazKYBN+Bqt9BMu2XG5ZDLN2UXkK6EHjmOSC018RaK/uDmEXjTTIk
ILsdtX3Hr/GshxxHW+QjQU+T0GRVchlguTtOcnxIlHwacXo1Llh0HUDIN/OP2G42PkY7Jckdbdoe
l28BtacSd+1KWtd4jAywPTWu/sY7bU0cu9c4tBUEoBQ6ZxxO+5RxiRAvP5+OlRkHhhtFnHmd/GyX
nQeZzShLa67QxZvuZgQ94OiuqunK3F4wHDEZE3X48i5gSobD8wltH5h4sgQKy+uJWE2fs28eP8Bj
U0/U6oXnIojn+S22FWDeeMvUHDvuiOIvoJlhNBHs0jozjCDryYna5uambf87A0JA2zGAZNlZV4B0
Ow56cdpHVA6J1VvxDitvopcvRLXMtSNep8SHyl7aN2R2T0/Li4Z/e7Kxo1NuWkm6O0boU0iNn0z/
KSQ/qGWfck8pWUtcjpiYQQXfF+3fQKP/HcUhL1jm96PAumAoU7GWSLyYA90kH0Qi3VRl0ZvrlidI
kPA16gOXWT65LwMkfA+1Pn5QjD9wFz7zpHAhcfBuvjl8ovWZO7HTUwGlXPQJLrTgM2mZkffM98zB
EyWoCIZpuHVK+iVinZ3ddB+/7daKLqvbUEcbBVCtaRca/TLJNDJnED8SpGugXa6iO94TAPaXEgvH
ULhEfZH0tQUY8YyenKq5mbmhECke8cc/+2PPizKyB/i4eWCbhyoMX9feI8qqAKmfbb03ocUWamrt
7CE/kPouWi4JpNI7cFo9Ine60GD7V7pa6Y6Lw2O/2+TgxrodW2QKq/YZYSuMT89o2wEdpTZM1zCC
RP6KdbG9aUH5UARvF+iJw0UWD9ZAVHJlTm9LwsZFJtuj7RBVaqFe9Z+1M6/kGoD/JdPXl5OfUBNd
hPZWdojCFWOiq+/phTqH2x5Hd9owe+WUcD2CZHeOk37LH3iIKojhBAC9X4KIPTQJ10ynb1LaqwpR
VZHas0U4Mu1+yYcfoZMGZhyHJ4l7nrHd29KLhSQ5zg/Ahjj/ywYSFYkGyjH0toGsvMLJmqgfNnLn
Ht4g1urUmiHtgxtN9YUGduYoXbkyx/v/9UBmnLE2jTGqInEO3iGL98I+l1QyKL4nIDplBBnpXk42
nKwahN+iwKpT2NBFrwqqG8tXjsol7LQQVNtRyTIVzleewfG67oS3eja+FKsX5tdEAVsFWcM/ltKU
tGqICmMco+rF/iupA4aP1CBDiHhw1j2ujhEH4SmiEH08HqtPr6zBuLfeI3ZyMcMvoQ+XbQ/a3AbK
NhOcpw8zqbtldlkHQ0TH4o5AkdZFYTAHmx0fuilj3rQx6LMgooPSsRuVVR1NKf6jcENb4ISLwX/Z
4ZHiAa0hbxyumvV7YZxp+WipFuDf23PVczHpksZSKfGMH+U4Kt5z9fyp7AAnmodNHHWl4fFR3Bcz
RQVAcdlMIkbfstY5ysxFhztsR8D5HiS5hpuAP/TLXp9VnTU0Kezp+Avd3QHx/3IUkuQU2EhhYRfv
jE97gpNv7HSCiYstwqTwVxMe8Mf4QhZKK9gRgclXNX/WZDnk/gxE4GODE3D06WZi8Q+CrsDNJpyi
I6BhpB8U4H3w6SwzdnMz2SkGH/QNLm9QNT8mFa95VvlM9EehrUj5JqqS/jbzqSUVlPIbxyGpbRC9
h7w0URa77IJrUFYVIwLywdf+fvMk4YJq2tzzcnkpRReb4k9gLKa1E8ZyySEi1HWiV50SLt5deWip
rIZ+kTSwWeuDYnPzg66sEXA2p8A5CbijnP2H14L41ZNk68X/wht6557tjur8s7+VFQNBy6ww+wJU
lQKGJhI/pSgPmvdHm3+f67Xnbg0h02ax6X7YWnT3rB0X6QR9bc6ulThrDDmRWy2dtAvaSThXnYkR
qHtvH2hZSGko6SiSWFLgZLvKLtHjVVH8Qx3vmnU2UWRBsQs0lb9yaHdoF77J2v+1i9FrbdOcp0ST
FUTQ0QfZ6OhNeLlh6qAYBxBwOQ2nkWdOSJPP7wwSTTGLbRKCzLqXu9FGtFPvCiuacg2jSfyw1m6L
cv7A6FCiDmHUe/jGvYssghvLRMFEssTSARrabU3+cn0sdHUmH3xSeoO/PZ/C2bMZ2Op+OiFBeQnX
SLf82GeO2PsySXdwLMKD7jaqv//hziroVxgMG+VCnQ+UuE/2Alo7suIM7GegBdK09Q0q3Jh1UrMg
wD0S35vYbcVU1t3rzENL/92bLHI/qO1A1JNSQmvZHUnbHCUaUQxF30RaZ1V8YSq096TMbEcQWQ+y
PGa+1omvcpy8YZFWXciIjESolr65SH+3AjJ3gvCAhyNSIhlCFQ9IPfWohZevi22ZpxEI4rj74V/j
UmKp0RDgu7EFouMzYuBlJ39fbsZ58rcyIwo/y51gqOWlT+aBCd42xUJmOsKlTYLjhgc9qM0XQamo
1zHNKWuDl6oTByhBmGXKdRLtXQmbxudiQKqQVrXzCBqmHtjysift3p88wAEsA6yLdGu9GxXFmp96
yCOHdTxd8cTsEGXyLp090ZwhxYcDZ/hh0ejMLEV7/66HTTj1ABz8tG74h8L3fasWZXY8tCxbiacu
QneM1C5TyZ4ia1V+1Ei4l9tWUcixDbntX/8XqMC+6T5jZPdTzdxCJwtcaUQEmR7Euz3lf2LwOt0x
OpKYjVwh8hrzr9Bp4A5XgoZeW9dEVYvwV3OdRhlvWE6giU8IiDiiaQC6gISecMBxMpCs8sEnRewq
p/t4GoVTG2poa6+4hKBkdzGNHI8HDRz4uKkpcPLcL8nwQGhCujUA6StDVvYDqwGAU74bhFbwBtBt
D45fHLYA3s7h40vxXRWkGvt2wPrP054WE1uIHZe4Ag7OKh5KGq/p4Jeh2BR7YVCh3T+8/pAofRi9
tOi7u82tzORp1wvKMhC3ld4tfXb42zqkcFDRRqcKZXnPFZmM31FkNCYDl3Upbgl/V/Hn4qvxMfWU
Pbi1R3gHp9BBwUGm+D5RExkD/oDpXtbKjOa8gXKXRN3xPMRfLIsHzg2UA9t1SfdPkOS5havWeIU8
DE70Ch9jWbpx6fi4GxnW045FTYuARN7xGkaGKvB6z3kQLWGvDZ0PZLfMkVPy/qiZW91xzPcTSkk1
h0aC4hybqUrzxfcd3aNGm1igUudxLOStccyreT3Y+IA6EBjTkk8zmkVELX5WoEw5v3viS6LIF9j9
CSkgqsGfhcLLhbV4YEF0m6CD8RAc5u7MdrdIV7PxBQC77kIsMjuzelRzzmX509t+gPfq+z/Qd0FL
R9RSru+NLMjgs6OlnWjBL3ili+cGaJHgILK5zWsW0+acT1WObfm1HB+XBFWMdJJqxEkIuxOSwqfG
IeTm/jqZ/mNmmFO6lX4TUbjU7+3+Rhfw5iR03440gQcIXvzJzJ7D+/HEQQMYGH/nGLU8zo8VWW6t
SPGyETxW5UwhkZM1fwTIzxG6kCfFedYkdcunLBMgQloE06oPqd3rhsqPx/DVbDFaVvPc7YlTMdfM
o2ViKRBYrBYgX4LiIkPpxtFgY0Q9dzvtBp7ONgFkyFavfGn1XWBVHrceCrT4NVNMXJlDrol2AwHv
49VBsnnsvmnsdoxamucJ7mdYGVOrrmz1PpmD1gZ614lzJ8RcKvvRcgeBEBLdrtT8bxCJjfGtA3Ku
824OfuNkKiqJsP1SGOjabD0BS4yU0MvH3vEcQoy78BJUNntEJuEl0x1dnZGXADrYht0OEjrgghIk
J0KSGA8Z+WX5iXLKRpJ/k0FCuj0kit7dgripTMzBXB4dNiuAMCTDV07n5jlyCEZWKwPZWxt+niGG
Q9UwE3BsEtzYTzP8sgMdA2QCoemBn0Yb0QQyHqybxJ8W62LR3mczl2fqCc19hIEidVTZU7bl/sHs
LwakdkBiXC44UZR6pTxw0wDskuhWu9YZuOiesPzdaDvU3Z3C6woUqEKh6ZtUZzrMYQsW6S9FLEui
Tv3fiAYGmT2CZH/X2NeKYsYu11EBZYSb3kSJxDC7OlRZF5r2YgYkrDeRSZTAEIqYJS0i3lq+mSP2
AWPZJSHrL52MxyyVMQxWXqom4JSRWt5ZpgvNHsHYp/lAZTggCUYsa1JvYiOV1EKcZQslsEpuDpTS
hsv2fseGfeyCW1OmvJnG7QkdTCoId45bNLOLQew75YwXbwftnQBvdbXtCZ3uqKP5xZ4SMpcNNUFz
O6tlAJ6+/nJsvCRoNhgBiyGJLHXY7aQ0nf9b/gkIhRZLrlCOOHvnM4pgJd9EkKX6Q4I9pk6roOFL
FHTPrkL6JtEN/7x+3uM1EUoO3FCH3zK+rQcTiLBuLFHzA4ScHrLywTk+MiR3IfFKHQqAixY/SN6m
h1iFO8IZ9ADbTjJMdlUa47iwr3kb4Vi7WDyMcR7rkwVcqyvAysEkPgO2txDzaqcS00ET3IPr7XK1
KefzbfradombDW5SFnJIh/34zg6Jb9hr4fLghcLk94Cue4QeMSNHhfe1c7A0eUiq3hPGEFmxIOzx
+U3jkP5ASFY8nmyvchsKBsmT/JYdzySBcsNtlP39pb4nnXyAeutdAhLT01l6dQeUj6yn0xCaejZ8
h2202Oza2lolrP2Q+9doGjHwW4GO2Qev9IzBqg4EL2jTcrbfKVt0WXVF0UcsZSokA7VVm/YwoctS
Chp3Gp5YEP4Ao0YCg/30EynYL16lMgKq/ZdRBPr5I/ugB6oElGv8ffasYxelpeL+yUqeYBMvGequ
NHeFm0tX0nxbrbNLg7ry7vyfsu7uP71BvPyQVIHIEi2R8Zduvrp6qwE5bxpcOLUrx8/QEAfmwMbB
Ti8JkXzkVuDLKhhk/NCri/yQe1sYnPuEeRuOJneBgR9/YsfxGfwWuPLsRtSZIHgAKn2vouuHKnU+
UwZdVlyflDD4cZKLDJ71HLR8rkmyitPrXVaN7hqmYNIICfd4IwnEmcEvWYuxXezk9rCNsTA0RfKg
ISWgl1tAHA1I39Aac6pO/F+vYrXQCFojSEI1waOFD7GYpC0aDfubc1b3tNk8uozkglFuUeY2nVT3
A6rkt9ij84iNjc4xQUedG/qCEOIOgWnu36Gldh3ZF3MpiWDkFrEo6H/YSZLn0U7Q7AbhYcwGezj9
AZ9ZyGHEFHrGy6g4KVy00aT11ZNwKNmp68xMa21zOctrbffdlim0xNAcnENKTd/18Hch5r2fYMh5
lkLRzppfMdmbGB0zvpf4GGkUQ0eFz6FuX7Zb4AZ3fvePQ2+rOJkNynMMnnAGO1B99bbmPzSV8QZy
uSX3hp1Ahp2NK1lAuhKWkUfWgyB4jozTpPbny7OM9lRYGQcmd8qOCELrFhZ0FfHQ8Pg1zQM10cuJ
dFj5Q114I3hDQWfysUgsF4yuujkGWHnKPvg2rV4zEgCk+PmdW7gIvV18ZVW+UDquzv27dh0pLSvO
14YpFNXEyej+MpiYOZn+fHiv8rlFVufBXpqbwhlVGowNEubvOsf8cae0mdIjO3v61PSAm2HjFsws
khyJbKxWwX2kYhpSkioNw4yuIhptJqsQOOFmEj0I5iES4/vZPC5dgdx9YaE83/OXlHggiz6XLdiC
w+WWpsLe1nDCzqW7eOFRhmQZX8DmrzsDTYl+6NhlEer+UII3QGY90u2IMH9nQzsEeeWg2Or0iwX9
2BU522yA/UdyKI6XgBQhwnT7x4dKyMOJAfcUGUAUGoq3t4R6ObLTziz6n9vAfbfi/GprA1uGLc9p
OD6pv9HmmiCD7mKcSXK4tIjQPhJ9WexFFp63Ep3cyA5+w7mP2qA/gCuOx7pUR5dIeRqB8E/9z5Uu
w66aWig6wfH+bAoAx3I1ihDsY6HAqlTjrc7L1JdyhjsD8ZdVOFXw0WCiH4x6tmzaXqsgm5zeuHO7
oVci+3qu1OZB49MgWMW0BzYIdj1htp4ntV6AIx1yGI2TeJRvcvNyo7m1fwhqgNdFvnTinMTcOYca
z3VeiaW0PD1qqyI2ikwPEA74pLbBRJx8bpN9fHXAyfqYtpEAdQi6b/c3HpjtYt6FFlpVc6zt6+MP
p9LjKApjziE5cxb9XnfGuyC//UX4w+JNUX2PY4CkWUfWAGJpeev+6rv5L3VoTRrIOOuKaFVWxxXd
LYkJ7ClrIi4qy4aXA5k0ecDz645uXy5UFUq1h4r06Vsr9w6V0axxKZSUcAYVcr3AVumBUIBxhkun
L7r9v8Bf4XzjdrAN1gAR/EikbjKqEBUlWltagBlBX8vJxK37jHcUeGpBgDMz0n2VObgkx3ylKd2f
R794Sx9y+x9He79JMed7m1OwcMgd8i3m7an5RoLtGrYqoxe2CFw41sklg+RV4HprNjyBBdsRZSkh
wmmHUcLxP7AKRn3Tx2MVa3eIJ6fU4XWszIqUsXNmRyiyIILdLTuuWVXSGKYiEgeIdHVqEyYjoqGh
TmqDi/EvVdN4feY238OihJo7bk3R6MJO/AxxtIAfmsqNnXiwLT/G2TiHN+/Z7wS9zfG5AaMcufOy
TwZKo2dSEqBI2Q7lc8URSlT9KnVfhgyPWy5EWFWAYTzySUcHMcv/SpDT6fLa/QsfQ7aFxhTXzHP3
U3bnv/LGVoXdn34FcI3h7DmTGse+M388n8aegimhT8TpGk3dd/CYyoZ7exjb8CwLuWDCNzawe2Xd
OR9nBDDlwDRK+9DCfFdsOTpWeLt7nhlpdHvZzqIyDH1XS5XR8/RAhV7vZMJKD4pO2r1kSleb7P+L
L0eIPiEJHqw0XKYm/ivPxLK7V5IBzIxZ8RItPyy8+krIkD75XPK8RuJqbZKhmJUMGNEgX+FHCf3f
B2zslMF3eY0syGIGJ5J8RYIyHI0cdwComVd8LhkswXE4Uv5I3HQ9OandaAe7zvQaGm9QGFHtVmFN
gzB3ZJlesT+J9CWogWk7O+xzYU9vK0SpmbGUGoPMlUl+BknryXJNaPxVAFUGLIRKv7gdorHS0y9C
USX6yY2VjQmCF1Ktz2xJqWfldML3V64wRLkNS1fBwAM/4e6XtUXQkrUINNhX8qTvWARK8NZrcWPL
8nA6+ckbY9qHllHRPplFTMFPxmxSQSWbfVG9qiqsrrMW5RCZgcNS3Ts5n7ymz2YquB9u5SLs1xeu
VGO6fQJH2etOWKrXBYMuOiOHThTJWjer62hSbucFHmLx/te2FvJ43Yu3zPqob23b/h8S4lIo62ic
897HmKEeVmoh8Ox4O3h8u6Z1e6LFofZU+Glef0+jwZ/NixJ4aAXrmCEzPoNk59N9FYtnkDYtN+wK
TnQ9tKzCGQexlwTKwcahXk8mmfVF7Nt+pUh0WIKK6N9P0kLG2MBk3MmP/B/M0oghbX/gkaysqCrv
ts2mzs2zLtvfqdpIqaFrXlZTZVsPIgwTwT6FqCysE7xpwzMA5LlnMUUdRRwUCcW/gl/2V35mC1WO
F16K4Ea0qVCtMB8Z5ho1/WQbG36QWskjIfZSNSEV+gYlho5cdhYXuaQ19JOlM+VWn/pXHAoso27y
GfVIuuo6CAvsTGE01uqysUYCRFaoAx6m9vftdJc0ZruzZJFvnV2Fc6Ip6ZOMXylAXAID2Dz71Z1V
UtD4OfB41yTITbG4TV6U1dKD6IVFydVIk2URza8yE019y2CZfNuSJzVURf7h34SEEayTbVXhMbi1
qql6B4f2Na9yeaouVJlaMuvTF1/xHAs+mEcOA95gfRzR+mZ+w3NL5f9/zC6nIBFczNdt8xzPHQHi
7Jr0XB46MxpjgZQqGRFjQSIT2U+z/cBENwdpc8SBAGnwhyzeDt18U+z8GHaxnK7azOXreFNM4ytG
LRjENlXvEYo2s66/4niOlES1X5FEmW+Wfz8JOSzcmg9VNtFQTAeYdaI4A/5IPs43EU0KZ4YGxyVC
EbiBJ+3apwJ820QhTEpigrk2E1/yho3keR/w9sMR0Q5OzyKvBkhMQ+TXuR0gM1wLXGEWHLQ+46LJ
6IafhZAAdjYc0+Kie0aMnMdfzAGba3nCkSpS5DuYQ7xWQY14DMzmxAJf4daq3VxkzC5Q8ciyHuov
zyutOPYCy/+ZhRHFHAfyLukRQIXaemIT73NtJLP+10D3vgaebfdq0q5vl6ym2R3GBPO2mQKwpudd
luCVlG29tHiXWQW3IFEiER64jcuyJ9pxHGF8+8Y5b6lOsQYs6/O0vYUpl2fpQxsIULH4gyzLZzh8
4XLjhXLSM7xFn9vQSXrQbZ0o4GO5BlWSt9s5hKaHowetfIYTyIFZfdH0OdioBsczywGQ15MHV21Z
fLVCf4KYzHR6CgBrQ8gL2U6875SXxEZ1nZd+NeCKo+0PW9ZRSadMX6CSwlZR3oe8snmhQ3bmGgkA
Z4DG5mBsnDwa9v9oiiY+txszdqVfGQucuKwnAZfz7StHPNiHpM/CN1d3nkPFemLYFh4ksfyeU1oS
OWZG992uwFF3xU7l/PRvRT5gQ7MUzABSS4Tdx6Po/+WNLFYfRGL+69MZ+qD4cbwCWij0xkMAF2jc
KGL1+UEKznBut4EOiCvdIzLY8Ni263BAbvFMbtVUSojR9L0+i2Q8nKTM6YRp+6q7Hx0euH0QCjHp
H0gfS42aVcRdA78mw/6rY/YG02ueTYyBeMYvmQmXz3ih74yk+plE/k815dgDjNs1NTr5Et20GH/k
Bz7SaUYpfbL+JDVlaDVF3Y12mByT68hGhD5wkhoE8bVGNIsbY/eubqMXRQezBsx+e3aycWB7Kr4J
PxS/3ZO05lK8xistUfuDTObWKmsGCUmV/37h31Y/HmC/xOEtT8cAtzkmUAJb5W4Y7cbFU7U10uYs
AvKouPMnLmjqUj+YiXVD3d5WvTK6i8XHMHgPnA5O/92QU/c+xx5mue3tx5kD5ID1evPJRjqHDNn9
X/Lxi/F5Or7P9PSz/9ncMq+QiELklHBiJ96RORFsDj3zdXEgn9zgegxxbD4QAUog4Oyvi8IAZSoB
h3iZzwjmZ42U8urFVKj3sRbxzC8mnA2BA2FPbJH+utte66TLpQ1Drb+TN3O1s51/3o6RjpSZ5g8E
aDVQCrW6KwvjFAj7+AyDICySSJ7ZkMZm9VlyJk0U00xt99X1CCTDG5oONB+PRzuBXrBc/DPMWa66
1NDAIttVRjrG8G/XJytF5W2ltW0E0IvFCyvrRCfm1KL4km9mu2LkDT5ebPnygsmeZAksiJuZ4thO
5dnFINWNNCnDjaPCsfNfCUfoseISy4nMiLwVcncmOY2goAScX5vRPHcfmCrod/xmUImlp2wWb5OV
AvEfWDKJIuci3vJtbXG9vOKTLzNGkiRPF2uTA2rcF7FDvlVqIte16BNzV21f0Ql2ZnXrWhNKS1QM
rEunTVN6bqIXNb7ZXiEBgGs+Ix0USJWelw28B/3Nhr+A08OA55K5NPrjm0t7CLBBBuCsfCdiPG27
i3p2zx4fJXGvs+nFWJL4+fH6JGzo8VM3rGg6esZw5/6M8LA3i9NYXQZw/jMKGEXMyJja8mFr70/6
fzLGZEzbivcQljZDxCn85ItBfdX9jPQsVi1voZ1gq9MHACzX1AXiOOx5hkxO+Xs5u1EayzkMzh8R
fRJ2ddnwlKWEBoNu7Tlvr2ft9oYdTvYkEyYqJ2TgIZWJtXgCkhT9QxJH5Rztviyamaz9onOnBDvJ
Eg/Zkp+qZ41EbLg/iX215aj+jPRRmChb3I09MRduvubO5yPtfZyTdJBsWSeoJFro8DFsGhsNFkmW
HwARMw87Z7y26rUx3z0QCxBRiKlVUAb0t9VS6O6Tvb781sGrZyAP/RFGQPca4Rq30j+DUUm8WWEa
P4H9MlB4i50ueDYT/B6I3sfIu/leaxGpy/4ywha+SQj0PDfYhmZBU9WDK87KKv2J/T/R0/NUd0mk
fp3/xVCh9jjKwsmdBevTiV/r5WIZDNQWVBbVO2m4aJc0NttuUPZNMWO+4xmgHxGIAS85GX9GevJv
7jQGFURhb7SwBFoNs1i7EIuUo2dVc5mVDGbBS6G+7AZWMENyFvxsZZRiVe0rwb4lbqTl6IbCSM7m
n2D+ogT1rUcMi3FPTiiLJi1R5bvIKNzs9EHPeqrTelP5LUQd98l4+OSBDnbG1I6nGEjEViWLKc72
BLDU+TJo29o/c1KM0BWWKWezz/vImMTU3jJkU2EQsTHYaUUckJ+hYx57cVdY1ds1tZBLGBpTaiQK
Y0lqvCk1mRhWw3ClCQ9176K29lGFk4kHrLEmNitRfHO10LTglbSqjTVjVGdIIi7HFlfuMoOyKZ4X
YKZdnK2THqX7/qIh+sj/QAS9XbIrMsiQjwyM/SDcSt9mqOFJRamLzqSQ2ctQXzjnqRjqd3jSJ/la
+Ud5dC30+VVtsOig0s4RkbeEAI+8ZADUHUjpHsVYKDgdQt785Wr33Jm4HwlgPdxPhjBxnjixWugD
Rrif32+8CJFG5BB8fs1zmb7txu6Dmpqnps5rM8Qrc8vOEcY3ECOWmyzbSrVrRjHFDGaK+pYWcxjw
azSNIRV1Fe8aGaV6jxVh72Wm39h64mKCAQf+9ISBSvxAscyzNsr3H1fAFUJcONcHOjjAWt5WinVP
fKy7Nj4Hw0wQgcm3+g6qDsUvIhU76tDoGsXP9Bt5XzC7lr+9P7J+L+0yWUCatxloXOGHVopqmBSl
Bjab1Sx4GW2JH43+nFF/kK41ZPnDttDzvRAONrSer0aKvoOQ65CwYfEgsUFl198aD6xHXA99Uwvz
B1S73QAHKUNlM5jZ9s9IwCn+QSdB70nMiNrdTfUhQbjiXfBs4IAT0iTuh99qLPLoKXAKNlf0XAXt
yFimxHMmn7rzWJvEyS0+eXutJDPuLKE8Qh3b0+/x/G9PWgVrNV+EhmtMkJ5W6ppSzAyxFV00XG05
ZwvPIrvOjEbAL9SK4LUF+3YNb930mKrhcjylJQQIH7RFijFzWxI+6GQc725ah9tcJvtOjeFV2qFz
2AUHI9wPnLzoWl+fTyQq7ID0n57H45NE7w+20lW9U2JP7Zww2DM4IO2PexdS1sv4QrPYt9yxsLfN
b8uOpY8d3trVPIoZRqYsr8pIWTrApAb1GpNAREgwCzxnoypyktuEV3AHkcq5HUdBSFLed1+7mia9
KtqNQzC3Otq1J5cN9g09ixA8pUvFSLN1AV5ZYA1qO5Y9nHwFS0tviNVuUWZIgOsaAlQudNZ1d0xJ
PU+sdZU7oIqRR1q5IObjECHdgXY+cYGump3NF8V/LJwMlRK0YoToaMZW/FNHvah001E7XhKkDbFY
3UY90zDoOGJeHrdYtR3XmTcbhWN0VNPhqmpaAXweyJ2q7Ojs4afWZ4H7LhRl1viRvHX7K2A5X4/4
r5lVQ9Xrv06MJSqh2qKcM2VgFCW70/cI/Tg/MKjTnXd0IkYNfBj2MyJ2j0sRC+4KPW1VEgJGxdRV
gYJBy1zFiig5UDNPOdjoIolb5qjYxcq9BZKC5gR1wJ0C6DCY6E3x7MUsT8s5P/5SLjID27JT3X+8
JzxHDwyYyQvgjsXMBhsTOwcQU/+ULQx7OcqK0WzsOUMv+3lB6jAAsSbb7titEmd5Hz8KdGIBjIlM
qkTkrc6MCcVcicTcsYvJZqrohqQrJQwIH0QTdINPHtmotZlaLhxHaWMQJw+5XQBGtWsMW5+fDYLG
srDY96SFvuuyKsg8YSwhl1Evb4B/TJ2NbgTpCOqVdb0BXAXB1fna/s9RhswQ802C6aLsWZbOYlAg
dfRHle0s9C1jkwJxnMoXdFjUkJLHH9WJQOzQJA2ZxY9IpTEzsVViLxPpVnAc5SCdPfBW4l2XHy1I
TjTCr8oiMIFh/pnZRW94/cRhWzvDeHaau+7nqfDLAz3/QxS3QKch4s1OMGwf3pV1ruQ92bCVEK8y
hpjYq4aUITxvRTG4To04/G3ZdJivnODS/nXJ4hGUTX+MnT/teQ8Oq7MkBs5nSMiOeKQ6+LAENcAi
BlR4tB+2YflIs2/7bFjmhrqFA2b/ItlaNEc7E0mxmLnwbZxa/aN/9G5CUkNjDaOmrY3JChHgt/wN
OdJOJ+Wyskg09R0f5D3co6bi2bK/+WrwjRn4C2AJS1MOCrp+0Y5sXj90B/+lF4YzGky7lWB0A/YI
/2gvuEryo5FxJbuyZUpHHrg/03Qmg++BL0hFVx1mM5ZlxQ/X7Rbf9lvLwfyITWtRwydS4Ya3FbBe
y2U7qOmLO0/a+u9sh/AlsCxyE86SsjBNmnH1ir6g6b9NmvAkEzSrYH0lTo9MTNFqxRPbAJhw+pHR
OFtheVdI5+VwKgSow1/uwk2908Rm2gpp8U924eyYuwwK2qToVrhf8DP5Rh8+Z4HvKsvn295P5yaQ
ieE7suenQHVdz5XBsdJQRRhlpMNHTGfLzhJfz1Wk4A9FNUcjaVBSd513tmLeQ5ncL7UX2w3Eg6Ki
A7Ircbb2bHc1xNIYq30a8aG3jPEnBnmn+63PHx3KVE0wmEtBTBeDdEWD1jSQ+5/AEJIBbWaLJRp2
qQ2f8jigJGrofJy6w3qJrmK/hogVE+7y5TZp2dSSnUky8bSzO2f56SdGOYsWsLpGh/UIS8whas3o
BZIq+SxHh4m+dau5W/D7py1xmy5lZRvCJu9PxjdYBST4GZv2Gq4mOznch44KYPP5hRRr4MM8kQI1
zmHjbC7S8V7IqtEenjVX4dlLeQcwhGmV+W8TA+TdfwwjNSlbGxbrewrSJ2iPfNidWmTOm8BlhcfJ
5FONzZv9j6hwU8XR5D9c3UyDdrb1m7htn30mIFezihFjSGcMqwZ48VrmgI9jiKcC5rNFxlHC0AWc
zzR4nHxNMGh17xtdEP14oYZRq6UdfC6S8xEG4vMt4D/tLznflemhXBph6bTGFwg4L1b0yfalNdFU
OqMy/YFHeIf7oTzeQ/mgLzDUlkU9aAFhvpQt7r53zfTYkGbv5sLIUM4rrOJgI0XwjWxDU2GmfUSl
k2mC88X7fDX3GX7+Yd0FsVnI8LrRFRmfmyDRd85DJyA9xmkT8HcJDp6s+QRC5QRArE+GLCEBIEPf
MIvjZMQEHFyAthN+f47arzWuxkbI4hjlCqZbkWgPecrQENVHYOTtGRWiZRqH8HBG5A5h+m3F2Ud/
qm7MKL4fwNksy9s2etLDlohvLUFiVTETfaDPD7C6H8rP9F8r+wWI2RRJvvFVf0QcdlEesfbFO7fL
2v8XtN81TIksGf+aq5cUTRLGiz527Uxf9o8iMe8AtYW6wQ31rpH9I2EXX7pijzjSyNiAbJNvKecI
7DTCUGaaYeoRs4PWtZofHjqY4HLPJ/8HZjCoHIxRuWb+cw+M+iUWA4DZzm6FUNNs4hxoUxsUKxcS
pQhntD8OMesPm7/Hxp3+rNgfIoGdTm86VLy2wi92JEoC2BZxpi2GSA40888jKCZziMhEqx9fZG5B
CXs+sq3gzf8UGC+NePFGfkH0RhBkg56XkbznmO/5xBcgEIMDaaWniALGRg6t4DDzOOmQ/m7KkKAj
gsG9EqsM45FejTFcDVKIcS26QJ+hkYuvEtU8tOpDdENPAmay86axf4OTm/Tero3ZYxUjezYowsc7
mnm8af0ELP4e2VhG3Ci72rHPstAC/Oz3AWzABJurYn8bxFQehqhWRhtyl+kZ05i54GVhVdZP4nG5
BCieHlEcx9fT7PY8ErVJb9QAM84GNt1zqRgGt/93+wxgxCxGCYi52RVpvNJH7G0kdi8VHoWjj1il
TtzKdZT9/y6wwun6dKGWPy31QJukYe+/PTaqHqLVrcor33qPkSIUArMFhDZpv/GhwTUkAdnYHiHI
bqTFSz2Wphc1AIntKUitFkHfw8ao1WK6OesGrGvAlS4wkfH//d8PFeCkKgmoGJQidDM2HnRQIRya
npom1XTHssi0cFFbRnQ8Vq4mNey/WVY0a3hwTcYCPwR9u7tL/O8yA1rPqPHDQMzHTg/b1Cq1DCss
M1Ml8jXRsRj+MwLOgYRT+lkaE0bDRGDNm9jwKksb5iDGYQ0xJrpmVVc+fUOxZ4l/Lm3ABnQHU2Rf
zDTjAFGKndQbB+c9OEbUFuqMmPOgdJj9GmpYnBffswXHjYyoyVjUzhux/wVDkBKM6MuPcpGDBp7b
Xtk1r0I9+JGX03X+YYDApHw2F+Qt4082VxtO/iCeqgtWv8BAhX0A3/lBEkOu45YbOHQ1QBIQknAc
my0VEq6wW9F3kCCAD6BTJI6BopEJuuGre72T3+5sIsuye1TiToQJOlkUSN9YfGMe7Sck85KK1Y9P
BNQGgkALYhtdIgnNsC6WkhpaOnLxVIY8rl9IbYKAMXAKiohVi/DWL7BKajV4jGBLHm+sNJYFoil0
iLZC/RhTWZhm5nq0U0pzi4WURIGV4rpyYboqI8YcndWHW2ppnbh8jox7LdOpSv6oZ7UIV+gk5083
XXYLhCZKR0zkz8oUnYgBKKrE9Dg8fnMWujR4ntn8nbeOnzloYXwSnk/ftAm/xokVC0zdSojmT2VA
eLrXLL4JkfC/kKZ7/ErO3Dj9Q8FRjzJ5YB+ZLk5vhpmxcH1xCUrGjXH9w1BffupQoP4Y/sc9Ls+c
hVzXp/E9C/iKOwv40rXx+hh2X6fsV8zSBIb1psLMWJmWtt9lSz9N0Cck1I9l7QDEk8lmywfvmtCJ
vlw4fcbyiNE7wNnZ68DYTkuT3Jm88LCORbnAa6XqxuY0pKESsA2CVb/rg1DjU7NZkGUAPL9LaZeT
/KAlpihJpc0PMIu91NzLhX75P1TjePfcTgsMNIyignzlQ2WkgaT0GJwh1oso8E2tiXiI7s2CmM+6
tpO+8HiQ9MUmAgYV/mp8JWzTt8BwRSVm0/OvxPtV3NKTzEHU9nla6CWSUQiaBvT/MtSHacmHWMnz
JjL8NhfpJFIqeElKxlAFOgtj+VogHGDw6zmGWtAvBYw9L7dJXVDZzW4MRml6Eh1HKIRgiy4d4+gj
CtIpQhzocjR8bmcxBWH/f39CcJ+wGePYhDG5R2i8znQAmX7EedjAML1D8WkucnrH6W94waIxG30r
ZhrnS1m+mU7C9+5mE/CubrCZWlcuBB/z9cR7zJUr4V30H5HkssIGJx/xPCsn36qVuORqyMDUcjWT
HnXtkT69rgv0MQnpF3N7CQrQ6Kli6PL4gqc2l0jHXd5QerpS+6zDRjqN9nPKT4KLRlRXlZApNRhe
dAXnBAPmDMlLHnlgMx/wdebWh0n/u4lmBxOauheX6EfYvEpq+/4ILa2kfekJdKqMz21ADuJyv5rk
NV+1c5Bp5fPk7JvsCtkb7p0UYbq7shnB5r7EtyJUuKUZ0TSLfw79NJKXOnj4lXByifD2UX6DO074
e+HJv+90IbGvd2UF3tyJgG+F0+tZa0k9G8nZrbIQX/gHi/YcYEFXCJhZKGA6UBgPiumhukusVDGK
oLt+DNLaddSQ6qrHNumBp+RS2MbYwQcJO6Kj4OpiJNx9yF0hzUUkfqed1z9+AUtrfqdVM2ptkkiO
vaGPXPuHmn1t4XlxiMUxWiSNeIQYek+bUTE0aUcuWLS+Z0Varnoo2sIvfF26BdSLJJM07ihiybEC
yW7cliLdz04Dg/2aRhhZGeNEiYxvJ2SNJu1t7Fxjdv/c9DxjfleUegIDSe+BO0kPuwa2qVqRx2/D
4ad43g5KQelzDlfhQHcAT4ei9MOA9t5BXJvX/99EdZCTZt5nBv4ZJC6W+2HVK29mZ+Ap4YlXepwp
NLvIuDySyW5weHPz7mUBmk+xEdsYwWoAN+VKSfG4YmI4RC3Pk7NQL23VhW7O64evqs0YnmEcXyiI
LQPMP1XH1Quamy1Fv+XAuZeGLogq5EmuvSGEM02nd4hnOCu6IBAe0gU94ufEKNT4KjRQYscNSxp3
dspokNBrmwvrGk1gmM98o9mNNXo1QMnGXDDfQDH63KnF5S4JtjXVHA3U6UI2YERIWBNDTq3YHG7r
Zvw8+kYuWqZH7vV71lPZ/4YRVmVYLlg2gZ1IrJyMJz8pWwi2bCN2OKwmNtlodM4AHBn6lAdqJMM6
NBUnz1rLs997enQzQYno66I/g0BUmseE8nq5cOFIthuXCsAaALWd5HvTQykNHIESOVOTNjdf8QEo
0ioS9/+sB2AWZSmrwXL2OHRJvCiI1Ri6umKdxthvHLiEP57yZEcRrT+eaJ6qrZruikt43p+O8EHA
bbauR/zmhlgpG5ia7gKB5HzVQoau6UEoKQKZJ/WXAvStlMCFBW9zPlDnTxOIdiMdDRVgus8OQmYt
OE9V135DHYwcYJN8tzFo2Qp4KeGcMnMjcKtE7NacRO1dbUGhOvLMk1xoSo/UF7Y+hTUb07wWU16a
U3OYy8D1PagG2dLOl7HOyBD2vGz+dc/608Y8FQPpxgyCJx/mRhFrgBsyDnIBiT2lzbo62dnuSyi4
68ZyQjVx/zRpQr0bfGSZ8+8FFDvRdG2Yp/p4/9TCvQIuiB+VOuxdbDWQ7GJjlTbGzaS5rGrkd0p8
GF+6zLmkl08u1z4HjJuegxH1+OJbLbVk/IhVytl93HfPeTiL1Z/oFKXvTELEhimm5x9oXqL38Lbd
W08PSntgdeIQAlvG3m2GK1DTXSeux/LP/vrmIhQd1MJjr8Ka4WU776gSqftXHbUanvQkixnFFrEf
qOQ3zBoAusR0QlPkXEeWJO0LNEv0saTln4cJfl8flNhIivTC5LuI1XYa/+D4dDl4XgOM8OoGhL2C
4lcMDGfJYi8sNlxZbrdX+okEmqNHuxrp6BnZ/CPO/PKLGFfimEyPudLVbAzhzK2+aT0TZxhhRW8P
WjSP8KhLiZG0X2wMwjZmkpOOgXObaK6Z6oxplhqlgRdrIKUWIsl4I39d76c/OQ5BVvuGI28aNSuE
+gISYHHyc4NLbS1oWmi39br/SMKvkt05Ppm2QdbJ+GGN1+VIhwsIOhusE4CSAwZl3wib12g8eZ/4
pdNpKz11r9OahhKXXoH6fNvU8aypDRRr4sNhL02+zdEUlp2n8K227nU3t2ggsz/emR6JekR0wHEZ
GP66PTAzGjNKx5i0xHCCX4ak0LbXORtYNzG6XHsFobXxrmNmz749KdyRX93n6MGb5JQwnIbQ1AMT
FLT+negVuIQXzCf8fsDOb4U2ZUZrdik0efLYLs0IEVR82pexxdRbZ75nSd3X7u4v8bujnIXqgkqt
X6tOexrREoVKFToTXtye4UvEvUTefnkCKJ+2wG2yDHaM5rr4Qcppo0E4D+FrHCO8TOg9Rod/LIm2
nneHpLyalEtQzxdXeXJXkRknoQ1S6/Q+3GNbrUzUyUdcKUW7PTxUTUhYVfCZLiCHrWvmu7WjvTbG
oHhMIH3jhKtwomggDTniLmX1mPq3UPqT8F72KmS8jYi+jCV/zYPHOeX5l5JJElugeKxCUIZm4OW2
73IyYctUBiP22OtM0n0LaUynocOXJVlWLr/QXc3Fn1aADNT60yvt4Z1tLkCrTRcBaDI0U7/dNaal
l6C/uP2hXALB+GAB30qDKBYb97dYmDBFh/eGHct/mwA/ORrIEJGMeqKuv+45LFWnpgTFnEMH7PjR
S6IVcrGgZpf2bZiD+mUm9cjv9DN7J6HaAR68zZcg2zzpdH5SjVy3hKLIe8lQEuDELR2Fg3d8ntGO
lysFuaA2TlGFIiKApwo8YGE6suds2mQxJBGPaHYy9GDI5U/YnzKIX1juCnLSaFevxF21dj1cR/Rm
Fu6fwVN1l5WvNI2eep2hZ/vYcIRBfqLNM+mhAdnMxXEHTEJs41s9hNZMMkuR4bf9qsck78xIqqdo
uAYFJYA6Lfps6T3UAG+N6Pw/eDcoRrittFhcV3gePrgwPYLMaBBo6Vy8SY07ZuB70R30JAwr4153
JJpWFUtFGWku8Qv9x5tHqwEvMJSUisx/GAge5zmNCpIPTidn7cnHOcVnFRh5iigJfp56jKoe4i3w
vlKhhP0kKVYGiSffUQ2M7Q4rVrPRxRb4JrUrS6ttCcYu3qAA429sxMsPQ0FhgEDUZZL62KjKmz2d
ARunXkBPUiviMFpBoaKGPMyMKSteicvoZkt8uJ7GOOoJWE6NCHmCKgXaQ6G7o39a+JZSLhiGv6tE
GUpdhDWbQEAUOsTLG+nCW3eNqwdlUh1OPzQIEOCmc0k7VUuGGSwlyHhDQHHz3TiIn+gfXtzy9ksS
8G/WoU3WOPJ5L6PXuRK9xVgx3W1UKuzAuKxNMuGbA2Gl0jZ4HSh5i2ui1CN8W+sUnIVIAtrZiaRo
euveTNZpDj3yyhAJvtnq+cpbMFHjXAN1oP/jRn/NYNt/Q+quL10EHUpJJNrtCh8Hx+zjxl5OBBf2
EY66CpXK4QSsEHqPHHJN82OkvWnd7Kxi3wQoFiBXa15RgINdvxEuKbv4sjgYWJNiUssviyQ2N7iz
c1pwGh+90mAzF81VZ/4AdpqEv/DmNF6WIkjP2WryBG5zRleLIUz9cPQ3nPW4jtm1/c7v1sUiwlZT
wVutBNm2hk0b+UbMStfAaE/HsBhWgPzF/wim3bT8BIbQC9fkqn26VbsjhHCiqutPal6kylWyfdUy
axkzDUkdenQw20Yzy8mnzjE+VOhUekE3C78cFwA00nwFpbweLfqTSVtJRxWm6gZHg678SCmB4or5
jZqScljEaxYiKyOFFy/Mlb+9Z2Rb1TaNPzq8G/N2hAYZm3V3iF+VkCaCK4I15q3+Fh8tiGPJL0qL
HbCxCZCas9WRrMa7D68zb2w5UA0QEc5HJdQolhcdJ8AtU6L9F1WXYMTPqVLqt0I4MluJSKSvaDk8
Z48atklNHgVBTmu6oikA9B1YosezNr6MkaiV9b4mz3xA4QZEJWxxa57RaumuaKIqS076TNGZD3GC
BL+NKyKkMKoSpArRIhzP9NsUWzVnztqKtGEG5Ntt/Ng2iY6BaUOCuyRW3MNEmTNCp1cVB2AtCPKQ
SqS5z4ydKGpGY+DoQOJrCQyCsigXin6iBD3C71yiarJGyTtfsfFA1TM8t4PvkFMHCPAi8J046Q35
op7XLLEq14BlAgwLPi71s+zPJ6jkZrKxgA22Bwazf0j7rnfe6opP5AgmWIZXAcso4jOqcshmUagz
TFIFetII7HLIoYoAv/LCMZCIPZUPAPLyzG6+H8c/YfAq1zl2mY96SMg3iS/YyVTKNKMwmeYyHFep
sm6vRMeD3cpAnrVUZPlhGMNNuqNXslB3US5/Bb8Vy2Mx8TYIdT7G7zpPIrbfeFd2Xa4u5EP9m5xQ
gVQMlOcmmAPi303cWhMenWUjkSiePDrL+Pp1b37u60/76tTZVhRO7Y26Icz2Zw3LWzko9thBMsQX
MHR+kmkRlwMCUJtvcDSahuwPaKgGhv8Mk6gT5/yVsRGGgIy5m4cfAvK5euI3DyuoHlayw1Q93svE
d5b6Xs3DqILc+LlOCJEvvKTep3/giyajx0OMke9PATUW0DYZ3ueK/r0dZx+7p4C1U1u4Okk2dt8Z
GPXzRXHEUPsPe4yIqvhAzmtGY4+Xk3M0T+7xJiYJjUUgndmq5eB21HiAVl+ovQkWwWl6sUKm96H9
qlNdP5E+airt3vgIgrwdcJijbfmldl/rFVVSzJOSoLU6Wz/LN73P1X57vRHQ/ZLDsQb2x7abkNR0
b5YKETHf5fBu30pSw275w1ICrPC+8+VfeOGDeAYAyYRXmhAimbD2PSMezsf4hk9wIdeOV+BP1rhU
isQbW7qnFJGuZhjroenlx/8ZwsDqSFkv80kS+k/QJvi1YQ/prxNqk1Y/Imqm+Gsj4ULJRFnjFE3J
P3aQAHAXi7q9OMAZ3b2rMVJbYx5ZR24js6RpScnX02SjpZLkn3wYi4PQwC3RJVErMWmCKCNApi2d
BRfeLIJohoAoUe+cmcE1+//iqlZ0gSLH3u6pFA5m0fOHiWFtB1dkgGQcfdbYze/XQplQyYm8pQNz
ZzcmctmOpMEQSDVcOmDTlVs45wAC5cecC1PaXDBR5Dfvm0eyx0YPlv5q4pB5mSeyzQUwi+pcRbLJ
9RZjSCajFgbHOiLSDyG4qwcORu08SSNSP28oZ9bIgwvJ9FWLGINjOsSBSC9OfSUcKzkO4Vq5Bb4X
nSVuCSCUs/mP99kJ16bTgDWn8JySnyPqxfyuLebl0WOShCR0N+EPWJ66RVcIGGvy+cD3HGTKptKr
ma6/G22cJU+48PvTOKaMOTZzNBQUONqcfltDKMnI830C+9evoB7bXVAI1SctQGDU56FlL2SDROBi
wQPxgHg4XAoDPbQFFqodDI2wmIT2N6NoWqgZ/Yvs8qCCjg2uI/2JdCWGlLW99zt74DTn5BXtyeAm
O5ZcnIxLKWm03bqvvYNnHWlfHVFwYIs17nDc9xVcfq0KISpJfLGvZ6wDcyQexWEQTfyLPGqgPxoa
m3JMncTioOeX9nAiUG9my6xJPkpdZa9666hpSyPq/OSYnJ1h3PfSvsEMU/65Q9hUP4UYkxcuoZgS
97qQOr7oRnVUxzA7FgI09CCfBi6pp7WJG4imqXI7RBwOZYseYXkLC+UVbsCUWo//HVQEmyhYsa9e
1q3nt5GPQRra6jECMbnadfViEuzibNOrE38wFr0EJZLWrzKARgvaUxuC8KWbJO4QsMr06mZP7pPH
2LXs7BMSTqia5eClE+jjq6Rr4UBCzo3eUpYlWGhCzFcb7Kxo3OiN64m7ldqkaqYpHsN7mvGgcg81
h/s6r3lBEbDagV8Q9KxNHIWyOzzCD/qjMVsmEl7LfXxtdkCHvVWt7pQKCXIdiBbujESLyLITx68k
rWvd88HJmD2mBLwc3Fj0lduICYVCF5AU3OG1Rzy4hV33K8bXbFDXyILOztFAITs9msiSZ8zsNGol
7bun2x6KcDSzVFesweqNva0Lwjgh88GKMJeBepm3jDVrmpodmAc+srevZhFEUycCg8LXGJ53t1vm
jyfw1dBni4p0rCw7DhMq5o4p2ZoMidEXaVn3RgUGoEoq91fLRvd3wW6Kq4dopDlO2ibRxhNL1VQX
0ijNXtRH3QvBMlhz5YHEjraWVavS63ycel/M5qfPh30KQo6B0LRTm4R6tXOlrjlQcMf1Qu8M4RRP
N5lZskZlc1uUZSIxVrAoWSeAY/yFQulylEQ+JU758Oq1rEVFLiAMlj29lwH+ceXhHSqfZ0lGdedg
E0UhVDX3Pvi2DLa3taf88SB+3PmcPbTQL3xcRiXX7wxyBcBnVMsxSea6VLzTebAYt6DMQP6mG84h
L/J8z2yejpN3WvgLVCGD3r1Xtm96bVd+FrKcwwxCVhC42NiOWbjEPNQN//K15g4gYGEvs9UZZJNA
bRdsEWO7XFLBYV44ihEM386FVmvh8LbhXOLR2pTIUosGtfb3xoxR1W2allGLAxLsmZ4Q4LCjVuEz
wpe7/FqzN3z3HaGhy8QFney7Ij00up+oiwLXIo8K2pQQ3CmRNSxHgbE8SUkjqQysWAcERou6mvF/
1c2ov1hQuCEneQofYl9Ixh+9WdU/YzDLwqyZRcXFa7tJfIDMdd4AnTXRfgMH0oi8utRY+RQX9rik
Vx5bk9IiMsLVK8Lzv/QnnBzqQccP7Wf1a8Z56g19uyV1w9GpY7ury1DRV98NpszKFLXSBfe59Piy
Sj1qESI8mGzIvhAgs/dZ3GoR8Tdb37XDWxSzx/Nx3aRekF4gQk085lllxgDbKpgs/iihJn0WcEVR
fNjN83fWFKNErGr109wiUEtD25F2MfswHOksf+yZZbzbnqH2/M7mjLbjoWGnJRcyOl3HyQE+UigS
TMDn7skgP3Jyg3IAHIoJi7+yTltIKpvqdAgBP4M/DP7ApJOidzNUL3umYWPILAd42L8PVH10LoFI
8xIB5Z6TJp6wdZ/h5WnZ83Pj46vwbVbn4lU6Q3RIWbl7c66K1jQLW3CnP59+PzXdki9VMMdVpezS
CAC1O5+k+gq3uDuukD3UYt4ERY5603yQw6FPbVruLy5pPZNh6QY0T2J7pJFilwgoiGyXjkXx1Bnp
TgFjNBL38+RrFHb2gJApo5vPndkkYZihiqUhzBtaD3Uh9b4yrQiL+zy6hWmQPtPq9KY5Rra5FIkK
DSQhnWXcVkALsJ2vLQJEpvtwHbRCcbdQNdbEWXEXRVqrgm8SbDsQVJtl/GfLvCqmNLgMyqK6G9Dg
xz/xii+21izUci0JgZUGvpY9JWBVqvZRsjz7KjF1S5o+OrxUe3kC5jvni9n9BUWKKP7qvgReRyxr
JBoc9T3CN/fifWck/tgLhFVXKnAMAgYgiTnol0Uqd3EbvJyiJEO4NAn4We48qLYE37EDLmQu84tF
/EIFoLZHlB6kVRyViQLMVjG1lal2G5LZMJ0ibhq1ChYy1kRfHKRSvcEo3Acdu5daUqVUBAnp/IdJ
MSlMsLPWQ4zSH0p9RAX+G/vyV/ImGEJEccw/jGDPnhzN4RSZ51XRdFev/ynHYX4A+ZHpR7DxrCdU
wEvA67UFjpW2evV7YVNUx02uNwqxnrKrjGoIkeFbMjk2jkfYeQCO6GkFxALnybQJolYKMeOPazFa
bp3mIePNQZGgM6eqm0gLogL4anTawoH5OFXeezSJXE2X6maJncN2StkrkmbpnDQT8Pl91uJ7xzEE
UNnBIT9guSeEZxiv5BuSWyL3CQiyvHjEAGNTFpVZlmOQOxlP27rjMgh5kzT7ydcNw6RcBErV7xFo
ALWz4bLDw/MHA0PLyuS6liAZR9Pjp5axLUWbOjuUhU/q6XMFnL9mK2QIk6oGI4QjldnmB0MOamyj
KeCb/2G+uyZxs83fd4p44gOxMkjTpmmVFDYOPj404q/4bgY1MLgaOL14e+weNnNmXy2ttFvFthUn
hbBfO/8EDReJHgoC7xxjtLifa7QQTPzbVRzMxT7bJhoq706rZJxrAOIR5i450MOrVCO2sKv54Hci
MjLXoxkDAsJ97tGcjsskjpo2BI25WJxsS9xVUd+HUQ29A+SMhNhlI7juCpkrWbnJ6JtR0N4txA4J
b/vraPW9oqvizpNRlAVdZ/YsYIUZ4mXWidOgln/tYG44fjjIMcGiFXEopas6wjfdMWDJeaBuIvZp
OXUWe0Hp1kPW9cs3ivSqVaAMVHicWKQRUHnVDFHZq03ZbzHtKI/wbNMvIODrW5IwuSTmDtbTZA2J
pGmgmN2oGRqcl/av5sPt1bGvHPUfKFMJRWiVf6Cc2lEveelLTFirwtY3NGWnMtedDOe38UGShJ2K
jb1jTFT79cf30WcyQIg62t4gmSg5cle/zAS2+rL3BpT1t99Lu5ysUPw4YN9iD15uT9DQvxLKUWdk
YlPClgxVeZHzGoyrv7OuxDdMyzsTEzOpNecQj3N2zb1+UCEa1sNZlCKrCeb4oDI1K1WJj4g5wQrE
RRYojvHocZjtCl8GxbljufNj+Iaeb4Ymsg5XEAX9pIqtYJFXI/tSJH85YJmVL5VAAtH7gIIY+OWM
JznvGmvCxXYL/ezhRFaT8TuOyZSl4hO0I6OGTaPG03Zwg58/mPAiNOSmnYnouTcrjw18uuii3Bbv
iGof/mVQwrXpxzCcfdqmII0oV4GcEhOX3t+zylUk4AwVSncePC9Nvl2ABgto56NT/vWS5X2suUT8
DjXTNvnNLNo9HUmei+jdQClJ0OgdNeRVEWUC8uaceyXEG3ERHprrOx2fwNNotwbrvezRuVcrTqds
ogAN2tfrkSTYjxLvzTTFZCUKZsttVje3Y5mxl7uHHrltzyPYf4bnCm8fPqHENOwBBRjJluxvuOgu
AxHIq12sECEUa19kImzoPcc7UOqbzllcNxp8+YJhYfq1gV8FfhTkMxNA3I79smd74FDgjRv/+ZmD
nPB3EwLecprDLcTnVpOtVPokkDZxHASlwPa+bxqCtP85cy7Q1eeWZHLGMBxPBzIcIrs+jPYjsgO6
1n4BSFXsTOjBkEWs6Nw/xSw21fzoi+c5dhuGGUye75NKyTtlQ+/QohDEEk+Y6EnwiPDty9bN6EAo
8BvzU3A6BQisVBIYgyBe6LIBtiDD6omegW1rdgMDpFh8thdLJ3eW0v24RCYNSkczgqQcS7Nx8SgU
8ISSwLYcNtKUY06EnZTBgGDrrT8b+unkcBMlKPvh3NRmwVoFkoonsdwcIb7DWonbcIxZmlGOXe64
0CPzMR5+x0fnSen4N4SL/kiR23WQiC8SUvBNigy+bF3iXouEHpV38Z96FXIuHM07l6K/mmwvQykr
DTwDZhfAqhxfxVlM1veDSRJITPtJ+y7ZKpsGyWDVtApK4SFmUQ8Ws2LuxlFriXUFZ4dZ0TKj7CY6
gmBfZcia/J9RDTFM+YA1hfOyky4mmQBuPDeqTs6frPFCnVm0OY3jbxrYzhcXegjQfdc2APBlaqmY
F8sa4FFI87sKT1eKS0flRCHaziylwOZ8yVhW9hHR1ywOnb4mydHDdNXCu15M3lTSbFyxV8hWpEJD
LvkUvYNkc3sFU69z3JVLt7mO+FNIUBS0T8jaTdaDECI6kfk8X7j/1KqxAtx5n8ffJ7yekt2wJVUT
ptEzvKrSbdKIXSBpF0oVACsGJWm2aVOe7R/iVIvKgRcBoZ/0/jeKT2f2Za2R6HoNy847CB+OLTjA
A+b2c2rDmXABW3fzAV+VucxeH/y9/PNwAEByj++3PthHMaTrjArIVWsSLaPJ4KruWdvUVYKL07Hr
yZ3f2J+pTxnYDUMpeCruDl/XEQQDyn62iNGs/+LJ2efUpxYK25k9bA36fLCC7duXpGMIx6IZtfta
1fYHov6xPNkuEfP0CQF4yvmfiDxvU4GC0l4Wpeonf6vPd0SCuSjcOQtzNhTcJP6XuLcSYuq+/Q72
aUc8StKa1s0QqyDDtRNAhihR9KLiDMwaKrPFJ9+aJih1iWcIlwVzEWl7Guwt9Yib/lIexLmp/yVT
PPCyB8+qzD2j5yTTEYLBTAsMOYf1nh6loPmrbIV2L6ZkqdqaeXykt9+nZH1hkk6KoC0aILoR912Q
VJ+klgCCufXwDhXTSWNoctv5bRcS/yhkuekRUBh9acvICSEexR6YK5FSdUGQRK2E9YXng/kKvicx
0JLeSOxMefrpMBAaVHC1ZPgc4cwMhPmYP8Gfch0nGQgSd/GINzfU/zKbRcCzM2IJFnTF941wgwcP
4FqNemQl9mCikOJW524I7TdClDBiHrVtny9wnLBDddgVBtObnyEW0fObRcNMEPVxhIYk6Ed6mbjC
OGftlY4MvmI+yaTZk7mFc0SrSmcKMG/L4bT02Lk6AmJYUixGxUWklyJzHe7vTvqYNFNLySfG7A9B
M1E2vPrNhYpDoX2OToTYal5ZOXLMb/p89rJYEv1RWZ/4EFZWAuOHIci0lylzuFFtjAdfLYxXZh/e
55HLUpxnpd0Ok2EM8EKr66RUEBkU1bFDsK9jUtbN43dC7qbF/iGw75qvMgy8YPzJby50Upf+facN
NSz27Wev30Ag0FnqzGQt7PzUeeZthGJQj6CSd/nDzljk9aW4lZa2nVeiFI2ZB7F3D6+czdvygEqK
EteV7kG+byCRjSIbplTf0JsTYccDT5R0xh4CDNoCMXyesJUiJEqYyW+3pa0EzfTELK7F9KdMduDT
DgkaNrPwHPuWTV9/c7FvHDtIGjF7dNvHzIZ6AfpVPFEHmZEge4oLpaPbWNg9hozdVcVIuoTisnou
pngHJjHP12m5kc76RX61qLmo7Um3bM73Dhw3OtV0Ule3R9+Ytywon8qvsmAZi4xUscCE2o0XOo+l
YKW21K8fpRTbgb1L6hZvvbU3GYCcH57e/VshySfcdyE4g9Kk301Qi3wt6fMAfXB09hKSye5JQE8n
mLF/AcaIgZTJf1GTmumCy+qZopENBvsQuQZR5UIkgZKf2rzRO6lBX2L+wGlbG+8whA223GpRieo0
VV417yMWW8Jybd1zMz32mJLixqmymYZ1qLnnv9LuTR6A/qHFMnQ+SN+TXs5KRo9zmUSFA2Rr2U69
GWlvLqBviEitKflyuZympH0Is+jVmT1eoww8gdzttJ13Ua8nsz9zQddQmKXmckofUbkjXk8cA/gw
aUbsbWvFGegCND5bcH3cFHkSRnIDysJdvyDrbmLurMDkTofeYe8qEl6VxBwWuJuLKggKxh3t1Hfd
AV1vysUImm5GqPsdz15IRdv3PjPsOw7LFDayKidbHQqmniVWrcJlD3HitjNbYoqxJQ+gnu/1iESV
ZU5Sg5aGhJS4T4DwBptjatdSc+UTMlm7+BQFl3hix3bzJzVIEEnWp4qYsJXelCRcmXorzd9Ijd4x
JTnj3+RFlIfVq6W5kBT5/BK5dQuHiefffHhaEtHPf5AyICuQRSKuG92b5GsyicIHW3KvRexGuP4K
RSnVr4+q1m2ReBjHa29mc2XOagcyxn2wyM215fQ0OkG5WWhiDb9bcDToXUHO2R5/AAa3y/7F1Bf+
oFnEeBDLH0vtou0L1jXMvOrZeAO9fpz0IePTodeYaUoXmps6B1g0J35RbsB+aD5cdXdndvfDHVR1
nDVJDRPCmVhRDEtLJF5813aA9yz7IjXpmP9yNGZAQCd4EcknAs1c6/JV7a/3l4/os3tf6S+nAfAH
ZZWkTuuu+kmCjw4lOUF5/DtRwaH5XWeChD1qd+E1+uDtb0cdHRqJUtuhij+7hVTitQBmDHYGc2Pk
zoISiuAKUzulMl3K70z1TROunz8dxBlqFnt3Mv90V6k9J7risKxk5jgaQUXkg2jsyLGmCVjQXdqI
K0TXZDod9Sqk6QS6eIzJfJ6jfONCMMwP27DEdx2p2cqO3Jp/tZlmlczmtaNLpzwdTrHfrvz0InKQ
pM9BceQH5PyOytBviDYHg7vbwzQkUslQkN46rsnV5kU8qxqMo33wCRnjtOz61LOqd4VaP8iXaTDM
7v/l+mBigJIBHjV273CS1OhHjsiO0HSOx74+ltSNUaOoTa35KkBJk4uJ8JqrnHBwDdckS1yNDXkR
srilqGuqhfQjbCL7O1+t2vraFCDGPAFT57w9mOGDrO9nI3QMoI/4EBhDOrIEkTSxl08uaeC/Za+8
7P0zKScpVvBxFhBGJ4ElMsraOBjayfp3wMBQPVFe1w6gORdIFj2gLz1IIzUUAQ82DRL1auhiadOP
TrrHx76xfF35Kms8aYixLL+0xb/vAjFdAHqmMMWE5o5/TbHpsPuvTelEKr6iPlkf/5p3Jomg+C+u
+IFfm+eI8lu/wDt7Mm7d8q1sMhSSUiXDwFPwSfL9n0tGRgIRuu2mhkuBbdBET378VcMKkBZpZXs4
ngmieF//XMtp0Rq34YWUb2XmieiwXTlKzCAnGTfNuHnDFYRbkOf6sIvXwzFm5rK+xbsXiwVeNJ1i
430YPLyrWBgSJWnYcKHnexPF8gmPZSVSwJt4GqO7CcoQgMX1VTy4OWN3ybBJwrphsUP9lYioLcd4
5zAsmHUqvwCN8tx8lTasF62L87SDszS4u8sPTHMDcd4Yk6VB5J3swhYOFQfdBodNnqT8CqnzhU7N
zK+vR2UGKRlaWPXGn1fUyQPbrq/wYBNVt4H/NdlgGcYiwSY0VVG8YUnbpLguqLytL+7Wuv6aySd7
7/vxGaT5HvUrJ27KduEMmI8ykNcUzgKPv8IzRxvE2NgGovf3HJXsux+AX3sXMCirzXgXMqRcXUMF
fUfYf33l4MUXosxYNLqNm8og55F5syoinCv0wC+4YdYYw5AbWgDnUQlLeOZk26asiZiBr6sMVC+8
fM9+6q5tZ9Q65z9XsoEINUxmugCxxV17TzjePcsXw7J7ZeTRdpiPbN/bmk1ln0v7gHM9fRa2u3bE
5MPorBSLaAWINzkxUkboZgBCkbEaEQnYjxRsF994JnbxcBxauG5qPLV45rPH/ItM720YfJrr6ZE3
dNamGzmxwE2tKcwHox3kbdwZw3iqMGAKwfbbymuQIExLltLaiEw1vy4mXjDgrFNGU+0F6i6g/+Zx
detnBmrDRBwNRyNi73xCyU90vOF9XImgV2GrtwxSFrCZ/R4dtuUfNXezkna1tohUup7Zp46emrP1
3ok5/LZoy4pxm3kHp8K8Z/O+HTdn3IsNdWuC9jAXhn3eGfW+6aBoaU7SOkdY5ucfnM5x7BYblF8l
HpnN8bUcCH1wyhq6Vh8lAUa9rqNlUAgqhu9LHfwkJBkF10VxYKn6gAkHLDvsXMkRydNrLXQ+yiu0
cgU1gTcDeCAAWBX7LiJ8ovWo+6whRxfKOr0wPYUP4va35V+OZOS/sDU2553+qhjvHMZR1fwYs1IA
5nAbPnZY7s5koP2lHLaQm+Lt/EENg2nTvozMEEKMi3SsVhHmmf5qZO+oE9gY3WUmHr3ArLrCy08/
ALQLSvkI5WkdMI+WaUvl0b9bTiVxWEjQKUcI1Mvm6HDge+M4gF7ZMQUqf+19mbAXo1ofa6wyX+05
aDOeksO8h09dK3OJkUgh+G6R9yuQIFCoOut3TKbJ/a060cd+ksUHH894h36lehFqw1CDkWUNEWyW
4aXp4MY8/JSB+NDrN/Tl/5TS1KsN/zbXAmmdELLvFV1ip128RUa0PPfr/rR47anWGRwR+WitgfJI
fFMd877uvirH+/pugwhmW8aPDYlFdngFVBFBrhU6QWO5Nsm5a5b4rJK9672OqPRFHm/3yZMTcg5x
31nP2OFLsqbEO0HP4D/oBgG6YIOznMubJTV0dJ5Qd13STuH/pR2jcjOOxMIGJVOgZo7UlOkl11jH
AcnoaLjhZqK0/Z2l9ybeXbnFe4qAEdKZE9elyHuWQp0LTHUk9i36C38PeONxguU4/pcLFtRjYmzI
QoPkAiXCXPRqu3DNxkBRSY2lZSRwFwgAc404cF1eW8YfWttqlTPhru69ANuz7UdEBwni7U7Um5C3
lUUInPL0qftsT+BBXvLT354eBixRYfLFVtdq/osCBTS9DbybaHqWqHkZuu/2uaR9mskRa8Dck2ba
3DeQAOgLRAPc+gLRI2FTV7uvMZj4W8kTNqJw+9qG9mklKxOer+jxI5+fX+fikvZA48XWlhCij/5q
T+nHo4shhdrG1IUIJ1x8oWgdL/wr/xHzEEOEqq8LnIEdioRV0XZO2pyCbBXW3tnZRo7kE7kR8sVu
i6UowZ9YDq9ZdKFTRs42O4Ljsmr6ZXPZqM6eN5qH2281IuwOrRAU6hHC91KVZUEd6gvvL7U9E8Va
Gb97nuWklISR6LVhdFWsfVceMkcOcWk3AKwYLAYul8LwqhKEy1OP8f9CR0iMQQywHjE1B6/d9bNt
DxpG+xxK7Lb3iWAkdRjMsJ9N3jWbsCF2kJ+lHCcWk2Ol4RFWcBv1zrDcp28FC1bzzSGQkFe7qjpc
fb33SBkWqd5Zw3UB+Up51EuT+QGJDhYgQTTGBSB4KmUQgWQK9+axaP2Mv1PRVVOedTukhoV9XpI/
Tj0drPNh/CaLqQyvDxCprrg+GpfHIAkU1LNFLrxhXBHhonEu7EpLOxx981W6pKfqsg3+IO33CbVU
Lpy2lf20wxkeRgx/d4vD/Men+lDhroJ5M2Ea2lZwKCnlN8AcrLXTNm9l2CfFaUYSVvY3T/E0LZ2W
6ZzXWgQqE+JmEQ7qNcqjkkfp+N5NSl4ZSFuEB3GFAPGYGCzQ6mzdr/VtnX+TUQLDftZaC5sJ6qBy
Mc2+Y4NCyXKec6i10lBAYZLl1OSe/1Ann/0zO7QCxzF/mlqwYpCI7cDkTtvx1E1AYBtMwPJ7QDA/
kQzU3R+kjOliSc6khUETspJP2jGaVAfGqzhHA/gJIqkJhd7YhMRYtJZf/wNet2xDVBffQJQDHm44
Z238xwVgErvqN+xV/xWNb1Nvi3+eHcV+BaPORd0egdW9j2LDlNG4HLRo/PecdsVkulyrnTHO2P3f
Y69PzxGmIYw12jCCjYlWHUz93BOCo/KaZyLATlqcDl5GADKYiy80K9OYcTUnUSoaUJ8Zk7gVIvgH
LmjSVSh27HKTreWTmk/NjNGFn9wryvSwXA16PadAyypTYPH8rwOuQy8Oxn/p/FT9hXAgLPHK6SSX
dyc0VzEAUQZaO7PEnL2th6noFC2mHVZ6W+yKyEcKIX7zfHXeIrSHmYEg+040IVekfLODzy/HliK7
8nFqJu6Fe4voFBI9HPOtz3Ow+6MBXMxYpuV8Rl/wKL4nCe9ojKdRpQpeCehkWfbv3xsSeELpRdcz
OBSY9nE0b6lKYFHlPT5jM4/jKO7twYB3SR4Z1q1Pw25angHQB5G0zOswisgufujZPbMfJ2FH4/gK
UvYtEPeXBB4HHPSA2llsPJMTO/X79+S9QVdy1t0v1PUJ2KbEK1xdB01ox23usHyjjPfA4nv4dkmD
aM2DDfWju2gI235W9lqsqj5lN/bjrsU1MI72JtsjcgCNKWjskReQPiMSOzzDQjzlLPVIwBKcUa89
zi1vXgzvOrJm0vpGfOyZvL8vaDoU4eIs4B4Q9mYed/RR26WJsfuzWcxQqxSNuyQ2J7oQmex8VhRr
5nhvzg9mm3+34SPuEUyqKsNM49HHMKik9M23J9pW9YWVRlqyidGm3LRRiEdvaAomNPWtDl/a1CxH
nuFI60EVeIE02zXnokKdRXteR0tm78dm5ZBHiMha/nOmOGdCqIZbEiOC4qx6/mYswXQoobvCyh95
eO1VWTumaPjxgiSzTg0dt6EEVTAwEyJfqxav6hPWkauik4ZncLyT/v9hUunpVRk5HuZCKITUq5wc
bz+nyDoBBxvDqwTe08Ktl1m/7Wxgkc0x2ecXxXe7rM8q1e4dpiJ6IpzeqaEVh2XFmf3yeFs+G0vD
jhF2HpUtvpIXXltQNsvOySp6a79WomZWBn+1NvAt7+JpQ59hsXsP9C1CtD8CqvZ9IqJxwpzWv/0M
ZAbE40GYEU1PtgE7GlJXDa/GvixSNwvqNjKkoOYRp7lIgrxfVNoO40KQ4SCOBWlzJyMn3n8dXbeI
ZYFMZAUoOc3ke6wNK7h8Q5GlEwizXUTQoCUt4AusSFkLN6R7uyfw0oMsx98I+9QwsfeXoQHyL/kE
XjQvgtya6AAQXdhqsMDHc2V1ECYSCcx8Ehs/Hn7FRx2bw5mFUGXI8itHrzN18hDhCn+YiZLer6QH
YBxh7MuvP+TGoCmuaWtnkR8Q4HbYQcjTULy6h2SiTH+/1MxYOTouNxFcrrKYGDo07un5VQaXpkPt
46nhR4w3RcxIOVIOyCRmQSW3k2O3ME0G7e4eyjE3hXU6Bw6L8c7qicl+chb2HoFnLig95kZ5919v
6pwfY4vZ8x2uD4UK828cHz/qzblpNhfpignzLwy5ULeIftZDVl4w5kOdgjohZq4QwlkZmW2oZnHT
d/KmAjtV5z5qcfyYrL6dgtlLWM9dxdIoHJJhnd8iiiScMn8k/cX9wT5FFaogx01lv90EbDhfOlYw
EDouKB2ptDslRDr6fESpMnOYx4UkpmaOULsMCUeSOS83rHlv6Awm7RSBUZsEjLTRRgVRmSV8tWP5
1Ksb8RNsxbg96NIjFx0cXdsL3dGih3+LHzaVOoDZe2vYEwzMWsN31UXezuw6Xjy53wyN470GtTK2
mD6FPeA0j0cQ9zFT1PKgAGzBChXP5ZLTsyZ/jklkMW4WphmNFK+BI5hSbjplee3WXsCtWxDCnsrB
fQrDMg6450cBa3FJIz3xukDPSNHTNro+Ew8UO2in9YVGp963osuLWkfmlTDBrl2IFh59tyZ5y0JM
zq03lXedVhGwGftGpmUzMv0R5b8USODvGcgRY+cAbLusHi/EUtgMpN4oN9tdRn9TaERjML7M2n2/
++FgNV2oYSqWh5QGIxEeqqdq9Av3gE2ih9FopSD4XjAFaVzLQqJjSzhWQ3K8pqfrQIY7GIrbo2+v
BFwD+ODo0QF2vrNFZhVFNWRlP6zF/3n7pfeK8lRWZb8tK7AISLqkzpzyxPm8rmOzHfPdXrbpoVWF
ytF8cGOmacxa6zxnjxSh0L2kPAHZys7jUhyIIiaujSPgWhxKTUG+Pnu3eDY1mBHKUPwa6ysvQipk
7aOQR32WIa8lIc4jtnwQFvF9AtWVDvTmscAhpb0SLA6XDzGUQxOXokY3xCPMq4x2ismOGbWMirJj
36B4rl9ReAK/2TE5OVmfpViWPjW1VCeOfhLbTEYZTmVEfAMQHAQ9JS5letqAwtBKrY+IAF3epRVy
5XoQwOL//NcZ1be1ezdeeYPsgQhkToXxKmy+fiVRf+YNPHWZXYa2IUaWxrKOP7We1CUKmVUeBD7n
48wV1fhQQ5CH8TV7Ji9j7JzTRgBuf/kxM+k+ATFKmwCh6u8BJ+16Ec2LrXvduxRudgHBrC90NGcP
mfmvR4mMm0JwzTt9ZnsFtFlm081Rf/h0+zQDNkBwAbTVT8yTdGyhhLhIRZYj5niC8y3m3sYox5/R
TmcIFH1fGeQ0o3I15HX4CP+P1ZYUtdehhj0mCUq8VnXnRxk/1lvasPTxlI2H3cXFpKr10HhbpQsp
RiO8bsBBMQipGG2DrbdkXJmu3sDULy5RSvRbisCOt4d8eXoK0B6k1a7J4+aVZ/hr20iyILK8yEqI
d2LMHpZ1Kpu2oBeVJJwwqjxbnwZmkMHfvhNZO3gXKFizZn4+tUPA2iaIkDX7l8YglY+QTTtwPNgm
OiaaCxETa6S9Q+8SEnH+wZz/K5Tx5XmRPkOq5JWw8tRJ7MFCepsQYz+SyLXAr3pbdSAn0qjx2aGU
uZ73xFWo00IZgDjIDzSipRuPz0OzfVTMwK2QlWJI5ATRAUE23CMUOWnxZR77nvJZrvBf0OzoviUm
OpjP/7oslPDHGJK3s0AzU1Cf85I3mlR1j2HfjqtAMLQFNPqVzK6n2CV7/gDnQp98+D8HvmtnueMC
vC/7NbBM+76OuRsIwhIx17wPFNPpu5Ads88LAWMSdqzadlaCojzgyy67bHC3tbYjMRICnABUerlm
kzJpFcbfry2AC8NGmwAp+UIYGz92c9cpY4SmjaF2TLLCL4Gh8k4c74MyjRWAwg8QbJAWoc5OVcaC
e79f54v4m4e43f/xTd4qy5xxDnbcGum9+xzoMyuqs7C7yVBCdjwe1zf/GbgWKI6n/s1A+y/Xac8H
NyQi3wB2wUMXj7Nk3s7Kdi4uK3BYYdVuiS3vHM08X+hpKbuKQ4JF4bJ3ntZVTL6rzeIDyyEHwhuu
p3hqhl4DAAY0WwNDYbds76V2BL8uECJ693Faez8kn/uDji9DA6M/r+rLsJrW6fpQA7YWzyevYt1q
Mpi6JRbEVRZ/OuI69Kgct71Iy5HzbPbcFJh3UeHj3FGEVM+sQC6fXIYQ2fjjeLG412MrykwVbiT6
4T7rGXB4bu7PIur64OWKahV89XFpjxVq5PPkIFM8vrPJBP7T6D8GQE+RY8xZxs0t+Xf9jusB7qH5
ZB5ObopmjywXSlsDtkx7f4d8VIrG1rKTcJXXRQBAdj0oYdjfVFkqXlWNo7Mu2hHqA0Y5EDIIXViG
8uqR4pQVKtOtqeNm4TK3yBPc4EUvQcgTELB7YVH8Xe79sQYaPEhn2pvitf8i+fWl9MtfNZWYZned
A/j65l6MQMAeLP//SNswucJB/U4RUQ0x/uU9TgYvrNFB5SRdz0cmLH63fxb2HYNCQuoLoz2Ih0al
odY7pX4DCA/ZFYKcuzTL6e70hcLppUUznZqvhtAPlGXfg6QhNEHsw+Q2U2vv9nKMtb8VF/OOrEnb
PgSu+nGZ5tWMNg3tFXlp+PjMVSrBDFb38/s8kk7H2xHS6KOJ5/4R5RnDfUL+TUyL4UyozKhpFnkJ
803zd0sOy0oaeeCDuz0o+tS6MNZwiiXt9QxxzU3Y08rdlslL0FYjYI2OPDI9/kYXl6BN77cn9/sd
s7ofzbnYhubUyfxO3GP/FKNbEoGryG1zgiCATSpualCvR13Sqjm8ifdvEt+QydZreIHPqefH8mfN
caed9u/ID8L6yVLxY76L0yE0ZdIgpWVpA6k+jC4qELFkJdJUbjoaQvjPFNYqumtj8ZH/+bsIOqSA
/K4cXjnTcAYGBzHbggipTOWPiV49WSXIwVfOTUOM2uCH3kSldFIP9N++yr5dYE+WH5Hihac1wg8F
+UMgm4hTcJTDs/NpixPLkvUBtvSw9Q2iJC+PCZucFH8DvzQR3kZsZm5p10Q5bh2p20nb2VBTaSGK
Zgf83RkveesF800KiliCVIkfXUACosdtm9+ylj9Z/Y0DKvbLE51Zl/A3Z3lpVb4bV8qGMvaszoxx
1uKWFTlMOhPIFcn2ROR5QmiudvpjK9OMDQIcPmt5Y1eJZZFh2neOe58lUuqmG+Y57YrJ4/4Ch7LX
r9OxiAJCSMcZnXrbPNodMGLz/ZVCUoHIpMUdlBZullQ2gR+kdLD29R1E0GFOM6luZY47ch11LUZt
vlYDwazQadS58JmYcs5LMDaMMeO9SZSb7qNjvHDJtj26xPtd1hvzuncEEV+J7ikH1sXd6rPBNvq7
2gCf0PgKEe/3ekjNSHkSd7DuXiQufZJ1jOsW2hpR9SCnZNoZ2aUE4Cv5DAqAg782iidx4i0Cmfne
kJ7Pfexe84M7+0PP4B/mpjwzwFHNgI9mJKEgsIr8sxK3phRMPcaBFMcyQMVWvYvZ+9CPIkDpJOkq
AmmrWn36kNc66XZRaEx+3kcppKLPqai66AxTwdLnk6g4GPouQ22pK/vD/P2OI3MfgcNUvmRi8Bri
/6waHG243tZggDYxE6poIpuNC/a8CPSRnxOXmlDdI8HYqQlqGSpd5V3E5LVU2zm2avCar0D5zJjf
/6zHziAG/4QJ8HKHQGSn6tGxpHQP9Fa9OHiznSRlUSKsXQIUNq5pUNhLcYVuc+JoHsIIjgkr0VxT
yPPJRab+Z1vdWfkOBYWc2qE4xPiHctjNle5MuzAvgAJXJX41vTsXVMcsLBxPhEiol2dGHomRfIZS
mslPbpEX36XofOxhpByiqOT9rggS5qHGDsCXcKK2nHAkAoxh6zkXXxB+xNZYVVxDbxR84H9awxMA
X0yPDiRsjXvmlG1aTFHwaPWx/LUcEhCnsUXP5z0Rng50ECDUR44m5Lm2mSPA7T6+nVpV6Gi/wyb6
hG6moDh4x0YkjBKg9yHGt8NYVyyUzB7RLIqc8z2qTUcwJPVP4lnuZfHG7xBsiD+YI73Nx3dokf3k
H/zcOQEZ7Hp3/PMTTJ2QEJEqoLT100UtyaI4bL4JijqZSb0sIzd3S009zfPkiXfIjwv0vsjrGfhx
vayLPZoEz+LPPJmgh+v7hga/Oq0E38qz1KQrLepbJ5SdMnEc950dS8XLytajBKyORjrhdaI3pzcz
9vnxEXJsLPkyqsN4sCeNJ/pD1SF10isUQmSkOKisLT9zZrzhRtku9WwGuBg/niR4tUO6ABKZ4OV7
hIe00X36xpv8jhfvgQqSKckYA9ULklXVLDXeHpGlHxKMa91dog6f6iXu2+gkwHOKx8QpYbEacm0x
KMYJ9sn3Dm86JTIMrZtRuYkrAxRZxjPPrY0SDH4/kLtzy7U9+vcTDJlysHyZWO3RxTbUiC28G+nT
AJtk23zbRUmi0OtDrz6i84LQMMDO9bcTiP+jEjxL0NAGjGxX2OSrr5YFNZwqFdmlLeWFS4ChecLI
9cq7eF05ZRDuumjtY/sDlJ64xNzmADdy5nxqm4o3IUQs3BAhHSBQTFeQ9+OPUZOhBKjGYbwK8XtS
8v05+qNlfArc9wajs68BCn0zdZ9SlzP6skxsdgaUJ+Ritoxuz+BDdZqPlUMvvp//91MpjbaIanet
6VEgKUhTN4hDUlDxbvmTffWvDPKCwlRll6d5Lf2jS1D7SnadIOSQvLS6w+YYbzX8u/eC+VmgV3Ia
VDPvKkrmroWfXxtGz33zEZoZZh+O2BZKgOYFRE/N1nWecBWtPUZM6yeTzuVR8Uda2OeIPRtgieto
ufuqAqRrsi/zAXI4y7B8KUx7VyGQlqagmFt+Dvpe5F8Z87IHO59ajmrIM1qwSk65s7jHGOwZFPBQ
vKjuNIPy6anRH+rWzOKoGmgFTQOyalu3M3JsJaGVv708QE+2muH8MLDUn9slJZw1cQNL8NvPhtWz
2Hwmto+90lCOjuVeYd0oiDuTz9vTXFYpJ4lQL6lPyvhrgE7y5cxybnQ+xrXRTW+OFjwyFt1/SrIL
BfaQFz88yOcr2dzBi0BVsn7cwPPhrI4NkONgsRygdRUsBWIQk2opWi0OgHNjJ38sah2/3smDUNv4
QkkWD6tU7NmKCv6J9yVAYkKxpGdX3imlvEMAEyJYJjoV203vBR4HE9GDV1sjia3/uGG9fSlyhMyp
1PjPTUd1u9+pSIuUpDJfiQsPYeLNTGD5Gjf8rLo/AsdfKwUCSewCjpv2ndRDNHIogjJSwEfRaa9U
W9WAP6lYdQCc+/V9FrubnTFY1kKCpiU+gvRsBw9QImGQ+QnA87MzqqYov6ZIuKKaLgK0dt8gc6yS
DJOtMLXlRKeZeag+wFlQ55qjOnx1lH8TTPDbAosYiBfUiSvmVgBdv616OhkmH4fJJ8ZKWkBjCoe6
+PeUxN9mo4yIW/52D1Bm2riuggPVM9rnuh6qu2RJcyoWIrBQGjckSjLSZyBjR/j/kcXjtx7g5mAc
8YlVLKnaalxabOEZu6vw17a2Zfs77sL06IS47xckdn15pVn8S2HmqCpzgS5ML4vCkHNvaN6BaSdg
RnnWDaHd6uxgIkCi4KTgmlfoB5du288lU79um5+Qrfc8NjAlq9unwP5ElMl+vUd93OBqLWk3zL+/
GfaZi0x9SYpBTaDQ2RQLkRJui+bk//r/JVnVaBFbLMpvxxeuJRyx9N4hJMEYtoIjyEcSXdZmob70
Km2V8NFo4zPry6XjLXB3AfpM5Jb0+Y7+v55D9p61ZtJBhCzro0voQNfj4Yh7Y9Aba3dkZjIeFO0n
Dz4xjOGkxscO11oIXKnZamMdFRoy279Roqi4tbtWVClaTYHn35NpuZQhfhh7mACfA44tdQneO8JF
FDubLVXa10E0VhJgXoIwMigMTyy/RdwonVht20SHU54AlJPg2OHcQ91KZPyo0XHotJsVs3QULtUD
ecEfF4im5cq8+28aC2GImILiEFDLBxQhYWgsJ56j0hqrPnli4jI7cH7ASLCWbmLHqtNBmhqLRcCA
8V+41cHymEO5ka8l9khlJgyOF0njIFNjvIm4X6p4QKpA+6W4TRAlugqA8hCfr3N6Xi0DPI40rE4P
1FaFswumLOHSEvZrv/gEqJjwIppzeQyoJ3EsoT7s0xgO5uf7rwXJVg4TQNb03gtTO7iHyp0YpwII
6mtQHZUuVKtSAHKYz5k8rFDydlHrTq+W5uXnDj5Q0fITN2Flb8RwkMhmGXcL6r9jGBZysvagXfxt
xTeqc4uyk9qhgyHOgJ5VowS8LAHSGGik64mf/Lv2LbbKA5pZ6ggG2tXJHhvi32T2AFKcouolasos
KcGtlLgBVo6dVoXLelxfHuPm9sFXMQ+jm2GABgQrdeyco9H2Hs/F24uKeEaTaGioYItckRcbOdVR
G/s7LK3O9QH0s5FcIdf9w9Syt4+3XmqXSZ3QdrHHs7fTxntMju9B+VS6cNSZpo0VTNZ8jmFsujoH
sQdlm1prvGPewWYEbMnsVQ2/pwGs19fvRYUG8EvgFjS82zz4wiso8zDe7uWgUVc97n8diUCjrwYj
iHS5U24fTlzwiG2vFcMUY6HhV8Fg4NnvHstYWoEmWYfm1ZHEO3B3MpwJkK1jSxm2ZZ5G0Zv09PbL
6NBnvtClYAg0E+PUekgBQic2R7W/UL/K5sTzm+TUChAN9h74WCnW81qCJn3Xj6kvrHoWuC6Rofo4
tuqMvuqcG0HAM4B82xYmoaBbX90Amowo7wn3XoFT9wnbo/SZgy6TM5WZYhkqNM1RFW1YHyhos17/
egOf8owVp2gdRrW2zkAEe6w0d+lh1V4ycvWV7L8izeqRWkc0LPKmHlokvXpEjr+2pL0PZrvb7put
TKk8NXO0DMg7sBxj5vcQYdT96ibSMpdYiRx2nyStdcxwBz8udtfwO+benBhaIJQNydPILPTNk8IR
PC0oHwn9ydo8szBcblpMlDQCRCfHrWxN3rf9fAnbkZqSVakvSnNnTNEKYXCxTxUBkaa4P1EYu+Iv
Q2E7n/iiwPpDBBcLmYpD/RcQYajpD5zFynsnFmWnaY96Kyip6Nh4nB/llBBTtC6tJdl2EZUY+W/B
VYtuftUN6t9lcrO2JlqxM8fGhOAGuCCFSZrhfuG2qImnUTGVeueyl51zOGX9dJBN+Gsl4haXp5D5
WQNI4ibZ6FpeoS/kyIMHLpnunk53HrkP9VhcQoL6LZ/ZfMaQPvqp0WmqMz2fsmTIVRjy/XcqnGDU
56vbe6e0EpWWZSHbaWJSA1Fa6Xfex0k3hMYfSxd20+KXlewEpFREkhCY9A4zafhE9TelXXDIvnU3
o66uhkCBvTDy/QsSUOOuBvX2BimNsI8mjOE7gqm0f3bZbW+767dohv8uC91syXdYi7Mfa1AsSixL
+YmynLPsngjUFcKD4le4X1NvAb2dmLfK8EmUNwLxIAO/Tit3/KeQfABEFJjYBf+k/vgh8gxeRXJa
M4XeVypnsxlThTuN42pmVDUyXaaE5+1KRdEp65Ceq6gbFRLljozEanefBEdgk4rOOiFizNGZKOJ5
tAZZXVgVF5avKj7+f3GrVsq9X5zZ4dz4Ev5cfj4lw6wHzj0Vj/8/5tmiF+J2qF9PGxnslz+aK4dV
xYY0meHHOTehNazV0oZ3YHxl1HJ36migRFAuB2PsNxwSNa7vuNqKm0jg1+8eYmBM313elS4m8vDC
fSRkRj/4uOJq5p95vxHDmxq1IbZfoE7NntmOeNNxNB0y9yU15kIskZ4CZehIUhkPcDM/w7nUSJ6f
8u889ApDdV3QzJmkkyMgadVV30+YtgdIVAE5MuVtG7sc1tQ/vjFfnZdfu6KJ8jGlvCZ+W0VeMxac
kTLDIhRyBb1Lcf05rgOWTchoO1cxsfga7MWjtdHLFfz8o5QSbLSnebG2zQ8mNfN+Hq55q2Ig4IUV
6gHK0LfkFonTkGUWL3Z1SXab7IHOHGM+LScG5anMQlUCdHsVwex9wGyrbH/yrjV2fqUvJ7j5LKwa
fdaBk8gzi2GNa/m+EaMsCvx/q19xAOd4u/DRxIXFyIol/yTY8v8MjwAkcQYJ4zRFr4/NpcVZ+Ny2
5CruZ4EvVOG+h+VpW2Fomr0f0mXnViSLmyzaHvAX0cNlIg/lbZQbxRZUSejU4qt3VQwcw/ABGfdU
AFS0X5aAJ3RM+WENWk/i2eThSCt8pP/oq2cbebaiHTjC6M79FOqJmW970a1osTxoev1XRJVXHHw4
tFF9cibEnK+t8fstkRWk8yqijsfmFKgzpxLDOENAWwZ3ewUzAmgXOxF8P4+3fImhZ7I6OakeK0MV
iPUEbX2C/qbvzipG4zTE4plMfeOceLrjh3DsK+Dx3fTm36b7/4MvXboKaDWW6IwZsOJ2Sj+RQ3mD
lqhGqNkMxHcJranqH25/8S54Gh/7+J1iINlnULagSbGcw3uATJnkaMZI06ncwS5/EyOwAuLaykdK
Z9LprokeGlMIxwroo1bTklH3YUVPReHqkj7J7FkqTz3g3KI3hmkIqoLvMwZdDXzR5E163Az4H7bH
Thj2jS4PbQ8ZirRdNGQ+4i3bhx/n0ELvcW0SB0F2lAa3xkUJ411oMWjRh6r8IqQIAqzGO9qN5fU2
XuOVbXfBi7weADhlB0+v292VeU0eFBVzvZgSYV40/35QN7IYDCJBX40MVWQ3EnnEk/kW3bEs7zo2
ExFJis70b6QZn5FXUimMPg4+mWaKS57TNzyNvXuadQ1BCobD5DjmTRREvGhrDcVP8HHaNWr7pMBR
wpdd/dR+h6UveZfAH6Zx8f1jd+XOswOjySF2PBPucsWZOA719ukRIopTvv7edQWTnRF7RfohaEcW
QpQp2IaocQ2p/HTduktI9miOg+i6xT5MQLT9N9/QHCWQsrVH5TAiUfZvi/VcWtEuGLmuyNB98JX4
FTe/oklaHtF6FD1zlwDfHJt908diIWSyogtJA+b9n4zuDjV79oImAN35FVHfO9z0CbesWlz+6S9h
BmLNyrFIkhuo2wZHAWTDr5jm+vF6JlprkHkeb6xLvEa6ru0+VRVJjCRVC4TTuy1n8C4Wy3QYhot3
nK1gJk5yCIt1uivwENYk0jTg0AxAhLG0fLe8OXPhRkxV025xRTwsBJtvYJuHt9OTDA2l3kclMVSL
Tj/A2HgTyMC3CiVyv8v2CCbjVefvsCnHaghn2alIuuXlwyTYDYXOF0M17JsOzxu1o9idFkzzQFjh
gKBDc5ZtOlqYmF8mhWW/0JOysYcYUEBmK92feRcDkmNgIMly6t/87DewXCaAHPDsRKeCScoCEBSx
GD/4fdTeS6yIDsCoq8Pe9yM+KHT3Gq0Nmtje0oXbsvbdk1ZbpOoqbXL8uBtVfW2VTXw9HVt3BAy0
GFBHXwQ+DISWaRH+B3rJ+qc1izoKLyJ5N4B1mDntpIQtxtj490G3I9Yu540aae1cX25Ro+MdPR+U
DFUUuG8x6ngKVn9sgnYmLn2TndesLAtJXFzHILRdCZqSK+6i9gaRZCjJMAZmUS3YqMqxiZIhnsPq
u2TbuFn4mwMXqls5fA0acdRZpf2GKOaBByQbTQbi/coZHVUh+VRLgy+QgsgFG1ef2bgTPYhIO6tY
oXqf9c/JQc4iHs2KEayFvduXvGk651vs1sttWIxfxvXBjTxpK4CUuleflBABOPLYrtpAHPBNWGAN
3RO+5MdwU3NRzV+rpGDLnYg6LIbR7zMmrrsI2QsCP8ayB9VvRVtgLOseTA0nP7/5CUgmJXWSKOij
pYr7t5Dvps9G31/L6Ux9cETSNQZ3xe7sFwZN/CDVZGhKg/lut3aTVrJN4HC0Igm8omsmc2YhX4V2
AWLpPaR79F+SBUDnyX5ufdpJkFu6tNrY6iSk/LG7oAVKW9SLjMi8mdEFW7iHOGl8CAxoxcvgXzTv
GV7a8EXlw30J4DWvYII9cTQneFaETkh+n6laQKzANm0LbUJ4+E/98H5xY0GiiBMcJIUPPLhdWE55
dX3Mup2QFZyqAEBxM3pC6LK/AjUcn0I/qqm5UtQslAmpcGMvOFJ7mUiqBdLCnFyPQQVte7o1YuVZ
kbebefyGikMrnWPyxDK+kfaLyD8UKjcB8MBMJIsHwlWLQCEMuNKhEU5zu5wnjquzcBhDAKrlxoBj
UFiTP0nPqhcAcNhbJTwL25BvXzc3/6qJdgzBH3DCxIWOqdw5f1AF5A53FTNpYNTKAbCCaCyAYnzS
AXc6UbQqTdnj5SPryIRZ/zuH+r6qTMD9V3qyPfS96aGtoH6IRibfLG3mQ8LYTi8izJJ7tNLUPxWH
gcuE7qodWNo4uKt4B4pPg2ofiLrErAzeb+GqaA/c8pnru9C1pRPdCstrpuDg3yFlIrGjhWgH0PMV
d1OjHI6VsXPkv/TMrTToCwEX8/qcNOsujk2c3VSsDDjJFDzStgF60MbIYquY/fgYp9piaSgJYoMD
uuNC0N7iw2myF78SUhD1T+ONqCo8N9mAmc4PDjCvQT3rLjiNm9hIGkkbTC3WnAAi0BX1ySRgizn2
WBUb2r6j+1S0MK1Jf+8zmoIAk44hTpzKDxleoqIK/mYfmC+7X9WmUDgWSLs5eireVB2Himw0Aczf
GVq4sV2ymxnz99nG2x+rTcKIgN3tpRIpL2EQl7FfCvew/73knFSLuLv3/yXvlOGaprUHCVgdTWEs
8/Nzllwy3tPPQYJ012QIQ+cjGHFdxO8gEHwKz2elZCG/fLJGbmrHOWbKeneaImDplQlPH/HUTglk
HZOu39NM9l5cq8y0leWk0bIVnK0lRGtv2ydbuWC2GCq/RoyGY/1zTC6NHtMcKi/qaStDB4Hou3Iy
NYzaFaVN7NYE5ZdZo4OFl92uolgL1ht7o+c+hNfJb5EI9xHRw4Mwf5WRrBFLiYxKLLKT3cL7STOX
c/fis3MN/yH8FEy9MOGr5E4P575hUJa+zobFOEKNls9c+yz72Dtz7u9yU0VWtY8eri9HvA8lonj3
sLhwUGLESiGVV+y5SEJmHzyRe3C2pWpOCWe2+ZvRUFS7YFjjsP3UbSLe1O1w0Q0aJliG1z4fcpFo
nP+WME28mJKRSca/wpM49LGWF3yerxWLHEkG6eSX0z4M/O9jjr9HwUobmjiro6KnIRp5AC9QrOpG
zDhanSq03wBPCbjQdzQhmcC1nXGwH0olnGzlvHysHCi2L345YiHLheJk2ASFVIUx/9lrRy80oC0q
sL3CBg2K3kr/jCj6VbmoE+wUUX7+wO3zqq0dVe/cbFKmchH1LYbl8ezPd5D03iOZoYx6BDQhnO/r
Gi82cM3xDLVG6O/9QZ0gJFU8xA7RwC40D1dFrQ+P3PIlEavbIJ1JumPzdvzgv5TUYQQ7or9mClx3
AJoweIoiWpDRCAOBU09VytTF6u7zj4mhCcT1pvzgmnCdGgXZKw1vgnyxU+XMjhc+OGUgKf3NIvLU
26mfInKv8Pw0XwwSr72oQHIjfQwnCvuwqNskhmWxGQavGyNnPU23jnaeWLkBZ10cNRFGrOBYioKx
CY/tI1zZnpPRJVJAFdvjwbv0yoMXxB23s6QaNLbvJjTn0dl8Nl+J6QBJtpss3LrdC2G0/6oAFhmT
+j3TUiopOTcpatvO0hgNPKmIauNwqy8aKQUMYk09oAhLjmcQg6h3HD0xOCAqJvqLf+MggqQqTeDW
kWhssJARa//HNabRGoI7xW64guNasJP2pXE910AKeELj/eCGmxFzSxvlwYSS3LJgl2gQUhGYNEdv
hLeGTNVKBDayOjMe2NbF5+U35ZOph1lKN0JvEpCo+PYWP+C/emKUOf+XB0BK1O9pwwHdJBMz1X7h
4ky+Tqv0l1w26dxJZg7WSQwBUeHrDrUMVviyFJj9CxuACi1wm3rxWqtqyfnHIZLZHAQI+iDYxHyb
f8dzzlcoU+UR39j0/UWluRE7yIwA1bEm4BpfiIlR9OHzAdr0xhS4rpzHe7oDrVdH8oOuQfIyw6KS
Udgeck/OyXozdVH3TMw1s55+/LnPxlCrRX+/0Yu6iu+G7KJBUL1n2fMlAFMBRahTy9lX/W3qSAHY
WdcTzljBj4D3yhPTGiDNcUjCE+4gobTb77fKPEMB8Xi0R3xQCbAl94uYGQ+CMlRwf4lcFdIXD0sJ
C8TtKXlv8JRZXkOTKbFAnaOctsaQdjKxCoZJVG+eetXOmXuyV6tdG8jjnQlJmTMYM2fXvxO7sGDV
CyJoTOW9477mUO8R9S9NSq5e4NYqr95v9fgHoQbtP1Ou0dL8b/0VvX1QZ90LnHd/cZUe7JewaTyr
+Xi+ib0FVRhyfcQp6wH2Pn79FVZrnSrGblmfa429O+v2055JUumV6/q1I88rxjxxjsPXWNkIaryY
l+EKQJFhd960MJObpWUOmDgEUZNn1OdDc829O3p3Pk3MMAReZygY3I57MhuIC7BJKTF8XJCMxMpu
q4SFvb7hR2GP+jxH/hMCfnCwCoEl/9VCQ7HYQD9XaPCBH2a145KerSuELVdhbH2DvJFg+lA33AO+
f6EDSnVWwBjwh9QrKSifGZEwlWGCmqpvqg/vBvrTLFI+tdLvmvUGgTelO1TCCspoJ7JKUkwcOyxP
712EYWHjDdNkat6RcBGt6CQ94guBZIih5kaWGHVDl8Zr4Y5LfCwbQzKji9JLeEs4JHcC0n/T0Lf7
ZSZgoLdOoXb7pMBEjCERE2X5i9j7w8jk7Wq7axV+BuTiLhXh/RRwvHYhc21ik45zYGJSa84ceuim
BqwUaxslQdt6g5MhdBnCFvCtRjfh4/biBoJxBjycS4r4ozb7rLdyJrcGYy7/ermtU6j4Qc17TNWk
Ojw9KL5t/neJhQ6PN4T4RHvYwV2fFw3vdAMMrBl6bWdcA1DwFXVV1sMxjjmTCkPNfy05OSvkcu6r
Cl4aDfeiVzp8rm+77UjA8RHzSY2Sr1EixW6QYxzf1C00X7sAuEC/flX2RhDH+HemONzM6mp5vEAe
VFiYJeLd2//TDuSLaO1Sqt0nALK/q2mAF3sziFFnAkQKuA/HQVKM2TV2xyVXs5xILxnMKrdr+P9Q
/08hfJiUeIiGla5kRA++HkGyBR9i8uxpU5kx2fK0oadnUl+ilLMbD8ojYUYGtqn4WJdHLAf21blE
P5xP47UYnWkOkTLc8xv4oF0bWVpLjorNPBvo3n0P085b7wh/S2scCZ1ykYD3tDmlzm5AOZ5xMVvi
YAgE+YzmduXtEYS2kRAfRBS76Msu/DGPQlxL6EkETzQOnyfe6jHAeOHOloN+vw+lwi0zhQz2h4t0
rsQi5ZGNpEzc3QRyIAt9ujD7V33ifXoyxfkz84/Rbdelgl/caGIvj8LbOuucCjR36SAsdGwZTbXZ
+qJICQAi7SSGKSYQyBfva/0Vts9fOIAyYGu2EXwb7jnC5nGhoeGWD2qrNYozyT54jKXujdV+PfvQ
WkQVWDQEFxk045D1Z8fLeszxHH06PUFZkIqaekuquYf8xhRklPXsoaimqh9coEBtVyfczlhi6YV1
fzLS7kJrh8F0kkLf0hrIX5cxpjlYnNwlyHwClL9O2xyfR5b96Hvkvxm21yzMSFcm+BziWqDfTYfG
mY4SaI6P+te4tYY9atLrwTazNwIMrcSl3LLKCItY++bFgsSgqyK3ekKA3L/uFqWqzEqObbIshDwR
W4d81T4bvYQ4luQ1PcnqHTBf+qZUzQ6RN3xF72aCeNM30CJ78NOltjKrJRhPscl0gpj2BFfI72TT
X+EFaJG3ZEUWFcGSqlhZ2VOAKZgF/JprfGj0tPgceWsqwADhMIES7qtZLiFWKit9gYlw5xxov/4f
YMRWjrDDS/ZCuFdNlymDLB/GbkwxenGUEeZSekJAFyqW5YCvOhGOqJ3/6Fbl17DDpfytNS4PfD2Y
wqvPAocRUDl6kAMphaCLTIJBFNojhSudDmM1C4TqbVmxl19kKmmjQX0ADXQZu0bplGxbdiZkt8Mx
uJyARNBwcRLrz5TJZwdMvYB6zsUawCMo2o7lY0HQv0+9MPp26MNGq5si1dSAOU7tGeDT8hcivOjC
BVJhWYCV0b2aRYLUbhc7BWu6zm4ZCOm98gTNTjZoQ6uNSlwqTF1oBFHcMg8C5tG2sfdBjyZdUntt
RPChja+PloWO2lx1bEUz5X1U1+BrKO8DKaagvJO+STtzWJSR8YnyRXATyZ/nm0FaNLbk/uHKe38C
NkLBFRz4i9I4dtflzZnn2jVcCAY8F8v08gRhL87Q/xit/DvhwDXHpotl5v+FsTkKkCH/rsEYCZip
xyKmtA8WTLJyMOQ08X46JJaTogSUAnI4HBRlIBOD7F82cIoqO91lgha0QJ0+I2FWTEGrzOONXOIi
3Gw5dFyHWAXBRwWJHhBoKDzMGjhfwBFwst5Vanh12AMz0v3upz4xeMimHvheP2fRvfxy1aGCBk3w
smCDPmZ5dgcYsQyCgM/6O6QdIQFAWqKya2FGjaf0TRSACfMd1C2c4KD/kIISbqIqMb623uqUjPkY
AahCaVQAXCryY9aEcvA+EZLJQOPQ1haOYkNbNJ74/B03HgDBksw9OHltR2hx2pz7dANS+p1iBvjp
q2fRNSQqo419JRme4t+VKCBL+BTX4NELCz+2agGHYXpQei5XmCHj+dnDFxej8Fy22QsmE1aMFYqJ
N7OYJ2x+E0Q4XhFBiU8O3/7KQZnps4SN6UcV8Ra7ypUEc9KdtkY+kQMLldFNGlkMAMOunYvyWj5o
eOg+e3QlkucFuMu/Gr/gXAebrpx10S2CcgM36ApfIf8CscfJjdbj5egviG7ZhAVt1YbagMY0SWOE
iEFftHfjAFpJ6+GG2mr0Ecdruk2As5L4PK4x6FBn9MO9VNWiaxr0+/SkF985a1d3IXqqzST7bgir
6K6YaLW1A9uLqHua+M6qWBSZtdvVK7okegzodYVRM7nFFILD7SdSxG49JkY6UQRmKuVbVD7242jv
BwfNwwz9co0zttRg80pQbocC8dDmhi0PvfHZBrWe8FxOZamv2NWUdAWifJUWTQFCdIyn2sKeDnxW
2mYd0luLS/AXTmcxVOGlmUFzLbibysLfgo1EXBHhVaSqbILCFJP1RwW1+PNrds10WfEnsZI4dHFo
g9tPsJdPrva0v+Vc54GExlV3ytF/BZpGNYCetJ4NWv0AhAMEAwJ0qP1yUAvLSEpXJ/wrgTigvFai
ZLJrvWqTNYdSx+8+5QA2zsO3e2KMGkl8RTgFjOztHRiip+KUl2MeE5AQP11eHjYq/ORNJTGRJiUK
r+YwXeoUi4od2LM+wb9eCbof7bh71ia5UhyBrP8bJj3x2OufGAim4kly/Y5Ips5/TbAujQ20lNXr
HTJ8r8WotlYXf/ANLkuwLvc5mD8zkrDBHVHLAZrmpe0K2qGfLsgjjHCD04Sns9K4lUGuVvs0M3+w
fU4St+EbW+U/Sy72017cTT3HpIRwSGgdJ7Ps4O7jbFLdtJcmVF5XugrrpVZfBo4wNHrM6+nC2QSA
sgA0pGDqKLxtKX+7GHH7Sz7NM/2EGkkH4g6q4yLXa4I53lLcnOAAOZV0gG7XyL3RYNafuvnKD96+
2ZFUcxiBpUyANaoHyGn5wxaLb2/8qiOxUQREVYCxt7hLHHi2jQpGf59z59clUA4OKlL8vLehc53H
LygdTPDt6iSccp15WwqygkJfolMuQQkLkiONuupe55G2D9LlLOdybSpRnTGBa2nCgfT4aXkHH9W5
19HmFWS1fsr/TwDzwna/PbWQZ9LdgS16jLRUfddlaf14CUGkxyQQVZ2H5gUf5UixNrHYC+jZtL0o
GIwsTtjPd/Tj2UiipofPDzp+s5/FnBu5s9n8UffNr5hpZTCZ6hXSbu9SpaGsqw6RSsOHxjo3YlTI
2vgkFGk6eoHpchWcO2TgAcXTn3A+ZVEv4YTcfljtYkcjhKiCFfWfxCE8p4/xFiUIo7VTT8pxwx7H
SomdfcFvNJp91K0VRZBa7tGgrsqruDAYo4Cb0EzE/D5JJlMD8hMtuQoQct4DfM54DO/mi4Pbg0J1
BEG1zncQr1+zo0HIKGp0hFsGPJfZTqqbeDTGnIiIiQG8rzGCeIZwapUEV+WV+DHz/vG4S4FuVajL
/DtzVw5svEl7xw+gPHtYXZWKKfCIsSK2JG4S6IewD6ssPlSZgnF5Evyz4WSEnwwXqxzgGSrQe/Xj
zDEGF47BLDEy/9MkXEweS63Jy84WC1bJzP6KUNr4F4hHNzEWrTZIDiVk6sLanfSap45JXKTDKQF7
qtjtetDlcfwiNI/H7Dkf/8M/Zth5ulkZQVt5ll/8hRP/PwAehrwDWANf0Qe9kGDMbtGUNgY4Qqms
JJ9psRVV33Tr2otFu2cblcKgS/FU2GwUBigLq25kFfXeBcro2qc67AcbjrHWN+Mi2z2GhvFrZZYz
GgsuqX4UeadgzaYQByfyfhLuecXQhga911EqsAUV9OCMv42ruKgOrLRQgLU1fLGiSUPlM0IUiHy7
ssP3WqpVvSoquVzytL+3Qz+FXfesdiFz39Vb9tzCL1T6ABmuhgI1ZiOYcSB6OX3pxdCM2NxYyjDt
gpsV9AjXJg5xYOpiWW3cDYx6LhDDrsbkXKaz7jtiPCcmRv+RFmLPPffipZbLHMcCa8YJPWBvqOt4
cmH1+/D+zW7tOsQljJiccUoEAoHIb3DN9rzpFl319akWamvI4tKDwunAXdr04lsy8JWt7xulJP+M
Prl31RSMSl+sT9h3sK1saNl+8qfxl+7HSoSam4qY7lfXs9nQX263QRtrU7JxK9l8CX9hBZ8BCCKa
8eOsWEHFIvLRsebzbYn006jgmWFPKP3B9UuRsiGcKfa7kOIbTqc9xGggTDJJfH1afghXRXrCY2Dt
YrQ1KRbMXxVZkvRCGImEEnaIur74zz+KmRyDnnDc1yztsOzD8h8LWczFg+5nr1dGsbZMUUpt8ifS
qDkoTlUJgItfv+rJWS/1y0e64FVel5j5Mkf6UnJ3TV/MacLbY2QxdxcFEoW4H6dICSmxEl0cfXhk
iNkpGhfyL0AG7aw7ml+F6bTaWsT63GVpOkIjkOLX5LkbkU8HaRtqsjAj/1yWcKFCG7bFfEGy4alM
FbiNzUicr0ExDMXrbGsRVXvC9ewA1/nFxmSD0QYjxNhOFgr3A/afl12G9RSQ5RB1ogtPlKrSUKXO
cHQiWDvWoJIQnSzmrAm0+9C2mfLvEotYj04kCw/auwQniE9GCC0zlLEpPam0Y+vAsHLG4etSouTm
VpGzfIGUIeS3Wl1vBdCgoexytoB3c+GtJrx1RkhSBxmrCmonAAxVEqe7vsKG7M8fjmJsxCLb99DV
F0EpJTviMoTNTMzJZkGWfpsaYplwSERrQ8UesiCj++DkUnhgO0Om/HaNVL1hFOi+mbdmWfpQHpie
9Yfejjdge8VUHUI6BUUPHk9dwAsSM7rpFQezjRr9PsL3R2a35TMyhyPP5ScGtpdV5NUvonN9+pI0
XVxqPH9zYkA9TCVsqp8twDOwDOdHd52PYg9hN0H6VZbemPfTKLDD8w9QMiH5Cc4+kCDdJEjNEiTy
k48zVRojWJ9vyAoH3vWh70K7igkXHY8QTIddusYnZyMz7sxOxoylLjwyfSbk32AsPWkyVVEoVFFn
QYpbT/HcY30Xszs30RVTNVRXwiREFcypi7pYJVjtQ2Z29vaje7ii8/zN0L3b198h+IZxJBOvHJAt
g4xeuP0cBURIauPct8XEJqYSzAzvA7dFqx1tMMyVDx0zEvUgQgkSPNcLbH08LRwOvlVFx2GMXZwN
pg7kpvk3sXwH6AI0/2Oz4jovFDZNQYesolQhjle/E1q9YrjnjMd6/8sjAhjzgVhox7YlZs++Ub+O
dtMFSw5MIkGQiRkbb5U3JCXfox3L4mQnTBNKixUPt34SANcih3fgJbMN+bMAPMziYueIKPXbYkpQ
RT4fz7Aa+DI3VHJrJ05YkYVZqaWPkQTfsm7VJ9Nr6SV6HJFJ3q9FXTMuLpbS28qdRSPaeuB6fVyf
qVruE89/IHBarlWy7Ndf2mHf5wm2xyR8EIWsabQi4e7Svy+xJ2nRcXsY/pyTf9KhVvDmzEWTwlOV
7cbnoHqzg2V4sFyPjEzfLU7wpCbH5pAUVJ3R99718HoAsev363BXLSl3t5h/mztkCzRJ6XzwcSxJ
EzS2KNXvzzseNZBiUXnNbim0DKdWTFBryHRiaggjJJiC4Df4jBInqnGooB0CCxA1n0aFq/mEQcBG
1uRPljkKwsUMUxERTt+JoHzr+U0riqbupYrigTj6UJADZYexpLxIeIs1rG9TKNhaAM3JyOWdhWrv
ulf9y486+IUi7wKJwMEdkkZptpZcmDvgPQXh7WB+pjFva8l52MBb78CoBBOpp8J76W+QD7C5/LLU
Ybm3G7S25K+V+OPe/bDhM1QlCxetIiBP+ocLDiWk+KXwiTKTkvMBWrCcDIOTpvbTpXpQDALT4yyA
HWJq0tYSJmzz+5WjOxLm/0ZfE59AG21P2Fm5QpZ6f+GAyRtwYAxSfhb+TsiOwVvUcfj1lfkQoZg8
e2yhDhsa4rGEToaWyvhgZP3Tp3Kmm0XnaXpxDMZaAv+YLojx2qRfhaL2HXpCpe2phfjDfuDTrZPW
b5ogIHnWWJbBRYQZyEAI2rZUzd6uGZvtzWLk8DKvIEDjky8GyKsA+hZK45u1mZItynpQ6a+QL9Qi
tHBqV5MM+BwKT9WnvD0/44n5opxLkw+LpdmohsJhii8zEKFYL6b2g0ShgbQxmKWZoWwcxvO/0OmC
osyQ6Zpo2Li8XOQq+Ir5uSaSDAKpIbKMYapIVk0MCWSAJdI+c8uYGAofRZ/KObpUOPHOabJ3C/7d
sRGYYxPqEvI5VST72efNThcyOV2SI5heTn1uvTu5QUqLorOECQcMhAip98O7CF/wNBrp468KRcUt
jSgoHnxpuMEQoVIVZ3HpkfGzTDccjnM9hpZsuy8UcRnqVwRe+1AaUd3S/b6fHY/nZbtp8e2NGPnp
fCTgjcTeHQL9mxaZqDCwiGK1dz3GA6FqlrEvjAcetU3P/ioJSAZs4plKbKqWIMr919RZkrMk+pbD
qHzXDiokaldxFLS+F1FFgVvootaNyc+SEVJqg5xMGfnFVeWHqBqR8F6yDK/4V6hZ04nAGw5kISUj
McB2v0ESBS6KxsbIZ9JmDtXKbi5DCsiXg08MHqvnX1rctfVNHSuyOQo3oVFwjxfYzUcS+INNAa/K
cFU+YFyzNKa3qjxxY0xhPKgwz8/WQJibKc7iU38c0k2xrQUcPM/AzHwTwbOrVuVIDVFfuk+QOiHZ
urUp3d4UxNow/OGGm6gDYC/Xb/k/zWvhQojCpr/NAaytd7vZ9ILyleYNielz4LBGGKz90pAQ24/k
q93KI9mlPqvQ4D8DBvYupp5aTg9o6sK2qcM3Q5rbthZq4EIgsjnDgXZjM10tE7JxNDLXfFtTuoDa
zLdk8smLM4beb28YoHHtWihAzJmj4ZlFq5whiWcuM/1vBgsHJsoj3ZU5V43C56Pmnqfa/0rIUiJt
lsrza/A1IJi8AaHvosViETrgGF1mrn/CQurLul+XmOx7AJcS1iKmkmKupZ8rf9OIZD+ioGluoluN
fdLwa32K+hypB6x99ZCodG/wNOBN+N6rY1WlORAKi33L4NT8lhB2ifQ6j0j/T5ihGlLAI73ULnu+
R/AYqGj4utd6mNIkGlMk2eRJd8Onp6MzlWFN5Vm3uzHuTx6d8RLN/ygusrfgckWy/sfnSbgjkSHB
fA4w5lzTSm1ksZHyI6/PUMIZMhtkMHr58+60pu7DkOk+2sH5FKhfKKxejVoV7ljBrLG+2t2x0klj
RpZZDbkX45dDkeiRV8Z+Pp6M/9Kzm/vq5QAU3xsRAmraOL6nbwIKTaCQfQ8bA7wUxEthsG1h6xXW
l2ykTK/FCsdhRkAkdVgZ67DtcUM/Cr7Zxv73iA+Cn1X4tNzQp8k/ZlD3AJBUDt5UeZ4MjYI8Qsph
/k1e0aPCPvRgbRJ0QaNUSWtp+b8r8mR8JQ6NNrMZV2XqJO44dAhF76oQtLObyGdeQ+pjXNfihWe2
dQsxERL3if/9ttNxDxAtlGiZ6QDKxZJZlYiDwd4PAeqMpHjmRxI8sbHU0ajUGiRl2vhNmzR6Rtau
ReXaxfp8LyhQ3I9cjp3PGDVEo+5io4tgr1AyOs7QitGbDO30tBJnOaqVOu55MAhhGWHIXmhg7/bI
8yWh6rpywzJFfF5SCvofcm/MjtNHg6k0hCjGJpUrsj0zN2x/bpk3QhBZaFYWIwU+QFYZhG/anQcf
qrnXeoliiHiMcT8t6FAXeKCHUl9XD1GE8rdgdvLikT3IluNuXNDz1jfPQ3QQuA0w0kfmxHJgLwdj
Vlv4Z1xFMdNqqLSRsmR/JA8D1SCluFkN97hVJucP9Xp4PxwGMtiWdyitqgIUMy+U+EHGQH4Eot97
FrHNXAKtSobQhLnNriJHX+cj8vbADvMf+dg5CNPrsLk7IuoUOULUeqNaqLrzApYLaIEwdN2Ohqpj
f7sRS40RsVFMxHLUnyhjOYHuZtM4USUgt0QL0SOTZtnDbe4KMHNtbLQZcty+yOVBG1zVdLG1jFVg
Cmvqv94dP1t4n569hmd35mjSX0llwaSHvK/P7vA1O8SfCsLsBKK+YlrewCs8XAm9KbKjaySGEngB
YfWDt+LDRuJUOEQQoiyKtEFgz6+KzpYfGoqGSgtF4RVEK6J7VHXz800wr234tvOWb54G55yf7IqR
DZ+LfwXK/9oOw4Y+8V75PkIXE15uT9B59xsSJpVV088WsFjKJ2A8Hp5gOFjM/WsKUH1Dd7cjSoPw
hCp9WhjJfN4wQo1oNAu+FeN1cUomRLxf8qQ+kpFz5JwuFk5V0vNF/lNGlNOPvXaRAs8va6s1WQX5
QrgG8/l3STH9BHB+UWGIv0PnMjsQCmBJiNaUN+WLmDErg02VICsVlzXihns+HJOOsUsMI7Xix0Yz
Y7VudGz3i9rzxNxbnAhMx//9Ul3eqnERjiljmfnkf+dry6CfHK3Fj6fzS/oMeW4qikXbF25xsfW0
W6meokc58i5k14+YYz/jeRqSCYPiwOdSEuUqCCDJG3EtsFBAVdOvfHWq9yvlH/eVedd6yMsOTHkq
m5QmF4/r2n2CDJndSJGOyexNfKPntZwnsmpIP76ZoJI6Qn9m/ohC136xJ4dLhGWqiOGHA7kmFiOX
036ppPM6oP9qVlwEUpNQ3pKda17fJq0/rFbwM2Yi+g+lvhTN6uT94HlCAF/wp7ap001LPFulgGw0
fvwZFsv0GStY/rOrfPIPwYa3DpbbuOw3BS0PrpiSVh2gb24GR62XRy5C/plocvCwhIWoq6LmgvXr
s/hz0yZ/kgteB4VhSdj7I24m6CiX/X2CkyaU/NSEoaZ3Mdp+ttq12Ap/VD9Hq4A3B7xQtD8QXAYR
fv+Uwa3IMeICdl17RtOG/eS5npo2DqWzAflB+CYsv+RpdwzdLJJ1IgAA5nA3FiAGzI0lgcOjlhdi
cYJ0JJ0pFgznrekZ/BiKlSJmQJocm2irfPCuSi3ygYRLZnTdXrCQbKFRuB+izCqvavTPpr5bYRNc
CIAdELigFlXZXvrOLOeAgIOB8eE39LMBQ9ooVOwzTwwgUYlIbBcyaVefTF7XAidQ6QjdkSc2sj17
U3PgYhUWyXr24CR8YsXaYHFSTzHOg8g4o/WVgILcYO/N+EI9gc6XYIkwsWzM1nvzMqvww/IoCEI1
wP2z+TvCeR0TEhza1ZNPRZLrTZyYpK10iZxCO9s3fCKqXLJq0dlell3Cq3OU9ZRKllIQJXh0SiMn
Ikgv0t/D2p6tCcrhyPzasfk+Ypreu6SA8W5CRJYav6PPx5F+GUZrQDpJIZqtAsRieqQokhFx+E0Q
WGfqI96lgkdmvSf3vkpf1OMDhgXG1iyahZy3M1QzaA0TIOkHngBuHl+ZyMqqOxDYekqk/xtjXw1S
C24sb3rmzkeIhrC/sj7gJm1Vn/uhkTyE0W9xqsXL+om/ocZLeGSpLom9jBHCy5xlNk60Xh12Q0wr
52Ngd0pLkTAMlqujmnFEidY0urZwiFqYlzoh4XYE1dHn3aCTf6NNOx0vMUq2O+Nm6KhdfW2F+Wp0
UBEsBufwrdRgd8rwHC7oaA0aC6ZkF0aykY/vmJ18w4zzO76EZ0TL/Qo27VtWIMpVGOcEKW5Y6t21
cTszg+FwNbxi7pKZKif91c7Te9ph2Y4ZB7MHdlOk+OXJOwHPBj1xWgffbqoKa9TIXtPMSEaef3B6
X5CxJ4lAT5KUyW4/pEMvKMM0TPzNaB9MhcRfaQtxukVy4m6aS27bVkaJ1QHEjwAVom+wYMOg3LPh
TXI9M23XCD21uXgUrGjtD2wiGGK6VZqroFl61tC9ZrF1tMGB4GT4t28R84aIonqUKNfa3Vf3qR21
bIXKG0SRIkaIeWCRfMVlQcMMMmPrIC0VQHlN7Fldbjc2EhXKqGIOFvPdVuBRsSEd3jUwnOu7qC8F
4KaiVE2VDbj/Y1UetIlMaI9EhmKcjfnGUvbBL/e4TPMt5INnzil0MsvPS+7pYzPO9HHAFdUFtTaU
uSzTGgsE7q91I8GcAKURQx9xgLOxB7kXbk562VrQyRgVoKLivcEq4JRUSDMGzCzSjn0XEmKVQbbg
VkEobCPI6MVjKS3hPumP5ffnsjaTPRloIrzrAqM8P2Bto6IN1BOYtxBGjlgsadTuwlUIv/yKhJlr
o8DvdlikqTlMgx5Wu/2tMy0UtQnNpwWrThplExQDwuIqN4/ijh1t6qhu+2yFjfrF/WI6gST0D+N8
gNkZkRQuKKCi5mj5GKm3FCwsCFdJcuaW7UExO0cttpbrFObhDwAIO+LH0uOoBjsEMvQ6ibNP+EBm
Io4ilSBbQQ88oa0yj5tnjf3yVUsjlKPYlhTXtm6GBjhyosbDEapSYr/5Wig7v8bYIAfyomI56sl4
VllwYLBQFox9CyiMhwscBfTcHs99DR74ejnjIVCWg/ohl2hA7bzTa9NtBu65pGmFRFgOkrZgRvkN
bKzEA0iJ2EU5z1QWHqLZvdFkrUN9UuzH9BqZONmlD66/I+XvUY6tlqgNWyzoHJ0njiUot8G1dsYi
0pabGJVlrw9pbDCzH18NhZiwXG40Rj9z3lDZt59sSiDfmxgg4Bs+SGnx7RMX7thkBWaBzGaU2eAX
PmZN0RWcOt1foTwg/1/KpZPeuq3L33KXXKZ9jSNm+SHMOmSi/Kwf7OG2PbsHamZfUHYEELDXRJHC
jtpL7Dh339BxPUGaWVdnRTm4qfaNb7GYBQImJCDOZgAnWpkDrGPaEujhrK4jD0Jt6Hoo+MlKmKAl
T/iqy5f6OKYhpAV7SlhNrr5T9PZZXMKms9HLcXb/NG2JpoeB2lEI2AJycGK8B/Utjo6zDJnOUXgB
V9CCmIfDba7KPhmXzBR8a6esxCgvBoLFBCJYwwGWHeroXJ8PPeWcu1UTikUc15b2CR4jav1Qw6TL
s+O7U1QqeUfgsgCGh6ekuumsIFQ+ViVaBXe47gahizOYYYKgYrK3QCG67QKqU+phViDkuY/ay9EF
ec4fC/HT8v4PGpwhc0b9gSGJulFPhrig/Df5+xvT98utRBS8kXPM+f2NzNh4yqLtze/XI7SGa71o
R6dHRMVs9B+Q9fqOdEdC+o2ETDYNuvzFJSZYJ8vDwvLzG0koa8jitHTIeOkR2JGjbe8vI6zJ5jmh
U4S0XA68PoOJaY4kkBpvK7AAGK7R8xmoictyfzWv/NbI348EF0Fw1Fl9OlczwBBBNaDxd+t0BMQc
v1VA4tC52cjqVycG2/HqLuAwevB2MgDyA3XtxuIEf1JeqQfl/YzugJBcPleYMLM2MA4Djc3VMao+
x/bRiFAfK1xyPJv01xwQXgqfb79g0KZmBQshUx3TDugm/DKP/0K/S1Fb9FLnqkC4ttdKYjKBUbZF
2r2aU6g84epS9JbIpoBsMIF/mQZQZ8JZAIm6VC3Q+s+Rp7pVY6+EWmeswd0TRAVb60+z4E7RwRri
wt6TWpzHXJTVurJa40Wlwu0RDrYCvV2gOWhoz1LOBBb7ffzVkCIQMo0rOg2w9B1F6DaJk7SJNtFz
UBzLgD+FldXoetj/7X74hb/1f46uvkB7mqAOBWK9YkVaqeeP2j4wh56dS4HzaHCys5b/zedNHGUw
6XvSFzv21HPaVGwwdI+LxAE1GkKqCa4cSnbEmQWJg8iuCnfK4VY6TlbzayNs6ClLtrdmZM2YRXMw
yP+qSywcL1S2x8X5/7xNhCzuZV4vqbJVag0q+Pt4OpvtFhMkNSCer+tNRIw0eNyYXi3KFvZ2h2/S
gj4k0hp7PfjBXpu9pBD9Z/u3dKJDs1uMHFjkWhrCJ6loAGpN7nY14jdipyDXfuj6XkQo1eZ8agvA
Nq69L/Z96XJPdKohcmxdb7DK2AFMJ18DVnGJ6MpAsirbjqyAtmkjWJVLeLL/dnInQj24ix54YT+J
5+xPwxYhnLoq2fV8g7T/GicgUK+u/rnWj6+GmhADMNzDoM3SEmcYn8CRaX15qEly1oCjp/8FHfeK
3itaJvqIQaKPnhNv17I4jTOwxkgAnbPNDg9497rCXPZ4m7HMTdEkQHOIaHoPk/aTtb2DaX5EJq11
7OuiFtHsfBrId1X28GXXxDjSmPzXzcLeEfPj1jxozHgMhkOr2lH+Hr7UKSPieQg5HrorfO+qWa25
flmwE3WUlKe6RgdLErG2nBYkIYeRnKZVZcpbCfZfOzYTaj4539muo7jJzYQI9Y3nBfTQYu6VARhY
45+P68ZL9twuYX0DzE7V+vwErsbjafSc3ilnP+0fPULbqMEpmnboQVC+hEljJt77qcSCCTb7PkUQ
k1zHjA4o5l8dvAhqlTG5q6BGA3tDDGpRO4YYP9/7KGu5f7rg7SoRiS+Std/g45BOiHaw3Uk/zXgM
HGP0i5WisI5IdKZx+SHpa8rPek97Kc8m+Qzq5lTA/a0eP5gUyuyTHdgkTbGNQZXu00O098chOBBj
7jjx2LIu+GQOWiG8ZKvhfADX8bu++oeLOh6AK42R6uKVs92gRXpFX4yOna8LCMtA7thjFa79jC4Z
YnOKfqjZaamMgf5zUOK38i274RN11tw7sFJnIuTFNceCAr/ICfYWRYPTyJsRcWDGpIyJnGzyEYuq
6WvYdUWGg9x4RATxn35DIZDt8NvKgLerkwbuXIQuWh3SqOXjDoKmRSTg2qsNvyjT4HBEPZ8Cmsfi
4DNtJvuchZb/kdzBa8XgJjomowtwwHx7coHbVqn8DTTus/sRkPyBfnYSqI0Nq+LnceWMK+wzqvkH
xbMywUeIsZ1xpC9U/8b/J84fx8PsOV2lzdSL7Y1Bhqqmx3HppArCgcaLW/eS9CKn8VnQ6KKM8o7V
ZMqZgvuqGcWgC15yh4xEGRA+qbAyLykfLOEv28NeM6OiR9/Wm9uw38BxLu99wi6xhL7NLAtNj+u2
BswKRNE7gPYzjHqb6ypXTv6ntCmglKJwKPp9/uSGmGxLQd6DjvJXDgJ17uy3ZJcB+ue3DAQQuwUe
cVti4fjYT9LQHzcPvtiEYQKQrX4uNxuwT8VvhEPDOxuycuWGV3suRMLLt95cZgp3pf4YtPjvX2Nj
1hFqYKCk3sa9p2EQ1+UC2k5ASm1r8OLpaZXXFTab7cjw914xknnLl3GTYdTjfUe0yYo85vytilgW
Sb4Herduj7DpM0j+8/BNJDI/BSP8Q93VpWwRSXiFOg/3O6MqZy7k0wISSHr+paBJVsHhebB6kvil
jQGQRHRzttWurwzDVdCPpDD0uCGbgpKgR1HZmXNO9YwNufZcmVHIG44t4g2eqTlULxfpmkooM+6U
DKUyJpceN+wui7/9y4ZqHkdoF5oXJw1EC+IY/HU5MP4XE9gd6JNoYSFP6UcJIrx/EB6TrSk69knz
vhsd9XApogfp2MnVVoSShTGf+Vj2kYjIGGkE7ejONxA1JYqVTXYqhel8U7KIb8lWp/8xhFBqgUso
tt8Y/V5uKu5Pj1hPSz0lrTL00+jvLEYkJfd/NRAWAWh2cBIxfkXNMlD5ucyK3UO+21Dtk+Ke5gFB
VwnLELmyN2GKKPaobDRigmCxhVLLwiBGyR1Y3VLrja6F+G4IrXdAlR45D5CMV5Ocpx/dWlZ3wqn/
Kifx2xUuaFUJR0iYyLkUwAHW/N4Ar+FQZ2PLe3h4GMEXx15Pwe/Tey9t62ybJodKfOO+qRgHgNIq
lup/2LjGiRrV4k1fm7wgYRCRrgbD+URkrAsfrx74tSe32NfVlzDsypVmcYN1ks+sGfYoKqTu7YWh
dDzpN9M7EfmIRtOSVSYKrulaz38g6UF5oIhk/jHuGX2i7BqAq3vrYYQlcQR4pajMjEVmz4ShsCbo
iSC82MjT3ABFMV1A7QyxKU4VJKXdKEapHSSK0tMnOzbKcZUDkLD8uptionUOo2drWTeTjko+2mz9
ysrjN+S2tBNZQFwPcEpqWUYnRTmKIsEniA6fmHsHgwCcPb/9czGm5YN0xbIz8obLqGLoYd5qlIvx
ceYtf5GPhx+njI9h+aKga5uFJJMUWzz9FjfDbzNwzcYrM8AaLPfweewVN416QUWSta59t6LJ7Rg9
56nen5UReSKEL3PedlWGtFvarovJ33OCtAS6E81W3/bYFScAh5+HoNPANNYwu1wl57XTEZBOsPdp
QSrqye92Pa9EZoZjR/sZN/vOG2nYqx8Ti+tKOvTaB/8J/hc8bbzjMFZFWhMwyC3+TjaObySiIWNs
07grClpLnokrN5FeToNC0bL5oX2a+ydj0ETk8JhfxwEowg21HaBD8IfFszqPmOuuDd+Ue+3HFrAW
xULIjkXedqnxPFCYEnhU6LaDpKhU4SSEbiAiK8S9D246QaJ86lZxSoBTV9uNebRpK2TZJ5w7JxI/
Il8lHq8enf8wmv9BIxmTOuvox7ipP8/eHo+IA/BFCqKhFqsI/bwyXM+lIwf7AABvNVit8nP9kwoC
WbNyhvcbfWoK+LA7GxlJMnBT3G1l/rlsE9KSWsD9u/DqMad1iT5zEDxLqFdogBHaZFIjf0ZJn2+F
I+s277euLFKMkODJgxMlhb0+v2W2urfARAeNqQELxO5WTPHKGi+LU8/zxAjvTDY9Y/HTawXM3AWm
nU5dItFGNq0KXh0zJlt02fD1/w0dgpr4CRYb54TVxAcMc6+CT70w/OJtmdahSc9L43d6zhxw0Chv
axsJjgjbxM8oSiE72t3CsNa/B5OopHBYfiGb803WfZ6afkLsLKAwkCEBqxDmNi3F5vQTvlAEuMeh
C7YI3vsfwZd3iz3BUc4FC3VozH0E/75xZKmRxnltdyfYLajrm4DlB867uM8iye/YNIovyIpyoWCr
oDYiqzXdi8mZtfD8Rn26VHfPeVxWadmuEHKtniYIobQD3FZp2dU7Z7h+dNnQb1pTqV8GA2/BMLsO
AFmvMPP8zbdf/pg0TunZ9mL2NGW6Z8Rsm/MnqEvlD6LO6APWpLGvSUruF1z3xDKMAqPKiwzynD2y
8GnG8PAdqk9qu9k+zS1PmN0rRwoAvwMkHJk9tfoiRyzzfOoscqWsWAlbIpYr3B8MsguxIOiV/GL0
jNtM8x4y3hHhmZ5huKSHt2G7q61+CY4bLwATHcdYT66V2Y3dEL/xzVpS88W9GPJ3UbDIXdnH3TzP
bZPRxBckJ5vW/pIJCR2YRS5HnTPwlr26KrcwzPzeXqOFpcLWAQ1QR6MvKY+hKHe4tX2R6FPojDwY
Cm14WuIIhx0yJxStvdyUJb1U0cEMwDYy78q8Egpq58i0BXeW0FSf3TghfuyevCEa4DuoztHuocN6
UXtTNJQ5MjbOMaAE2Fqgj+P0u2YxKckZCYLrNykUAzylQ2mcLxyK72Nv3qKyMDDf5V7+iLsDwxRi
IZJ9z9cbuaOmVdev0wXTtA1WOzPc81WGRTwntRSrczFC6vrEUwrRSXzCiwMOzT5FSdLZQTBgIx2Z
YizSmvQTLXnJl4J/Yrl5aXwm6PoZhCf0r7Fk4mF5K34UR/OnJvmPO7noBSvnUQPChOwHJaKzo2Yw
kXlVX4J7QzYZNer1EPTvEQRv/Y0DEL/tFjQXvxF9d6e7VE7s+qCTPyAgSENiRZ3MUl8p0n8kkU3w
Fb30Z3gLdYKfsZL6dPE9sEypT+cNLjoYi/0eE5EuR4d5/FulZCOS0AZfdYaoecahziObx/Hkv02U
FH2ldFMdMsY21w6sih/ipTa0dnBEVFCD4y0hpO19ALT4FH+ajfnSTcA8B2LD6RGKvWi2LC5lS7cw
/Isb56xWFpmqUtdaNS4Vu7KIb37NVV3iJCo0J18w3gFi+/XhXTWc3QrYYJlxGrVCvq6ZcZ0iKAXA
+xMVOeRIKl+Hl2Xlr3PB/mZN2Mk2diTJ2iJkNKnqGpSJoMDgZIfVqPwXcxVvBT5B3/f0RsV6pFGZ
INct9BW5qdaKU3wiWy7TuCR3/EfUsJ90I1Eb+y0p/LGXkrMxrAk8tvps6a7d6kjNMHFlCtXA5t+P
u0MvNmkUSZznkKivRSg+5muohKCbY+aDIyZrzknIYq9uOzUxVBLPK6YrATXP2/FTW+tpO8jlqwM7
2Vya6OeAmuGlJVBcpeLm8iujlYeleB6QJyAqzYny/Y6w15fqZytIHplwcXgtKpHN4DPgyNmh7ymG
eJOom5kPPGwCdP7sHecrjfvO31jYoGZE+8wPFEREv3otzRZhWW7YGWpNKpfxRNHSYAcZ9+iXAn+Q
ozPi0n2GpgzRju7/npfhifpTwgQ1nwpcwiQAWXH64r5pTMDQVP7RFS2CwdRXjYIkwfOy9+xtA9+0
qb6UxVZmcCSuNVfgeqETcBU2lAJggOw+kVMM/hNQG8oEOjkZVcNmZbqzKkcAk3CXpKv4v1NBYbcC
N3DaL1LN+G00POgHCp2o6L6+WnANOqqf7IUf7Y3aIJcyz/LACzLWJKdQf8P4Jtm91gm450vmSC9D
Tx/86eP0SM6nIOHbTpr5YhfwYLlNSmPQIItFcpN0wKk33Q0v9rVDFj/BrHZwXoU7IS7zL76efbP3
V8ImBV6uK6RMdntRjYVDXRB2h4XTqHbukgkRZE040Z6zjzvpGe1lX+n/nJMq1EIeiAVIpL80plUf
Nf43XVuHf+M8N6+QAQis+sy4OaNxewxOptWmFxY6Y+TnhAzkvD1HwEDYB0PcSurN2gCJ18EwsvkP
0ydksn75McXdakcyXkDKjObV4WDL3Wox6kr9QTkW0u0SBLWNNuT9r/5Se2a/i1dTZlXMD1dK49zh
TwPsmVepP2AkovXV8pYOtDmRwpjyXmEGSI3Rko4Yb+RZwgnBsTbuaXWxZeeF6kgahYNCpoDjw6DN
eG9dXliW1VSFn25QbaJNAtstScxYv8uIFKjDRjo8wYbs26rj13qGvzRKP0J3rukZ2FFPcQVI8y0r
T2APn08rzkpMNOshmlw9a+1o/F04u7BZp5F/g6NSV/6F10XouwRI+odU3iWqLH+Jc8VsthkqKRhP
liAfAAynNKOIJ5uf/G+5ptK9sl48kDQc39ifbBVoyhkEChWlTvcmC07OT3iBFBS3uIBl2pmEf5cG
PhScZwC+pOsaoy939OGUCx63GgJ+UbfeuZ9ZZgxfiSTjIiO5QYdj0KdoEG39ZohdYGp5HgdDJDGh
4GidfwZsm1w9qtpO8Xly41cmZpY90cFlJrT271tuNdeShvFkstc73oiTLmDXUXJ+NY2mkb7d58ID
iGd0b1pmF41L+ylrCIYkXWSqUfdh6hgjdnG3IGA2tRQgzub4P1EnozaA/RuUZ3gQqLLNBMDRbL20
/JF89ikB6UridKS+xmm292fXoeAaYCBlsrKIzbylrkbZrfqWoLhfqExbR5hst98tTkpckCYTNPSv
T1Zsar4HGhHPIIy/+2ePpr41wiWhA/pH0jNz/Ouo1GBCgpFBEKcWQgDc955rKlVIZRUiwQ3dkHuv
lx+fLaXqbiizs6bObbNlDvMtZnl63DHwNaJxLJgZdIYqIpKeFnsvAddBPM7xWAsYSSLm62pXKdMW
mJOpSHF82Ce3rRMHXMZb4yv99gB9uwFCdvwx39h0u5cuBnCfiUqExMacrSaqFYU4aoDvyYgXUsQ5
hOpzH527jFf+OI0nVxCf5jlEKFH0Dp7Rmifn62MJ6hT4Zg0D9k79ZQJ/KkcwjAU7RCNNjBieiNdO
VAv5hEDbFpcDiQRsFigjCO60pD8G6yWgoWxgZ/0t2VnfPgzr2QixjDvS6/vh5i3J0KaXMj7ohR8q
/Qx5b+Y440ld1CIOvUyjTLTwoaoINCS1Uyh23vMghLi51OBXP6p27X//XBNySHdb2JF6xfzlq9zZ
/GEK2yXldNT8tgge2dj3ky7ofbKDwsjEperayQOfo6PnS6q4HhVGBFswCR7fL9/XwWV37r8iVxT8
/k7+6YbgHeo7F/8MFY16rFmtkQuFAQ8n22q+/Tw0uLkRdTUhvVpQwigbhY5uGP6CB4KBEiK5oasz
epD3mXWen/MyLXI04emmaWgmpYspoNDCbOKG1LKujQkG5U4opW+638GWqHD1XBaS232SpkuF9l15
q/NWXKeKviY0ZwwPkS1ind/WRg6mdmLc5jDqbBiwJxXFBFdpPWpJqjL9x1Dk4GThCOTPrA/bLC9a
9CHTVsDMKrQ5kU3Sc25yKCRPeec/eEr0ASDW2pMWSIN3mei5IL15nkxe/XQaFrPy4OSt2GnUTGZp
ERvb2ch6ZLFGKjyD6AjJJjyaWS12P55KIyN2QDed9TQhz40R5krYDSuw0S8aHkEeAObFmu1hOaLa
MTswVpOZ4xnmklpxU2Gb5Vz/mdZr9qeDPDbDB6LXoCShtWMi6aV2N82i1uIqi9L9GoCRKg5oiNoY
RB6/BEMnAjz5FH3zoUwvnF2ARUz1c8tUQUREbe/eXG0wRA7jnq252mZ5IcDAQPDoQjVRUnCfITlN
a7Ia9pJRKS+fSRjQIKa9ZgVicH5PavPJ6Z95wgEo9fWbdaujSY6HIVDC3G1uDNWXLaJ8jRK7WBP9
Wy/TGYXRfDuHYb1k2p1iIxU3zA3DD1hL7dL7CeiiNgUnA3z1RcLxeLHlG7Sc3QNkh/d8kHoFFFzN
ZcIEFmOr6RpdEs3U6hivcBsKHKL4L6pfaMSTEnQIygO7/0P+lACu5S0eTk3RClPFssltvWxx6e9x
ptFoV3B1ethxbKPJRZ1Q+VpM97rtrCWMdEXfjZ9AWZx5H6VMk4RWJpIJSoiL9DuUSPyxTI0sSWmO
zPPPUn+dxmwa5iQSBxYRVSPh3zQpTz0Z8thMOkeYhemAdHatVT+jhaPYbbU+z6uKkgPAsjqPVzMX
0I/suCT1kK2XjMOoK+r4PTJQGp3oQdA0SY6kp4czgP/HoKu8zeU7GNVWM0QURinetugiMYhxkp67
CWkMxDo6y9Pe2KWAIIL5ACytopaOnuGHub+eaDxeXQamLYAwgraRrc137UbwbiKCbQ697Pthnciw
YUsmoy3cDm32K6Pu5E3lFbMRaImG9EUfp0EXvgUUuM+T3SMELqxSmEsSjhT9CIfiFIa8cuo7VGn2
Pljc9Kk/DVFZywvXMB1tmKrSuPxGliNnjJj511pqzi3KlBIb79nJ19lBFUje0q9zhwcs43cVHAlA
EP1oixnRUSISmD+VI7xgi7sPpur3nhBuk1MJlItrFdspENqjbptcbOBIV/HD0kvl7a5KukhVEofP
7TM/sEv4Kb/eVOB+jcFSsCjW7S9+Udy4fLCFtmhuZjTR5DMWTBeJMhEOnNVZgueYr0tIALLoQdfa
29gAjPL7G/hymgFFkASVyKdLMOYBR9tk7CfIjmMExT9UhFhBvBbgxq77A8UOtvlvlao8BhvSslaW
unZTEYOOzNMseen6dtdb7m9oqdOcYvl5ZOIHFn60YwRKXSFO49ex20HcXayWhj7d4dqe3NNp7e1p
ZZliu6FSRywAClbph9Wbcu0xypyg9XlU4xx9jEGpbIjggEwrZxX4g3+ac1q/+AkHdirWZ0YzmfwI
GhsyqNs4ftaukgBmoSenfZOPW61aN7KVjfKi3WbUkKepD5hDKgarDXff022X6pSMjtvnsfLtxI+n
cS5ZYVHoWw6xR2qi0w+w3WwBcKPiCFk8fn3NM8U1o9unm7/Knu1KHeWTrYZosVQhQPtLuMR9fRob
2d3aySgR91ujIoBOMr9RTAF0gTXg+fzh1bdrE+wUNjdx4oV4S2qM3jdpZaOtdS+gF3RLCafGeWqb
FrXCIuNa3imqaxzEwEaiOBT8kDC/dvo19AceD5PFK+PYcne8fLDN0aAP04zFwjve9+bN/zKdu8e+
u+WRMaSAzEzLKZGiMpvI1jXxn57H9aaQ5YbsAypCwUnZlHXu67ZxVmkQYtvfINRku6AuR7cb6MyC
MSZJ9jwRHeqAk3vYxN3pbE/5qeOIpRzWkihxIkVrtNQMIlbmJfxxbE4ddzOSNvJGPkXG7sc5C0tk
xS7a5VMRI02f08VJyneIAsp2j6hYSFT28n7uiLfYbEKj5Ps8qAu++qUsLyX4yc4LTv002cZQbjuy
K5V68Klo6p5SBGobtJDQ2IBtLI+A5cV4mCMiV47+9YYZWHKGErh9wB+my1ebIRPTQwJLih2ddf9o
I5hIALdMfgNdtE5ZTzJlV53XYjhObLgo2OIkTgvLZuYKBd3OAHZW4+lmDO5VXFa9+ywSgfaw/y2F
7pjNev0vKzBRf7PMAxTFn5ElXCLVjeHb2Ly55JuZfH83MWywd5dhjXG8biPI4i+BqhtYm+sCixNy
uuydvD8mtHKGXQahDhJi0MmSH5P/KrgiCXqhbE8cjNWBdvwdCeTnFBzjpPM0PXT5LJZhWUPImm08
DJCWRuardyd4KAMMGIsOTICOQNCUoEU+WUWiHkekSxg4eS1cfoXRXPRFXjtdVxrWp7UkM/sANuP8
oTzVRSfOsQeJ6qs+ncw0nKub9/9CqsZCbXEDknBKJiptBWlXGH2gtiTurezwhdVsSJP8OX3BDKTD
ktW9QGrEiunKISsRaS2ksx5ARJeeyCV8H0I1LKD0YstX2K05MnUmQCxTRCnWIHNsPk3UHfuG/F9C
seVoPKd0Zky6OBp7DY0vz3FF5rB+CVnuPPJrYIYYHKhZEzoHlIJ3egeRaFZaKOmPrVZsoM4I/wxy
dhVK0FfgrTqTteKAQmkcqrejW+hbeOIFUN3h67Gc2UzZB+Jrav0OfVzj1YDm/8+b/IWJpfLOIpGQ
d3ZsgPtxt8q93JMv66bM/u/tG4MkV5bhvoTOEsyQBQn3LhD1hOlNkVtpSa1xo+aRGMGVNEeHUhMO
SYFB8YQHAWgw+afIEGQ/RwXHlejE1YeGBFKi4JlAtj07wZLPMxI76vX9srNhohANr1G4sOLrhCE7
9OuKepkPu599uJTOsVzAdI2ylvDaTlsqNGmQ7Qsl3gtFYTLN5sE8zWYmVdQnUROYStYM5CfNdtmk
aJPdFwH+bqGwUR7NYwBwzUNDXYP4wp8p/IhxzNyy/WKzK4aL9qROeAywMBW1jSF9Xk0QNe/LTCCt
Yp9AuKk3e9IX9/8+Phrv/FkI0Pbb23iM6nEUE8ZQMwcQSixC5+AMsl8p8/3sVOq5Sn3Gf4JfXOOh
rqSHI7Gmzr68uKLojAZ7YqnaWqPQY7zHEMKLuj6n9aPzUBJMw/qkQWXOmZyRr+aAaFSTpE4ogvvg
ymTHDPEtB+KsMPPEXFvYbbSQAN0DBIM3oIfwIKpK3F7i0bMj56nIiuYj260IMzF3Be+boI1QZYaV
VP48PpJaVsueHCTh4q5vaXvRPiuafMr3kQ31hPv6JZs5ljYbo3orQfHm0OazJhAo1qRZH91ILtal
txyA3b6JNYlAB96T9dR8n/pES0XHVaZOJGsSkUxBu2mzHUYMWb3o4tSH0a3eixyBHSEl+lMz9OtZ
EF15BZTNtqK9/Cna/BDRIxRtFXSx+1k4mdvihtgrhH8Co6nErMECXs/K2O7+63RqXLErmRZ5/6E2
E/PML3UzbLfr+qwZmX9lG8XQk2WtbG4PtN3TmqvcEsBgGsbmTalpsVNXo4gZ+3+wEO4+lFnF3eha
V1HqW+lCF6dNR8Z7n0AMaXioVCb1G3Qo4+LuRbfQHe4Y/5VKrVP2v1eCZCosKLjBwbKiQwzvaahB
NSNafDCavh88umif9F9dO5ZKET6TRzzkCKAuUbURxRtlRvoQGB47peYwO42jVC3Rz+XIQnKA1xBw
GQM5Y+O78sAPkQ0XddNmP7LASHd2rvjn35FZItevFAifAtKiSdhvy51cZly3LkJWslgNlX4hUCGW
fsqRMuJxvlxqJUCDxI122Ndn8nqybSge5yHqrxOz2T51gFKhX8a2DP9JeHenfo4UtLEUtF4Oc7/T
uEXfVvP63gKBsHvwE751qufqRHMuhogkNECEAU9uPakmvQupJz5WuZT7pGK9c5j/dlAR0NOSqrOi
wyQal7VniU/uwd6uFBgkVTWkW95UeO/WuADDRyB5adWmgeFdLUq0aJWqmvxMCWdKMfrMM/f635Gf
cmag+D352WlGlFnJJfuSJqq17PKLWBJ3DlSvWjlsfVjrdoi1nvXzI4kbB9afDEtNXxjGJIHrr7Pj
grhbfX/okyN9HHGKIZaYweHjT1sNY8TKuq/nXL1aXvqeeLt6ZNb/s8ABvO1h2NzVNP0Fn8wBjPYR
lW3A4lzfSqAjv67tByFhwAQStEbIgIt3fgaVQl6htU1efxQYcMaphecCHXponujUFqIwAZu5KzjO
Rv6u57Mllfb1UA2UfG6F4Y27XH8uD2c0kaDUm5095sEKhReZ9wqQajDEjvBqJ4Q9gDotAvzU9ZLu
DnY1TBYtJQ0fgReXC0LI8R0uEVnrtSsj+GQ/ylrrwnAk0oCUTC4AWuABtlrjBTHN8GVvopBkeujN
odSsOLAzLns0QX0hEbvnzzUQSJ3c+eGqMNjJuwFtrogzr+rh7iMkviHtLs3ypLrNwBRNFwVQ4zKu
xBT1kwEJgje1iMv3C0ok+A26n0ebnoltrcmR0MFybz8urwjCIiIQTvollbvAuYD7m911V0JdIr3a
1JUpyIClaMyhIw3vuuf5imA1COZ00GUq47yc5+BQ77SlnV11vtklgIZHxR1hNkVpPlYbUaK4B0Ql
+LxatofEfeY5nvUOdaKbwG8KvOEijLgBtGmSer2EmQSF+CpA8P8AkSxzIu0gFcJTKqIW6uqnvLxt
NrJO9ZjVJhAsDA2XgnKBPpQnbRV2k3ngBmhO6pQP7tLVHIYdcbdTtPVGhOHPNciZtNrGOkZeUzaQ
721Y3iRg4xLGeYuKTu3e5cpQN68uJX4de+XDpOzyIQN6baaXhOenB/7UxzZStV1y1fFBXKikdcTz
6QVH2pK/XkMM7ksGCPsjZOiPj89gzC2mDgHqtZ2gmmk8nX6DUnRy/deIS6sr0qWPN01QcZfijbY2
KN+P4Yt2cvWIml+JC2HTjoamu/pWh3ZX5O5D8KkZtIVaVZk6g033r5nF54Vk3nmFQfJ8fL4tPC1K
oIlp2VQwZvZQ3aJzwppe+UEJjtfjv+W3g7qyS8h3zjRwAMwZWuD8Nx2OoLImL3tQkNYCBinp+IRI
peCLwJAtmEDVGQDPShbKeXJ628SCmL/4ZHYx9s4JRPr/jSgsCSxlJBlujYbiFlhYFVtaUnOgZGKx
dW1IJxQXQxW/idlGXvFU9xV/wh/iFAUDKT1lXx8aNcT/Hx9RPbZlRzLoNvQxOuNxb7vGFVOb+Fh5
U3xzLakbazHony1XEctZ50XjUb0uCSsCT3wxtetinOPRUgs6DsGtBc8Tlj/tpj6h2q3TBmFtjGvm
C19atyJL09d3c6e+lSulttBG0qehjPchlyVFVysXlrbXvX/GJqhKsJZ8EGvNMU1ykcCA1GoHPdAv
oOLroUVn03id5Ymy1ENg3C2R4nXmIyHDQjaPA5vpIfa2y/OcJQWzZtsWNzeVe9f9ISd7COMU89P3
VxddS5CP6aIag5XHePqRoxg28RF3vnTh9tCab2UPOxajnmMxClDomoSMu5HMDPYsF45F7HjAoGYY
LW1k2+o/iyrkn66truYxjAQDVkHBSyI+EmbB6WEN9g80okwbYtZ5AhMfBOulikqjS95NxuIfhL5b
dfCyDhkMD2T5MyxBhwpsyiJ+h+/1MfT27cDxNs1CRpkGyZkH62jmk5nty6a8BfeTrQSlrc3ZeRkt
dwgZoEnP3KpC6tS5ssibai7U6nn0PcAJEVv/0S+pQd9k3w4Ltf1UJL36jWK+D0cEYhk3OZbAC+4j
CXsb8pQrUyxMJjlPRY9PiTLn2wj1AS4jvP2t+eDLWPpHC5cbKHE0RrMYvlc8ZEHWH4xzxvXvTeCn
PF5sVofpE5Xmc4ITC1OVk1/I06jAp60qrONsZV9TtxWH2saENBmBCpcwCqCkFsKM+xBzicbPU/iq
b3qw86gFqpbTfEagxz1nJBf5j2OK9Pp5uUPJFJKfqg0pOks9E3TO3ZfcjflGQGv2TWwGnGMu3Qsc
4ZbfAWVAyrvOCvcl+zsjaa9x5U082/QqPwLhyEe26riwBmSA/yrVbDTiomdDsY2rB7YATVfjR9qD
nIBPXP0sRh3xbySmwu+GPcpsbvuqVCLY/dLPKyKVKp+TolaPRF7ALv+oaMBXdlqZDaAEweACrBhm
yxkZsg+w2Sk9ekNXKBU8il+FpUs7OPWo7VUSm/Vsbws6IAUY63PhD204o1+zB5cQPmBFBsL4cYsq
0k331RUA7Hmff1WcR32WTyrNLD+iOdPX7toogxj+uzpNRQbIfZL3pKSOVXsu7pWhtY+v5K6b7AID
o9jLMI+g2THAvn7Gnt25kU9lh8qNxeRikbLrZEghGFqdAVOq/Vz+hW0Z3IOWacsZxZt8be0V25ZO
IQunwxsE7h72FFjomv/9SGsBkygGxuyQ1FL9Swa2LAz+SfUfu1WYIYEoHZo/4c1GFo6MrkSFiEkI
jSF+QCTwJSPv2/bh3UslDduFshkF9wEfgpO2TgM60MT3hc+QHDS+CLG/Ava+ipJSgA+fEie43tJp
unJlYY0hXS9prYfbT4KOpjipexTRi0vRh31mj0oJ/drSG50z5xFOMwYJpfctQLoKCe9+Y991jIWz
Y5XvUBI6PXuPbo2EgKSdDxC5B7yxKaCkvKfZ+wPfdnxvy/Bkbn80f0jRJUNgil/G5xj3d752+9DQ
K32kXd/AWB/UB8X40OmFRyqgOJyJxSMgSVCWBr7qwSVp6AXYf1+hlo5wXc8WFzuua+Peq/76+/QH
hIaPeHzK1LsHosAwoPlBtblUxVVjZxCWwaOvK/G9tTxvIxpCjumAJ1mcn0zUFf61odTyj6fPv60E
IbRpo+SABTzaigjWwnQUBXOmR1NAVdXR/jbz3lfOyKefD3vA320h6TzPpyf0udnjcyE/gBJZdWH3
OmvMTWuHwV1bo5Ed7PkJ4Mvq/TNbijOF3Sn33QSCdESdPAICdv9NJs2vuWhwwp7amVcLfjnDg1sD
8mFiLoiGNctzahnvk47LM8S19kV2hFjYeGLxizPz/QjfNtRBujnHm0wGjSG5MwIx8rl6n6o+Frau
+2zkhwdvtzHixyY/cLxxgQdo3q77UTxtXDXFeeelXICD6dlF6zLCTulx61RWzyAH+hbf1KZ3/A7N
+UW0WiEv9byBac0ksFPsdDBUviXRlD5BGOR0/ZlPjxfuz1C3lc+8dxIrzIp0goed2L2CBfDZIobU
Hw33ys6S4n5aXtmkFE+914ylzOxVT8plp2ITjfhmRt4zVKM9ORKhSdWMLoPLAH9YHn6KT00VACKg
jNeoxBQeHkwwmhRPfAY3UuIJcoU7ZGLT5IhFQewb6k8ym9zxoADmjB/KKaxuCznA6u91w24jCOQQ
gBZRapnAgOOf02y5izypCfdgpd7KnAGXE/ktdE0twLn2Lq46qSUxjnOzPf6Thatxyo8KP9xy7vD0
Bkmep0ZqCVvlFJBiLg8GtdfjS24Zly04KkSM9sktJkwkr4r17euPJtpA8hnTlOCCgMpHA3oN1KiL
q9LxVLdpxEs64xP7b2LZ6yj/ls5jvkCUmEBUQcoKj8EgtW3BR5esJsqOe7ySz0zEK91kXpw7oinf
uL4iK7WN+XxBZDTZJfq71mmeIJmZi6Yb6cDpgUGJ25iWHOOuz1z5UVhHz3TB9OfPox6pl80TxQGm
fHapitAD/DyHFD1PnpHGIiWkFu5ml5Usj3G/j2bgzjnTIFfXmY3vNer7/Tus2d+RJnhJXs2GmTra
C8HAtPQbVVz0lVYegoqJNyXj1EDir44RhaHYdCWYJ2gPnCffq2sCpTCD8KAK/HmQSasKFK54gdeI
5tuinNgvUtVWbMncKgBSN00VsZc2TUf3qWKDAJIxcGMGXKwAZRIyjzsYv41smalBgWv9PnSphA3F
aIBSczI0Yrcd1s3MD+d9ykhOExC8aAqSM9ODzMpPvYUwjojkjpC3kRHrAc0eEfq3uF3YGUFczLD/
rj+fJL2SIjUel6RXQHWpGfKkJgbxaW8zHgSRh46nByWK+cIhlt6V+omecSypjsss0bTjM/5BQM4p
wxSgcBdrJYz7Mfy531xU30P255OMv8eXv1l0JHz6li4bHB7VcqetWMdXwRurjZAmu9agbzEDDtHP
UjWhNl3fvdRY+Piffn10k81vahNHzd0T0dq6vzFmhnemjhns+Vk6URwObqXO0/ymSYJvPDG1Qq/D
Qy5OVwMI4VAwn1B5u1hREiR/LN6ICfVu8TnBMbXPOPb44E6ixrOwtwcYJcRmuZD3Ofgg8onJb1wS
TnIeKf7My+ZeaDoC0jS8YOsbvt0TYOCMG9jaBehTLh8R2YB3ofd+nJvTpKblsWdHyVV1oLd/n/8v
/bMSl1pwYdkSMnS6W5BiWVY54cQ/PGl/VONTHXsoymZn/Azjp/egx3SOIs1a8uzUoTKo976JxPHT
0tB8AACzH9EDbQjMLbdvY+r5SgwgNGnMPAzG9xDQ9YMWAP6fV9Xr2DrEbb32xDG4HjR7PpAROvc5
xYCQLr1cw0e5gqKKCiVqvxusEjLrgMz4El5qnToH6ZGaITdGR2XFu+gXapHSIeLMojCYR/wQ4taG
RTGto8WVwU9ZUW1CdAk2jHZgfwXENBW+P+uGx/ehFYgDtCmSei93ev8ViCrMFJ4oAq/eQASF3qq3
PsW8HLH0HOF5dHiMl3WCNb7+acQ/w9HkCcZMI3/Y6tB837vWYAaeCJsMzSBEPvbJ4cn2CEC16TX7
1DwOP7fRckx71zJHLj5aMJJDThO0jCQ3l5di80RP1Vo5VOdPM4PafOvv+EYFbQOs2WOYbjFhBv/Q
Bbu4WEb3h8lxd4x7z1tTcWPhaN7coctYCBnhYLLEsMv6+XgTgSKdPTzxpoFHRDhx9t+ExIICyGC4
k9tAYRJC+avI8wszR/rPvKJgcfFnefTuQJSyHCTQhoF8PoMXI36eOyJNWwQ3sD1FfOjiyQMCPxXY
OUyamY7AUmr0kR+qewcSy3PAvbxRqY4xUeizb1ifGIiWR3p6yrYgk2F2fWEe++DFawA9XJPiUFMi
01Lmzo1I08JYQ8to2zh6EZL2dD/XkGX0hNE0uuTCY+bo6G3StcdUbrBr9P7bf87h0gMwEKLLr9PR
izjBIQcAzey76Dub0bqLr945IJ1UAEQmIeMR0F3h6MEZkePVySwujwn1jR1WBBjUqhaD1NZws2XY
Yc9m4zvucnZFhpxaUOH++Ib61V8Nmbqzz4w7d4/sn2jKt5su7bb+N93e94VAb/NSdtRWvuP40cem
N9t1qfZ5rppufTywdCAOuCXrhWeXXqpyi2GclnbtbXYyy+gJVWBD2Zlesj3fAlG+nPD6tTntytoS
YjVLlypwpdrXqx/2hy9204F6qnLm8FSaJvODhrFTVg02GAupjmBkWKJ+Yxn3a9Owm2NuWuWUO37t
2Ddcf7h89KTTfbTI5G1Gpyq9sBA3od/HLnM5nXdj29FeBk3Z2vqIolrtY9bP/x0Zdr6L7LVo9KzQ
arOphlX0jqNxBvzIwehzQTs/WsbdyR3PA+/Q83V73rklllAO14Hc9zL1wuzZPt8X6jjhFi3GzqZO
Bv6WQIVZeYyCuGJL9BFBluu+SYaMrCRR1GuKlQkSwTpAkBGWn7kxcwiRqOPQNJbuW8hctsM7qqGi
pNGmVUczk0EVpb3BPtGAmoLPT6xzo+z39yELn05P3DrV1TW2Au4N5egJqW76+SznV76GPiUZC1TD
lsXRo1SGgBsEkC1uKRPhrHI8gF7hWHgNCG93TctBXVJamo4Gc4FPjFV3ke9r4mE1vdXu4YntYAqh
01BpMQJVh/kdRuPCDYRjrs5whhlmgMFpuB4eFFOP7zzwWuFlqKWsU1PDrwEV/56w18bZOCjOR3Mb
dZQruBA5r08IaKpAz6ZjzuMqL3l9bzdbOirDDW9qFfx/5Ja65B7oTd/kLoKD8WDoY2ibr7e5Lijh
E36xZFAst6dV2yFM5d11FqTN+SXSVv1MHh2LKoHP7T99U1+Re/8pqbAiEcyHO97olp1vRvBnYBMG
i6FhoS23r7FufzqrnXa9VbOnsoaPgQAzEVvCWmo7+etsfQP6XO/sOSvqh4lG1FIk1Sg/u9l8BFWp
sHoIl6Nr+OCteFnsjQZk2d/G3NjkpSugXdvE4KA6MSvwUKoeOvABw2igu8lfkiwsz4AlLZgKrPbB
HEn3U6aNLVee8gByGSvnHwoxMUU9Bp8sJtpQ0qzrNxsKzE0DAznGwZ1B1ncWt7vN9qs1kNGzSJxA
LFtHrxPm6/5KVGTxdomtPHh+VStj8e+RCaXU5BuBXk9pRepFemYQQDxK8R8HZ69WVCXn80dj/4/S
o/IhRL6mgwqcYu8xCnnn8Rd1xCe3zauzsrcwf4O8zG4oC+q4Kv7+D2XDWDxyQP68jSm9A4FMdQq1
OO7uX/0ent4b32Nz9wCP2UfLL/q6YreBgFnaYAKRVfcE3dvRl95Q20Ny82xccXm0UBrQyI32jj/J
yZHEqCsZukbzdsw5l7OflvbwDrf/jHG8cIZvFhqk3Iu3c7RwPa37NrNVJhX9efwFOv4TFiUgwDBX
F14dts2iSt3/zvgWSfPKiDKgf6NyFf9f5s8jTsLNrYUGK4lPhylPgrR/O338VGIC+RzYyb5RA9yk
2rs1BX5ZeGsCrbW11iV/6xmF853iKSjT3YHpaMMDJDf0+lDif+WiQ+ziORlvu0knB1rIrO2OUKle
+luh2upSISVNudAcCte7ug2yqg5lVZHZyB40h4afxEQGzn79WmGGZz6OqUM7Q/V04ku+sW0mi51X
+N+VBXsyKH01ehToABlt0GO52CrIXNHM/UPQaIXK1FYAlK+MR3Ig364rc6pLoE8WDDBDPaplQ+Yy
oiNS8nZ+aFe+xebyZ0aH+a0aknn8paL6H0s1LMvC+IpN7XRcCGYBTRkYMb69+riZrE68HZCeQben
R+0F61+4NcyWk8w2MBOEBKUnJDRE8NN6agyJZAAtmxnOm9RbJyuXNMCytnI5ARmE1pCQ86syYluA
wYvs/7uERRGcQKc7cgOz45+8zgLyDUU5hPrNYPbA2HhLF8c6TnEAGNu5WbADQgzWi9GHY94YY6oy
Mc9UeEfdfCy4JQwL1FJjgWz4UEcu8naU8vcggqCwE//0qZoSoWZKLMrM8KtDW7eoM92qwSDytBQO
xrtj3C0g8OQwVOJWmcWd5/XPmbk9NFfxZiIGx5rlxef3w47PDigOqqbbNpvuFZ1VlssACGHGiRwS
tDWb6Ailw/Js85E3A65JUp8vqKMeTg68BEzxQrHu9ZJBvfexXrzrAE3/Mj46pAQoD4kp+EisJJkO
1SGYBp2gy11vXc1WTSzSxz5zn93/V5tqkVp+ceK8SZB0WhEYbZvGv60FGBiCCKBX2YbW6uU1eJ3Q
K7QRh9OlOd+hmg+Cdsisz8DMZFIBFl8Ztwlwf1AUS7zq8JF6asnO4DpHrY5v2KMsO+DqX/1cJqEo
3miDxNYlUnsn5IAoxSpxQ+MO6zvUTgwRDbSrxtrA2YQDji3AxeBEw8lzTJPr4+eFugMvLuKZ3TNC
DB0vVjXbqryxg+Ee3K28Nh4y23huaF0Ukl2ugFvNtj4kABUFJcPi6F6lMmj2B4a1/DGh08phluWI
tfgbbKGk0ccyDJpB6cuYcoV7VAFkHNvTGDcfZLLMo3RafWg00X+5w5m1yRmgRoRfRtvzHQLiL96d
z5GeyYfEFtQTI/4b1w3XtPdsfIei+Kt0eevR7vd5amB4Q3W6+uUVFTeaaFlAfZE9+L7I4YaSDWDg
ucAugYkOlnqH/+4cBysek21ezY3zJXEep9YWDYR6IilATQGfzftwNFf1xmRQKQ/31+fOQIz1o8vs
gi6fu9TndFSa72rJpNhkqIpPTZpLyMbg/Am1IfPCEhd5XsBPZR+ZCZaKMv1ylrJf0lXwiUW71YcK
xW9Dnizc8frIosaVz60vKoVUFI5lr05AG8wzHifS4fpMbeITgHX84XwKTnARcqXD0pm8so15E/Xy
T+jpkqBbSG/7Mb+x5h8YwAzn/kW6CMMAzLInvWnXXk4FBc7wnUSvfiAI0qkLhUlL58Ev1KHpa4+9
YsJmztfd1H9qXg/EGESkUeGv9gAVDXafJiNhw8OoE945faeLaV8BYMk42YTcGWWeDs/9qOBnWDv2
a6IcMnj+XFc/5Ipljl6zTixPugBPXm56AW77/JwRxZXh/rL1MV+vzhbGDEChvjgK1SNqapCeSb98
5IGE8+dkPpzjvniQRP3EdVPHvKg4/afpru/vwZzKMpUrit0MWFNib/H6XbEqqexI8nASx4G2CShk
uk9BVklOTAd2K6bA3QyB/pmTCttRiqB161ObJ49FSgfmWCBUe+zJPpiRvez6MUp47gEgK6q9+ZYp
jHnnDurKED1gr+E0hFc40y30ZQZLopq6nz4Ob7nXEUcbhEyPjLsYll/kMA4Oa9tJyceBEKg6rcid
uQ9qCMFsCM0ZhGLRBcNyCwMNdEFuG1Xg1mFlQT6M8fWxGpuXiwZgXrF4pmtYvthV/uJaiTjvTFxW
Uk3UNim5bKnckrHPO0Bt5nYQfh3z0NjT7xvLlNQ7u07vBhTCgeH2V+p/OfmF1GtKLMiCzLzCFKha
csx4idQguODizyADMoY3Ci54XWkYWDC1cVnG2IVmql0pgZztuS5ZMck+F026sgFRMoKfiXFjUMGW
C7bB657U0/LW7gnCzXtylZG/qxM51Xu/JubAshvIi52/6d67Qx/DcdokCw91o5okcXeDEQzy7+Bs
hKYiTg67PEiIOc7J4LDK1sPpeWNDuqkBjwvj+uAdATYIFsJF+VlH902C4sAzb+UYVI3QvAY9pHfC
C2o/gxYOaeX+JH/cHPl/fH6ml2E/83rTC/50rVKN9Ap9smVLX6kP5t5csE69nCcRbsggNkB7iRn8
sLAoRSV0dn+8d+XgC83HZKJVnTnvPpyyGqO3lp0cBKp8NhPq7BwE6+aiE3aAauVAp4+C7z/fI24N
5Bk3cc+wdHV3bBE6IXa6bpEVClM7/j9MfPCuzvzvE3V6bNu5UPhXHL77I+nvgj09OehPBalZtfDz
/mMKJ0KkIjLGzSoyywtAKbwLIegyzCUsRNqrMswS3eYkUhYEEfdAtyV37OB/W1ijqOm9BPqulbQP
AFa9iOijzXHUWgbeqRlcdV5OtAbs0YOqNA5vySO/Abwkw2PODpmXiAzro9PKHB1OsB9NrnyxnxrG
iV0Tsoz8EWuKRrcvHLPfRsD9Jz/+VBOPDSKpNmg0xO7VZIhlpIXAflXdCiWSFXT1aZSZe3yVTyTZ
ufn/04y2gCbliUeS/cOCW2IoVC7/JSfte0+Yb/QsPHna6NvLw3p9um6sYIrmKji2RMqtWDIkmCFr
zXm5gGHQ9eDRnZCjw6ipe5UIjVwFOv0cTFd6CmcVwz7t0veGyXLD6iiA/th2PJFFmh0XC2vXCxmS
KlQZHBfG4rl2nuXQNYFzSLyDFcoN/uuTDwwOZSZPFXkdmw9n34J8WQH+WA2W5bMFyDsp8Dqehmsx
eOdDx+9p0cGNm4pySN0/JWixxD9Ti6RzidQtehpNEUR5MdRSS2gs5FoWAzsANydgEtjhpHzuKXaM
cemNyF5ZrWIydYG9apCj9ELEl9x+sCSQTFAh1RpwlUe9LaRaeaXPJFxLbxn0wczioeGtveccyEIt
6v/eojj4TiHXj0OAcddWF7u77cPNQzsJc0SNI7tItftFbm6Z3HW+JPHc986nSxzK7+YtbgXh6odr
lGH+9jdanq/3x/L86cLF4j0gesTwo+NOjL2yBxlsbwfaCP/xxLEfIzzADmSNGEWb1vRBnid1e50L
A2p0t3NY10lA08Yj432WVLS4Wsg07EYyS9YVgScAMiFoCirTMkzq6b32ISl1a7o8/cotmc1/lpl/
CWqYN+iw2fW+fqfZ3LoqPmGBrwnh6dkn5A9vAV/IVdcKU+Gl5OmEikkigt5KVmhZaIR76/yAjvfO
ylgpWtdmfvHgXebvXIu1biwdB7AQtVO1KKTEfES8dyGEflMF9abPoyESScAQlzeJtYB/oziklXlE
K2M/lgwmvu83N44OmotircJoifop70YhoXWqdMxYSNWOpfA4PW+/XCoxNrecfKO7Ym86oYQ9cTJA
hYvUp4lZi8oxhqIs3Oaqmcdc2eb4gQMygxAEBQv8voX7wsVILwWeUhF9A7N9xwlEIuE+JoO82nh/
CY6WpbYqO93jjxXuv+sUnTj8+LxYqqG+bBthlsaEC9sREf3mBFt7BM4bsUN3Jg6ArRG9uRIQFp0U
gcL/b+8NcCjBBJmhHBoBmEn5IIDDQB5k1um00w7a6ijzjbWjW9bfMNeA9K2eJnSt00ORQEjK+geA
y0XSiFJPbSLgxqZ/Aha74BcqB86PWfoO4Plj4AAFdSfcX/k4+Pek1bGZkpAHI7ycQCrUpqQkXMD+
WJwngS60ZP8+VbqwvU7leohgdkN5b/PzApwTuGJG9lC3ea0m3B25BrzvVz+5eZbWEE7O2/dwxDcM
+db2GKoFtaaIpQfS3XEg+y4FzseN4bVLz3xdeEDqqQw+VxVCTl7e5ZhxCo3MGX2NnmhwRB8vjq1c
wSWvgoT/ZKLGecIa5rq8O81ddq2MHPgy5M7mUT74Jg/RjBQWOm3UNrJwo3+05PJv2RU3OnZ0NP6Q
m6USpTmmpC5k1MmsRnGKhSRPGrLpSTVS97fs2qDYnkP98ddH7P36db1D/FGr6+fvsFc9t/wYRMwx
MJw5zVY2scI7x6dT/KfiRG1hhtbvuHj88O6/vINSaOntnva8EHTfTpu+ZT5r1/f6Em/WbLx4W+uo
WbOviTlEKDEUP047e70rlzKAtWs2FlMECbjl7HF350ayCNOStHxhq6cPMEp/dNDl1XW5IhFG21Ny
X7kSyCc72s8dUhyZVaN92/Y8f1yqWrzRE9tKM8X8HyrV50ZL885GJ5T8VYVhToqqOKLV/YBxfIf4
W6xgHgtYcVD6VIjyhgXX/ll1XAyw5D6PGp/ww8lRRKKN4M7Vr85B1RaXg7u09LMxiMxJRS61+yfW
twi8TgkKknl0+zE2y1b7ueaPod96k4gNIox49pv1f3zEEfP390wpuziTKe8OyUOasedt8U1ahjOJ
ZLpYxRXCVETSh0kWzcVTFNYTPcEwXlMePhZa3/dMLQMZBnMibJJXZ+X9lhTotX1a6GwE8NuiXo0K
T7bMk5nEtd/Qw4Ic8EVh+EMHMN9iH9m8akcJGv75bGev7ENTqhl1M4SulpmONZsxm6Qvieqx8n/S
JapSqObj+2Q2fId/wHyHRBLbiJpm+6oYrckrq5aaoiRPrS/FY2wARCk4UlaJIUGg0HSJCT6mn0/E
/jYPje5K48KDlF4BXxL0iaE8eUjncAzQyfVfOKo+bnVTt8NAb8s4LsMTWhQIRvySON7Nb89Wlx9B
tedoKAY1lwyOHllAOK4StVE3MLxC6nP4dTbfeyrTaxu3UIppvzzKxN5v7C+W8arobHRJxYTyqZkI
1oA3v7LAUKMPm720NVtb5EKucO18oMylNzkifFB7wfxZx1GoXgDuvI/NqA60Obf9zAB4wJmV4pYn
DffWaPdDSL4D7X+MO7pJ2qHjONHw1crKgZAkmly8nNH1jsHUy3CBRVWxQwgl07a/Ra5iQt7V8WTU
UvkcO+fTC6W/mm3J/cONyvrfCmDvvO8n+CuQncBjhdoxL9jyc0+ybnX2WRsOsnVR9Nczvkrr6DOm
aVMOlAu7dvNkwwYQtU/ndXCEJiprGao89cHnB4JNJ8yJa7KTGk24GuholrrD5KeYqttBRDmlxpKU
BLqkh1NZPRreaaJcVI49kutvSHb8KI3zWpppuCcgYHUGooo8i2Rnd3Xdn7BLSQL1F7umd2WEkoyr
OJUia5+xH4SdYPfLsF6LP0oqhIgXjkClOXentn056SFPVcJCLowfKxcpL5XOFuM6Iyr1MpXGk5k1
KugmRtFzUn9Xsri3P3kx+06yVEWzblviO0mSwx63HIlu7srxQcsnFzrq7njhYZoyPFR0sKwE4F+A
Jz86dBRyuJPl7MhdVjIsEAGNCtCHz3lXQAMk07RL7hZ86zQXZq+MVBouD82pRA+q7sbT2b+SyreU
HsmiZPGBmXuCapxWLFYxGA/RUzspBCSlRCeQeipJK4WYOokAmdsB4Fmj7OsX++xT3S9J42JRW64F
bRlmytQR+gREVbG2L6AKrOaxn4k0wetN5c2zPhHaBtqEuxy4mTx6O4lsPNoT0x/AI0Ad3lJ8HXAg
3bSKVxXFy/LSo+Oi4SZpTwKJq5Osdgt2gnY84sFgCw2HQUz6dJ61ppiKCAUtuRqOdG27mbjNVOC6
jnzf4E/+FdGYxTSuPRX2qnsPguVp7rE/MoDroU9+UVPTjtNYPesEbMTsGrRd826tQ6Mi8+/x1WZ2
//DJd2qR2mL2RDBnV9xmGoL5k0roycj+KSqPgFGVpJ59mRYVbKZ3PzHIpC6Ez0Oy6bAbDy6ZZqSs
IGMkGhPoSIqZFmr8+Jb0wdaWA3f77SIvyE69WcI/IILqVbvf8xweHa8x8RPpFpaEPE9EogBD10xx
2jpeL1EmJ4TIAlLhQVVNCwHWVeYbDQafAfoRGTJFosxE79puF88m7tpUkWpyqw+Qde4uEvdI55B9
v0AXlL8WmTUvtGbJUvVt2SQIuEFRv1LyoXJ1L8bu+UQmoR+YGSdT5TJ6bEbQ6l8w4O5JEsQBC2nh
dje+COUem75jwb3zuWa/ICjC3oecoH0uYEAIxbgrcMRlvzH9et1Xd5Mm2bdZ4CJGBAlHiA2q5DkJ
yghLjfH6wswoRDD7yKzeVEEjuij3XsdoYI+xVqPVmG+0Dc8cEtlexCYA4qh+683lEv1wpn1Yi557
uEHTuuvS55YjnXXQN4bf3hFm8FXl4puCz1Bw/jZPX5GOaC+CLowP/pkXbIiNjtebmDBD9Yo80BMT
DtmIuMwrmZsUrQF4llxmRSmRzaF1fU6m+Ol/CD4F/fPJHFAc9HDMTyxtBol88i2O4tcY98X1Nah6
tqf378eJ/EUC6xtQC1zE5R1j/w8bgVs1+/+7ex/l0OyiTn90Sm4ei6/2mIlxWnlpwIG588DNZ2W+
zYFBTG1DmRgoyA9nBrPxzLPmzO3WJ3FZVh0BXpnyotUpH+kT17mEC8ll2q02k+YLv6V1QnviFpSl
TTZS/fO0/8cjr5pFN4FK6/SVNU9ibz4a2hZj2QV0eU499rKnTElWWqW3qo0Q3N1ZpSAWGgMTSO+j
vRaA5/KEMj7HZC44Q0JWdHlg3bTDKvByNveNdVu+aJkAYjI4A1FHfQS73x/KbxcvWBu+7iCynore
Jy32CS5erIi0Wnr2l8UPeV7cJlroGT6g8dFTRy2VSdfSUEl7VRc2x82Y26QWQSbNAf0A9+uYoQP7
DU/VE4fLRt6ANj0au1pTJ8sEbZ4f+fYPq6Nnc5EyH3PjaQNcdYZaqdsdx/8vrga3xpe0d6VejOrM
/v1EOqxcRTLsZR27UdtQBkVxS0oh35W6tv8ZjJBlB/ucoUWWhOHbZJmHd7OR+EMfSYKQR9byAhLQ
Un2586gbie6lT/Y0p7RGzrjz6iX88hVvbZZDEcAvuBBZWS4W9edMh2+JMF65S6nZG6iXICZxDc8H
gTqCVf0E5p7bPE4muKRCcar8y44TrEzIzl19EmKVhMJF+neVrvOk4KWPoKehWu6rPQz452HpuFHR
QZGWbqcgHoHcl4f9AuJgd7hqDOXxa1lLnZwiyNrWZHpEr9vfu57oP8sJLtORr7S48Wli3wVi/k0W
Bbg2/srPSlogc9cV5x4czeoYFukl1bB6ZAKDpz21GrmLSScvy1mrtW/K0Pz24lTqxRYdBxO9IqDJ
pz9u5x0jXikOIJby8ghUTYfRe46DkIBO8vpKZDqdFSeoQ6j6dt8nPp+X0nXz3qD2V9G7E/EcxyXI
01MkETnVfyCY4/d52H5bPIxJpyQvulpvdJU3m8WCHftRu5rHowQRbHJBp9ScEsotNcX4FQIqXv9O
dO7QswakZz0KNxqpTCdVrJ4Lia5GV94oFOrRNNOcn37YxFSIM+fce8jmwPyY7lwYoOonGjplJSZ/
9n/HEjy1MUHr0WBwLrClpSMfHp+X7pbsobdENJDclO31jO6+uh9VbyRKel7/Lcc6TfAb0KnzEybe
XrH2N5GQx4QUyvpqhmZ+8b0SVSLUFw4ogKxpC/lam6D3uoU7t4coRPSW9SP85r82DjGh0XO2/S4I
DZzJdrxYRTswstQZcLVk3jRCyDojYz7r5voJlrL+sKKTIHkWd7gaH3UO6OmCY1D8ZQjIIGROuPpn
/JnBNSJpK7GTbMbIjVAM+k15sek3/L2/nxWOUmPKYe4YC9YecRTQM5/Z4jzr8EO7UNf3CfFPdtRP
TyIZAzqgQ8XTBafVSqMN+79Wy14WjIycd/09yGS4BYx17YLANyv0Ux8FEyCwWT2jbacIucdnOwp9
HROjLrYYotqx2l0UPIfgY5uuzxPF6mNJR59FkqyzSOhCnk4b4pGxQL2g/0dlGRclVCAkuNBydnk/
8zB8L/QbiXfK8xJQb/wOCz4mbeAhuKX25E9091bncSJFFDhyztF6ssEc6dVFJDD4cvvy5wtcV2xn
9XU3Bb73ARjKJZQTUbr/VzEwpo1skgCvHbtphSPHO6akhr4aLg/m6hFzsqrT98EZ+jcR++BvWJFg
rQaTionNvEgP41gzNqbs9v5x40bPMl/Tm50Y5f2jX0EEyPGhDhP2nmP4QwNVKwpONy8BUDjC5RzH
ccTlPoyMiNbLocgKdAtduFi3/7/jgpTYmR4Bm3SbVnZ9hf6qoHbUqWAIf+KmkcbkY77yb390Uo1c
BwNsZfW0rKh7g3DJXDTp+QpBi8GYasJ32fUQqQYFSIU5rwG55XMGjKObZsUKUfzjBnDiY/CZeAap
LXC1S6+gJebEptk1yssKi4kRS/hRwd5KMx+PeEym40f+z/X2IXxW42YRqL+VPyy7WJtzjma5nbOH
S7ldUt2y1ajwHcMmPfwNp/xS7L8cdPWGDf3VG0jczCRANgAxBwIj7JZ6Zez4HA6qabHLyj9ySEiy
IN+/T/IfqnBk8ORxiZUxZVON1lY/SJjxGfycqWIxEIGxDbca+hh2qJ+T9Tu4za3GjwaxF23wUKGr
Ru1LYyZ3e9ZdA6vIo6OB5SpjZAxfGWl9CCGwLrVhYj362zKvAQelrJgWSWYUUVjW1Z1/nT0T0T3z
ZVAcKCYQmhCc3fFAsXH3EU2q8qef7xLwzPIXUvYXVJMUnoUw6dCK7SKU1bMy6svHKkydMwZ9998U
dl/jjQeLV0Pepiu5lffs9zl084mDYNsaAtoqB25pz9joJon1M/oPM0rLrsjBDMRoU7Ip3zYKkJ9i
4PawcJCLf+3BKrpq7ubgtwJ/DUdWJ37h9Q+JJO1RgOqoALaEu7/SXRw+yT0jhar0FiRotdHkxtqd
XwCT/LpPKPaLrtx3LcY3EABMzoSyvyZzTGPOGtx+TeuvwgfzYxyYkMI9giiIDTeVr0uPNT4Q1EQ+
kdhkLjIA2KAcgTf7RUczKl1OJDv3V7o34jiS2Bjkc7bR2KvPvNM2NgaTGU0D5VbF7Kct7Vcp3t99
GpQz/bcaFxtb95bGQRrZfP1UHibptL2R9NLgwtfJJDp+DdS7LdWj+iS4nG9u3ryvUn9U/FPzTLro
Uc8UU8h0vQCIxu04hetgkPGVwN/1bxaTHVN+pMPyDTwHG8ZBOgPOe+pkPVoL/aiePtGMOpqFupGX
KxeKoD79zgWBK2KxqxWhm/yoOZn3cZEzZNiQPB2cMj5cPx5GtYcR1vMlbuixMkHxAyXVA8tLnqCv
BUUM3N6GAe7wrtlIOPfolsnYoBLZpBNytcXRfVBPAVDsJrswSJpR9xgJoveWstbnKF6RetVmn8LE
guTyzXA8RWY1p3m4UmyW1T8VWzBbrGIBniNUxEr7OUf4RraurBBZUR1mKl+vQvkNBkOutiI/9os5
Dp82umvHQ6NIYW37hX78pbp1OEf+n/1aXKY1kV2cS5AWYQvxUvLEEbQlNsvmplYlJxSXmsRJB/DI
EpdQQeAvHU1qp/NzsXtp9lze+QfanJzFPxeQL24Gec/FymMSZiXkKB12W+WX0oV4k2IsRwfdM3zM
3PYOajFE2BfwoyBB+2p7lAvChrB6rBxmoqsy4y3RcwRMatFNEtgMg5nzi0sNSrgfMC9MGPa4AzUV
uoYh2JBDkqBgqb2EFutdvO50VRd6D9LArABi18MG3+5MKyuVW51K5Uwph/+9z6xtOLGv0EPD+qd4
bNL7gW4CrICjX7uw98aIedJS9HuqN1/tRZjR4HNkTbVTqjPe+FQmik49OUGZC1Z2K7ynjjp8xrhh
XF6tLQ/UEEI/pldFr883H/0+2AqUOeg5H2etFSijUZVVtbVUyVQ0cucn7KZxnOB+MrrMBuUzT0uk
dsDE1t3wDBvTNc/AxQ3ThgDwWoUo0Ivbry3JLRHVvmhO6W/DvD3iV5zyNHLvE2XWe9jUg41wvsso
2DVEZPsyk7U2hKQax/EVsB/+IJUw2nQDh/mGU41pVNpa9YoUQjy9X0TyCJCqW7bPKtwXQEDlj4ct
2UcgaAo57/ou6Gs/g1Pa+ADr5UxJ+lOBmccf79k4kZufEraksjRznKmN3ssvgRaKBRL87j8ild11
Yd/7zU6NU8PQODyh3okJbNMc4VhQ8f11vCP5+DZ5LdOlBbdSoJMX8qLToJnBj+Fzo/7PhyrxIMTz
cXcaCjVP64FBtDC2eJSZoeokieIhuOSI35hLt4aVncu40po4qkWETRg+13RfHhqd83svk58EJUn0
Rd2Oy8frn7BGKNr7bnZWrceMaqALGrOtDX87A03mpykv3SVuXHq6YtY6kmrCNmwjQa/1gb7jFA+a
yX4lgs6dH3B5PuPLW/RmOffE9nfVIFCMQMEqOyppx3X0ZPTuOuuxLfmRQfhjWZzeRCGw4GziSWXB
xR0STruebnk5FkcUkUUMGgzorg9Aq758034wSlLM7ik9dT06GZOjyheZY0Bc8AtMLo48f38QVPBo
vEFCWocSR4ny3f5y4qWC0ZE9QSlOK6mjZodnFCl4SshBMgN5l7iAG3xWjjjz1M4Jk873cpLU+tFg
w1+crV2RDz5iBo0SW/5TIZwUiUiBBzBKItTk+ejC2yLn9bkTSRy0pnwKC936D9LwWUNRpvephIGC
/HowXNfqDbczwOyFz2hY6HYz68QekQf+AlxV26c/Uj8pJkl+6MAWLCARWOK+gwnpqG48ycG5A1vf
8qGiFSTvi23UItyvO+OICMeTen3ous9AHh73PRpj/oeSTiFn8MTNAJz6uz05Nnj1LbnKT6edisJq
LVcq37HvJ6s73IK6Grqj9IlyjLKa/nomVnpx7aUBh3v6nS+kOlwzszC2tlMZUe10Q0S3rm03xpoP
+VqEK4FZ7wv7D4Gl2kGR3E8Otm9PRapWPMQQM1KlZ/jxj/jvsLMwoTuNWf3PxTayCyp1iFUX3aBT
32+eO4LClzsDpMWf6gEjoFxMvp5YmfmP3R/jG3Z+bjxMs84HbNWyKA9IAWzXOglfYoxSMK0btvVj
Ljye9I8RO2zKWS2U0AJakiwS28dxOu+t8Cvly5bVnuWjaODRpqhrpyXlC79se+E8yXlGm0Opjacu
pOQmPPIplJe4WN2yVWyZDtnzHOoRGJFcJh+HhyHgHpuv7AHsUtqZ/2WM88Vd8i9LDxa+1aFCxkyq
U/iemnbJhxLi8BpDn3WDNuXRxoj5z69H3NWtYx3a4h7zwIDDV5uuvVA229JxDhQttgPY1F/uYrdK
0/7C6bNbxlBRL8+yh5sEZIaNbbzBUvxe4RSC0gzU/JTpBp7Gj1yqIqlIlDUNhZ6VJU4xAepsudZe
hsjhgarZjmazosjgbolUyatcCAln5xgmwewHxU71vP/UeOresjy3UDi3cGCUYzqGLHMq5IrBGIR2
UT9Oy08+C4cf7S/Uq6LYV76HuSB3a3TSKhC/gxJTzZQhtJaTDI411076X/7wa0v7jweFr75ktg/w
rUfqBkNSAEvaeEPKnTwjf2wDieAWGic9c9H0a13vL7M2qu+RjdsSBJjZzRZzLBAhCUzdjnf6Quea
g/sn3Ny6XzHSwfIkdgn/XySEJoOIbKCXxsOOSaSOyIbvM1zZd40xQ4BHIN1k1WDNUkDG+EifPiAJ
YAwhEZOs1g6qk8KGGCJ7ctnEc7Olkrqhw9oIG3g/wzNKIuNWitTckgclTJL5ZFBCSUCJ1FCL4MZc
NVyUQK57iW82jSfL9d20HXEEoP3eNRD9C4qImVPxWsU7yyUR8QHHDpeoc0gw0A7fIGaMRv/9F/nS
VEyyQN4Tkw6n9K0SZiKILQ1dbrFPaHBm4mur7g3KBpevzux3pO5fdQ2LznQ1WWWVf9jM6eNFZ3S0
BvuvCH6Tx/nq0/f2egYME3u083rHAYRICKsOgZDJ45jQ7uE5hpP7lpRWSDpCBhWg4/ejkYQ8qON7
5hlr7nrSw8xD5iKqcJGtv+GdpSroMnEto5cW3m7mFSH0LZL29LrLdCmFQ/6q51otmVPht/77GlLH
9C11Fu/8tS627wcWDorS3iRqesmxaa0Jaj4tD8Vo/nwuDWIWTAZGpNS8mJk2/nMAPE2GmvKU64WZ
e3NvkRu02SGuJ5i5lMNyvURrhg4XPCwbGaYiLyRqTKa4YY1aXpILSK2qFb+F7Jr4ujPMWiAAYgr2
vLfiEZfAUd3u1+zQW+WtvBTyOZ0hynjefkZ3TaS821B0dTt62mZU5L/2B2xPxLRknOkajS7aCN/4
iNZTjUjPIqem8ZT5ocULZ7IYllc/s/YLx/zGnn97lToG44eue2kJAQpXK89UzP1NAn+KfV+37qTA
lO048S2lL3QqEiJV7zINvZrGZygzVeTFiHqzOw5SOQI5wLBwB3v04fElli6rdU9gkEemV//E8ykQ
o/+sfHeDfCKvxYXmBrLWIhacR+TQicntxmspEv//sUtcw2OVtInnGGxwW+7DuCP4lR5+PClZf3tA
7tMzE6Lzt4y+BiTSP7ZU2lVlCNRnsfbeEC5Clm292K07bicbzW+Mbv2s+HYo0YTCm4OXdt7e0kQD
X7kxf0SM/LKPNrdRqWvtEtXr/PhJrVvXVdd5+eeMnirS4L5EgTM4qqtRAkUhk7fA0dKQOL07A5+N
aYO4wAveGi6gGrXRS+3E8oPzpp+Zv5rb/6t5j4P06S+EJGCOM/K2m2aFED/2wQTpkm0k84LdKzol
DeEktCVkxgfTPi7LuqeIurlpup7AQyeEk13w3c5uB4tunKxjulkCKRB4hfI4ajBkpV/fyUBk0zgS
QacweGghNOTBKNudsDR6/vlU4bMM7M1sCRid09o3U098Hc7A07e3QGC9O3pwHNURlkcXfXVCOxpR
pP9lr24RRpv2IPvBjhfoK/Uhq3B34pUHcyw/bTEwjC7yDoHHogMjieMHEV/HWjK5ZcAX54eZSZ/A
ZR3uX5NY6aHpTtKuyxOT4KQEYhj3gxmv9IrmHUA23yJ1RTeLKRh1LrUUXEB7SefaWV6+8p58cJqE
+FGKWUKgHJ1Be63+deFAl3m0hXyXHNeVuXxRqqiR/NNkjVqd06yKm1DKnoHVNVQyW/9ZQfPZNAF0
KE2T5VjnqdoA1W7XE48mBh5pSbHS9mvt1Kqrix6A3AkIksBUxOkJ4CP5z2/O4PjIcq6Ual3thO7d
YUR7ibtOVg6ur06Xlogs5tBzYTNkM19N5AKVygpOtKporSJjKA8gp6dAgILbuCgG7YhXiNNdgLUp
3Rg8+WfEZBaifpn6n4RC5fpeGdelQURy7GdOmGAgu3kXdO/RoQ4tkiZbo4v3IMu/mCh3Z5zgTldI
2T1Q2Hbjm8alRV07qjGc+DdMR603RORknnc1fLvVX/qHBmxR+5wmU1ODuST8+lYykbABoljHkY+C
x+rB7OtFcOb+J+OsFyST7wG7i3Qzijgf6ORhQoE43V9q7OHIhFRQtWvow++9rEII16o1ozXU8SeO
L7kzRP7z3h6IlUPx3kThxV/HwTiL3shaMPuYFqCzJ3UW/1s6v8qaLA4i5qHdBvlB3dBeLqCCdIcz
DyAzK/XGUjfjv/75jcRAmQ3CjeEXKxYRyqQmdzHVc53VlYTQYtF7519g8K56htFMloTmLfDlc3pg
VhoecEIH1ujT/DmgRRC97GYC67ee2cVilLCQJGi9HidD0ZehWVllgvyOGXtGJ+BSLz4UtagvSX3v
HoKSXLfb+yy5NN7N7XnoQfyxs1cNqWdyRsSBEZU6hppewAisrdPYL/jMDb8qJOWys8IvS7/iYOuN
dmpQ/6OQmgLCH1nYe205i8Wczh2l0b43yhDSWEOBisQ01UomYt45wPH+hpE3NWBDsGnAt8+xT01m
Oc7qMBdalf4pyQ6Dp/V+dFwLrVyfgGPECRgVPTadRAVEG82mtqErs271CEyer92M4PphC2jh3F7E
KNfKGyPg7qHrH4yPSIOryI3idLEsj8o7TddjrLlVTcVmH/3gtvqzWvhyH39z9oa5ydOZMUWzghO5
x8lCtTaLMKXwcXNL5aFoo1QPElEHllQrPe8KRlKvESvAQaamavE3M+xZ+q3jmdHQ8FIoa0n1ZEpd
LO7mefdsQIsmr3l7y3i4p/uW6xkk6S6xenTaThJxOcE1UaKb27JNty6g8HmrB4gi7ZFwgAVEujIo
HGRHTzk1FGJSvuJ3yScesCF5Og62UfF+2WgarZdGdD6j5b653LkE8scoGBoPIzDZ7KzunQ7tYr7+
E2LXsRYqQQ009ZVCspNLSJawheby9rlsc/bvauQ9hlQUDoSdqqUGe0E3yD7Y9O9+VpqGweIm3FAT
kg3zdZt8qsy5sFqyj9w+IPlIsx0OysTw0moWNwNqyvt2bOK1rUUqpNunnpZfT7tpjFqWIUUp/pky
ltyV+G+JyLs/BSnvKRwqssdIW+qroxLyuZ4apRxaYue/xd3im+u30QqIrWV9IY2Nm/xpKNPcuq6d
pGxphUgRgWZuZQBdBOcubWuK+dVTjs5rce8nMorV1rUS0sV+QYhN6yNXkWuU0w5RedPFbjMLKEry
0S6f12zmRukSQlpqkkKteq6MuTdCA+4c0o3bWuZnDEFhVGO6ztFP44MpNjL/UzISrae2DMXO/IFK
/Ny4+3BBCPWjaKicoSf4suNSt8c2jnD8Iwwiy/97kJVjtd3fL+aBYevQSnqZPPcWlK5HYxvZMwsJ
JZshszUU84RyVmX7N8ImF22rGAhI3c89QPshmrJUbDTksyFvgJYNuEfoO1EeKlBYSCUJQAyMmDkz
1++aWtRCR865+xOcH1VUMUi7uHfNSOuwtDan2m+Es39vzKy1/58/oOyAsYcVM0dFYNJQrSuYJb9+
gpCaq4c4piymAulPw2sIvyE54vyhTZx2uOYlLYkUUl8BxsrpSAiFIKzWx+3sKt9E++1sz0TPlFYR
ilZhi3GbWroXIlxN6eqeTi4jilqTRnGuDI4VdOQW96Uytw0PcNdYIGCiTK4kBGcFYEleaD9J2sLD
ALSVcEQqmxlT+OSystDhLAEudDY1HZ1XWaGyRFYpvOLhqWju/mxPLJy03FP9ht561aVUNwSvdV9a
lGpUdTn/V9zW6urrjBmZjxGtAicO8E812CXVHO4XMIhyGtaSGfg7R856cl8a1HCZ5Q3oTt8iu7os
z4jBec10FwCj+ZjGXqWmMdEpsjHSc1997jSTCJIm+v8jOp3eK8y7tILPB25ELa9lbCZQKgekYfp7
Z4A21Eux/wIsrSjaKgcSNbZgzO+yrMn65AdHpgWbAG+M3c6FSOwaCJFitKpzVuFDkPJg+ZBRwzOC
AsHFk1Qj0w220oOoE1AilglznqjLtBPoSJQkNT7mEyLXP/GbSAdk+2+3KaE+StqtOa0T2JLDh+08
Fh5iw9ajYKCaRXdqcCfeO+xpplcpcX3iN1dPu34S81VL/g3cAutWg1ON3LQfTl/qG8yV1acAKNDt
hAsusYObGScBFaEbPzgf6y24Ig93Ch1nDycPe0iL5x+uLlpyamrBi9T5ZP7BMSmiqzadtXS5Ll0k
smLvoRng0UoHDgNzjhWoWra8Iekv3ERUpXbQV0DC1aAA+KvlEm+7mpGtY0JLDsEK6yXmclB4dx2g
Iqy9PX3P3kpkCCa/VFq1DpJQ/TV1ZXZRN8RuGG9TRs9aptPD2TTAPoHl/xuaLQYkr2FmgaJH5FVL
tiXhmAdq6EVPih+h+K8m+Ju2Zhe54+VWnFwuM6zpfXxenuFINKs9yhgCqeIHYea5JXdZR/8A54+P
hTflMtxHRi3Helm45uIUnSfy0khNRGZxMXPpX6nL9qZauvpUT2TRwBqJZe7aEwYBGC0sI38eJ5kp
MM/+P5yLDZS5wtU5vIdQMTbwAGN4etgiRo8/DrXaYlU5dVlt76/Oh7dGr0dpxD1Z8jUG4EsRPJcX
77uknnj1b5Pd58KifaSsZW+OWoiOhJQmgHp0GO1jV5Z0k9B26QS7u0S2P0h4rBRHU5oNQ7dmn/t+
KZHXPkp+kNkHVvxsasSnFZmj15Mc+2UtX+43+t3ogZgUIUrFfioOX4W/+WFJql2aBQjpOutSiI09
R0SjmED+SxTFEl30GE9KPmCBSOUsEGbgWgIUYBhX4DQG/z/YfGDcpWSv4LPjwzyBZhmUxrrP2qee
1EPGL4HDoVis7bKzQYrgvc5sy6bi0Ejs1A6iMAafrrqlXtoLshfPNeVebaa8a6N0OoE01YFknFZZ
kWd6zSTohfjSFo16m1NJyuLpWa/qGDq4DEvroC3YFmW6dnALSesSg5j5Y8rkZ0holEkd9cM5yoh0
O/t+4iCECTbuO3VEhJMzkle7zKsCwkRmxL5xWeYCFbDOipCVHk9ImZsYN2MZ4/2B0VtgTs6IddAI
rNeS1CdFwvBYU2Br0wfMqVKRvGMvfJ8qGHmTqGFoiq0j3ZKhz1wheDVfE0KAFbHO3tTyYMAbvWMx
HkuX1xJCOFrWB52VJ3VsFthJqxvT5630oEq6rs7gOY5C4c59BSLuwAeyB3WTQfcW+BHSQQBZmF14
hx6z4jzfRV++8hUiE0/JERzweuZR7LQdP5QE5LQE+1qG/1xRVhpJlvyhoYJKXiR2cuhczDXzZBM0
QPNz8gMYFSKkJrDg5i88HVAtq5tomv1hHuKLXILUsHsuQqcJRd6Nnx8rx0GfNozdHI/4m+nb21G+
qKPG1IQJe9ArWsmTdaqd37nk6MT9/Q5eSMWEejTn+5S58Fsq6AptyJ1F6eeIuWhdnrZzRB8bYF57
8/hQxQ4Mwh9+Ck3QZMUSRytgedF+tttMS9ZsClP/nFQDNN//M8vm9J0R/q3l++kEHzX4wXkETJwd
i5YSwcJeo7goNly9GyWqRkYdeWn2dBgnqDzv/G/0ODlWlZOPgZMHDoljrJr8ota8BFcmQ7LjmiK9
K4PPQFan1Bzub1tWjJlJCYyJm9+FRyn3aC/JJFDendWSFYl2ibAEy/S/Z4/leFqmSO1vbuu7Te87
TbP0/F9dqCkH3lF5rPcjVGZkhSxldxbjSvujMScuwAUXI+1H4Zkn6X9iWbS5t0PU6UynYS0h/4My
IvfDB1a1e5P9ZHadb/SkiTniaApPRAMBjTwsdVNSU/FQ1zP8/sP63Jb+i/z98PN5hyavOc7oKANz
8pG0WONT0by9kUYyTvd7Av+DPkPFaQtqWxV3cJ+Y6GSU3CAmnoXJrvcBRgmXgeAhtrnh2fXGH6pN
Muj7/ARNiLqI3Tekitz8r1jyS1x5cIf//bSkuoD4S4O6Gu+iCSiRLthG/32izAMJbvxe3X9GfH8Q
JePtKWCweE9zDEV9CfsvvRp+xLbswBWsBorEG0KQhmZ+q5Fvzfi6f1bQCrY8r7SxIMkneuTSbAao
tZLkbsL2aMdz/WOJGCsCF1IypOt9/LWmzKs71yZG0XXBFZsAX5OEcldJwWZhXlR0KIhG2nZKY0eM
H/ee5Cpv0gldeA4+ggLODy0R3facQtQg48TP8VU0nzp2pe0VhlPGTnjdLKKjYcNdC818mA4f2MqJ
gfCrniADCMkyq9i3JLt6GJn6qKz1LxpqWFQsW1uwdqQAa9hiFmFjnQRvg4gLppWoomS4MqPYpnE4
iKNOxZU4ckej9MfrJGneQg5wH84UuE1XOmq/TjItj8bh4y5g81tgUwVuysKYyucRmOVfiD4HJSBN
m/EHMjEhCvOL2ZFC0w5Y+4jNOdJQ6WihlbEwuLa3/AyXjzFJ9HoP8bjfI/G7tk020OsjvVe6tkpI
laVD1YjwSiq80WbZCiDO/g7GRQqau1xsC4oomx42QDCjwdIwyfpQ+I11jhGteXaSVtV7fvOClZQ1
1YkRBN7trNZUIKiF53KsDvpJZqsmHa9tRoTDYoSEuVewprjaI30eaxVdHQBCI28G5FxTP7VFIfK/
Gu2AzPw8KmhJQtKTgar+VVSZesVtQjuGWrwznERNWg01rUR+tgZqXQaNBXkkfUYN4ZbCVvrLBz13
b/FBYf4hqDT6TdmacxozR+7XF0WlrEnRH9tO4pTfiWX9pJyQcy0MPRUpV64dZm31DRvxURSi7bkF
utqsn5sQ00+19J8+Ts99Jek6oaxX235gr2g9sv+RRkh/eoJTkVSXGUKE07rvA9dc35Q4uIJsT0aY
Z80VjHoMXIm4isX5DWPoyTvlB/ppnUtQdenLNnkrkD0Iw6Bk3WjBJuz2FZhuBCNZDcY5ipG64cZf
SVObJNoPItacBp3m0Z8CpFHph/ou7BlHH+1lNUgppcnsM4UVFdevl/a/UsAwyEcBvL4N6fE0BR4R
sAkJy5iUhtasxhJYln3mIHWwxnfdyWDpveUIJWTqCZGm8bDI1FjNms79WFG4/YMu5M3rb/CaoiV3
WYzCkNPIE5ooqOpa2Bl2IcRl80omh7MeymaD0Pej0HXOwzijEITidRazceYyJhPvWCG1rJxn43bS
uGU/nkJKz4gWV3fdljUCa/3j151JTIoxsffRK5KBaJ3mDsNvpCmdw1Z/amdvGX23saj0PhSC3b10
RAmXpsJxD7HhaWozDvUrZw0H5O1Sb57n6dsgYA5StodRbbL4+/jsaMQNBczlVt1DkegVlTOwZB2X
Jujelvw+NAOPnh4dJU74iT/E06cMPlLK8OdNg4RzuQkN22ueX2oXKpfCRJ0jck++hSzegdh2qc6h
jnZ0l4rmPHor0Svwy5arvoTUjTsUuLwBHXw/7/yGm00I6BdV4Hs3FPIxm84sJJOv402M8QYSSyn7
5No/3ZBNxhFKu8lDoLi7kzlk7iOJ5zaPhkurKYE5uIuCgfKndE8UTg2yg30AAbl9nNb7KBW0bk56
r9pzfGQNJI0e0QUYAJOfK63G6rcNncSJMbDXwKR1MZAfsFTba/iwGnBCLirmfCtskQdJBWTFM/ZL
Am20OjaE1w/c6hiuW+eL5Y9opZFmoIhuqTQBMOBL+6zs9S8JUK+9EsjlSJlhkec9FN1qZ1HbiFbf
bW9SffD4qbCpBavn4g48FUPE3Ct9AsZDYt7SQtChVLZGYqXwVzAKbhGVbGqmtLzuf1fG+BtBK790
R7a0RkKiGB1A4ZoY09e0WFhwF59Mfy7+EsYQzKuZ/+/RopXEfkpIKvpiyE4xWvUTRmFeq7Xnhj7L
B8oO1XGNO8DrMRLAF5vHNiLB6y0xteQhu+Bc2//fzSx6duJsErEMumodLFwcy9jfeHLlW4xCuPaV
Uh25QkuVhS4iToar3pxKaCNYzXZOp/cXiY0GL7TiT1XCDx3Wit0PCPibzm4OI/u25xIL2ovKGaA5
Be45ZWxYJ1qOm+k6GDONwLbQI3GzfsyIvi9J9AFVTxU6/9IkgvV9EovFQOeFJRT00cQXyPiHNK7Z
btsDFh46pubkgJ0GZVTZuBCedvLUBDFi30aLXT6KDyErs1CqxkwaRG4bP1iCJm44RFdGZrZTWzxp
6iTHLlQ8/vnEkbzEjeY2SyXzrsPNblbgJ/0E/PVO2EgLW5Qey3BZ+BA3SNc87OngqN2SI0KwlO2X
nmub/+iFhbf1RMn9LtRda4FPLJRkP+Oz4+MSq6x3LQ2J738AG8v5aQ5LwdJFByhHLWuJ+om4/ZtO
647up0WqRkzGvSQEps8vnJ3yjuRLr6qRrEVpbXnY8kSg4HcE7JSSYIBJyrFEQpb3f+YMTV8Lq2/j
e8oxX92tFK5Bv//x6sG92hNZ9KjpXGycS7HxKhd30I+mZ5YkDVdeNBw78n/cMiP1rs4JcflIiryz
T6yJ9pg9g20gkpLplH95MxE/UYPSiFFM0+TSzA8cUiGnMqnccqsCeWUBMFUwMq1aLSBeOFfK+6Oa
G9gOnwDStCtKUKKM+lzclrFt+5+4/nc+uq17K2OnosgOwdICiX8hRFMM26rHH/dS2TH61p6sW0yc
/hE5etDCp1EIXIl5AM0LXQPZZhCC2VIYh8RsYQG59rRpwx5JF8DZFVYdNW9CSF7KzD+OYu9FGfjW
0j7+73vzWbuIaLAunYZ6lN5EXXKN1KKjeO1apynVuVORxWsrHk1cldV0h3e0iQC18MQse1lxoT0c
tB9+HgSderjnKBU6jGTS1831At/mCxuz6z7OdJhMdrLTct158A7QgrgSC3w0Wsi5dLTuQwa/ZRRD
9aqr7hmoujsJkmrviklkBfEVx2tq2BANRRFUH8O68P/9lR7Sbidp58j4uFfcSAAYP1cFTHjE6g5i
9MUMk3qbCTm9kD1GIHrU6MU/JzETWrbbMJLXPQDgZ46r0iSfGlJC+KYGjsZ2Ynr52OfZCMjOiBPw
eqJozDeWph6vToNK77KZG3oZBoXTpTwQe6F3+6/eynLm4LK9ut5RpF4UpAt7U+U9S+fXWQNBm9ZN
seOsJ5Fn+bIhCTJK+ezb1NPzK/h3f3Dk73map3AsU3KxYMqhxHirXJLpZukbofBhbI52bG66+sXE
Eyhfj1LtzVQPwq9lxdj+j7W0JISROnuVWUcjTwLwnUOrfHbZi4dMD0tcLEngsqdW4lOrLqI/3XG9
E5/c0T9wYimRpgzRjKtEBMPxderERG8T/u9gdWuHVkHhXKb5jp4A2zMnhvY0KmqPn80YM4UxlZW0
ewri1RZDmYWsyMGM7tluAfrq06Q07ULGCUqdRZynKZc5eKUwodoZQdQdOSue0MrjSpSzh6M25QnB
yeiA9PBcrMELRYIFzlYWX0MLdzD3RrfavUpD2k2DH/l/hOSE6bQL/pVC79LpWkhegSvOVI95XffA
yCekB7hhWIuqsS2JbnHoHTpT6JIpO3kDJ0PVe+qzMjNCTeqT69a9+weMhwvtBVEpBsOQlQUHpRm9
duxl4q+gRMqhLQMiN7r7rHimhy0n7kffgCriFoYO+IZHBi0gri2fC10oVxhgFN+YgoEEbA2KqEoS
RW3CuAxVi+9pAv5byod7/VaxNCRaBWjFR0zfPoy0/fz66GPjuMnB3ZWmBKLuAfq2IjoGBg166cjb
6FjSatY+hvSV9PB2TNkL6Irl/rtajyrZPPjXVxauH3CGYoMl+AYAsiNk2YKliVSM7XfSrI8zSD12
pII8zudOwFHFBzsy/iq879V2CexGdo5KS1Dh/csmjy8i84FWXM99r/qJ5pGOyC8mgxCY5ToCAAOR
hydMGWTAcTGfFkY63zgc9Cf972HMpz+S/fdvOCjLepMUfR8s0DqhYUh/lshbslyYB/XSPiRMMJ07
8bmOnr2mrxuoVOdKjLI6olrqLx0BZT/QTkUmJS2huWJ9NjAxwgY9fZ9VeidtPZUvWSAjQEWHTXNN
cgNXYq6NDI2IeOmxaE+6Ti7HJZ3X24rUhl+gjrO8IO8IYUt2yttOMl2buGdBek+3ER2XJtE/sYoY
pBEQOXRxWL7ap2si+AJEOGwkJWC235+uSXl3nCs4Yxw/uUFuqssmwqgzKRFUbLDQH/ZnPe1VsnH+
0LItwye2E47cwRrkklvQkbjV7i8Rn8V1XWWolRcnMiGNmuj6Dt7HlTSWH3w/EsvnWRRtv/tCzw7U
CdkYjVvZvObfd+MVD7Q/QGSMNiFYUFgEDUaCEyaj+mhN8aoOuEIG9ZgOAHn3ufqKEgrRS/M48q3C
54Aevkdb+M0iVeDMeTBKReHH6ruRIlgmv+dyadtrNqCYdgeDylwElFc9u7ze2dIFSbkQS9oYdp44
qYvEEENW285bEfbLqfrNqR70dZovUwO2vUhleabIwx15V2WaD3pM6UJ7OdKVhWIQ/uqLB7XyKns1
AXkx7lIXdAvak++e2ZQ5HKLC9XUUyfQBTro/GaiKznDyAoYHbyLTRWz8BiWZSN0xQt6dezP3dM5y
V4n6zOZYHZ5EgxvO6meCigxMsxjWUlGbkg8GaKcRQmD+okm3Lf9595C9AVT6VwtVC18V58xpRKjg
13nnleORS2X0YAA2fj2JF5zMeJQQPRmy12AsOPU9qnjoE1rQYZriS4QKA8PdeBKClzIPxfAvmPgy
hyR/R+aAGb9EsPCMVD2EfvNHvLvi++CdC1zmKH4HFxWVO08XYfqzZyWOmOKuC4u1ZxyFIkfOUFVM
euJHO2SU9hFRuIJMU/4f4P6djrmIANO6K/A26vvPrmMrK/k5FX6jVvjNT1lRysjDhWqqPJTKL/DS
xxdRtLpvqQO2TKPV8cVdScIdSCVybkhpl65PXQch7RWudaIWj1Ir6k9Me+2Ci6fMijy+NrtTF8kv
7xOF4FO1/8qW2PjBUikzB9hCyNA9WsniLSpX17ZGacpshZDxZv81ImJozMsh9hPY8pAqavjL7iv0
ssz6awBaPSY44KKWxjZsVaL7QynGai6FN3k/NJO2I29iz1FCX3D75z6e9IHFyEEm6UvFM57rnSIT
+yjNhg2Nr5SEdZdIDNV/pgUbqhfgXRkLTokeN7j6iQeoeNsfsTQzYf06iJex+xN6P65h5eDnaYyU
JUdQv0IjuYwDtLJpGAM5NgJoSIlP7kxS3nQDPINDsJdrcB9FITmRYxVvwXYxS+V7H81lIIEkNEhT
bN3TX7rhKZJDuPhJ5E8WyjyMTQfGkOMFA6eWfQctXQAVhqRpQ9HQSXzf4Ymc1mS/dCVYfvjhp8tS
r+TWzpVg1OX2OomUpiC0tumhhYQFiFnwD1qlwUkXsljyyPUhNUXAVDC6gU6rW+SaI7fjF/kcmCTO
gaGNJp4+4URMFzKT2rQkTaYg1CiHy8pus1arhf7Lw7x4A7kU3r8uTgmnPRMF4P05FKPDvswiZTqh
Xg125lJLYU1POUj5r2+ly1TZAm8CPcGv07GnaZKofo+RItKYIgMj/o/Mf3vg+CUtuCvrcXC6+q+g
tjhWGi4GTKVovJRdjZGQcIKbSEHPrDMP9YZougcTknz43IPttnis1W6pNNsWa/3Pc5A/G6y+cf0X
dAowYGKKUvvZJDNgNZiZWDpoIjG3xKqCKJwP5dZ8RA4opdzfY1NMWmCj00j6gCroI64O0KHfjwTB
PdpKnAUImAZnHxggum6FsABk8/CzsO5iGWM0sbDI53xlhB1p5OX2IE857Etzk2n8f3B99PBnbmVx
Pok05iGsvsgZOXqbFppWSYlxW5i0gGKcRmHuEgqd53qC5Fs6wDkYODufV9gP1Ntb1gomAflkTRxL
KpbaPmGGEv93R9Jj12EWRkJZiXdymkJH7CmVJz94FOzTdEyMTTfrXiY2pEYwX0LImCjSVyIaxjuh
3Y8JIc7qi8SN4dDsZh76dAHHZ3XlMmbF5mJY/SP4GmB+bs/+xOf7mWtXtTH2X0e0igFcg9u7Q4PO
eKqN1vQIrNYoX8Wtx5piYBdypBGJ1nJ4zNPhArPTLNosmMEBCFFm0MbhKIeTN2XMhvyElplnKc+d
hjFSSDIh3tTvWXAyaFYlFvNBQ59BKaiTHMtbsA+52QcuiDtrOST+V/NL0xo1VDrFKuG2ZbDX2Xsn
eFsfNiUj6hdFVo/1Ap58uboR1c4g3SePCrdcsszXLySKYsr82MM2OyV0pVzr2U5pruBarRvVEe3/
QVqx1YdUg7zOpuh2Iti9jyPob8Ho6MIauDs1lBKO7uPyDXKLW9piby6EFzJTU9ivTLiNRzBJBZM2
rj6ID8SGvcvCA8MSbUIwvGRGJT3k5c0vw+nyxU4/kvrNnDpalTrZwO3uQLE+zPiMy3OYvkVscPXT
WeBItvz7N7oIllhRTmnNW5X9hV+z69jHx0pWXVbVqj+V/CeUjkqU+7XO8P9YA/oeA10wc1fgTTAS
04zFuze0L25kgW832SMfwdmwdOYW6kS5CUDvdGTHpUIgF5jycE4dSA/E0d6MTsC19oedM2SZkbcm
LN6PmIMNDJLGpsDeNbtHu1lat8pMxhQOxusfHKG8oHNJChcxRUkYR4maOJOPOo5BLbLazAQjRxX/
UDXPur9ZgpS7aO3L2D4k1Fqp6M2xJ7TikKb9BJYZGasmS5w/aqQkm10zAEyW66qY8ud6JO49NYbN
PKgr5myWE3WzhT7wG4Zd2uX+UEA8wLBB1vSZNI4oWA71jDKw3Z6fBd5hXTdfHK97nBQZh4M846h0
bSttTQJFOz4osyVjodSGzRD6q1ZU2wanuAz4lI3tDbfJQxgDhPNmcOUxfLJ1Uc8oXEhJBrXHk89C
f9wA975ylvNi8iKWEMojztE7XckoptDjvUWJKe8P1jHy/h+k/DPnsw/MHv5rfqdCtab2vYrvVC+H
kD47MgscnMZ+vZWBGYUFb6kKF8TVLbIK7VyQFBukEyvp3Bq++joiivrXpl5r0UAr3QtIx+gWYdqt
z1xKt4dF9vUnGGI8bGfhdWu/GdvHkE8gnd+PhtMWb0rOz4uALkv9LERA9+hg2DnUG7j3D9zB5HCd
GZrO9TFj8MDbbyIz9xSDx7MJUQbcOWWCrTRbYcm3KWj/YDfTlkxl2YjZ4rPX7MsbSUqQmTls282k
4jrylsgYSMKjqUvO8rH2/ivBZ1H6y/SXHX1vXRJYixb2dWka1Vk4CZrze82SCCz2qtEhn57P35mM
JgPDthJIOJasfe6pctLW/TySzoNTRwzTYuPzV54mlY3jWDQRSGjoMFz8/BmgxsRG/I1H2GBga6/A
d4/TR0ePivkXoQI2eU3z5+MJBvIfTFl2eXjVlpVpMXq2DN1cRlMASauYVrmM2eHKf/V67QBsf8sZ
Eio8QWNfg+7D4FnuM9lCkhvQt/6I/74S0FD+Vzdm8mzHsfRWUfTMvgmUmdSikc2OLDM4Xuk25D56
3WLUO8VEErLnaGZWE5vEWxIE5YJJ2eeIaZG++9EuWnkZI6DfLZEkE6wKmTeCmROBwG+XgmXcyCFq
x4HAKCoL2SD1K6eVqVwXD06b3z5vC0iCBzxEPoLnLcUqkPfghj3FDgu1hDAqwkp1rNHgq7/sgCpf
g+k0O5kDcMiak3KmNkD2e5wSGCOJ5myYyUVbGZ4+pBQB8fkIknFBy+pmrxrl15uqVVGZjFT4LUg5
9KWm+ShPfWJRLwGu/C2KAxMGqEJyjMi/7GAKaDdDeB5+YAvbu2Evihe+mL+u1Liji/L5Oz9VRAP+
b0H4WdZfWllrEcoWEji4gn0IssEKK1kXH0XAa8Uh3feGAlEp//izTjzlGBPgJdvzoPY7TFj/9NlM
SfGuh6oNhzkj1L+XM9C/By75UUs8qeie17FWCfH7dNeV24IZDjVnmBztqN0DrHTYUZLhmrzoKXCn
6RqOZKvQT23UBqC1tM16SEwugH4TdJ2W/J9rcrJAPzsT0l6WC2XCLMxPJNR708zzfkyW/kP/HLtk
OJkZIQJaoBu6mdkmHWqqKIpqeMUVT2//kizNj/PcTjx3sb1iVOda2E1KkaVOItqrrNfbn2kmyxPu
YHwiTT3ja6RkMCR49TTeWsvbAEckPpNhn4QIqbV8y164chmgRXt8UNHQ3GgM4bbdue1jh48kfzmT
qwjN8awaWFLy4j83BoS9vwAPNnb3PQ5GwFgd4v3N5zFFIu3FAQG9qTIKk83zntRlUi5BdfClH0ih
5kqWwTP2eT4QAYPO2F1MkxmUA4uC+9InY/vuQ+HYOp5kM30hvVgVcU3wiurL+mR18DB9C1KQfQOZ
vBGGLyKzZhgfjwDrL7AnpMltUJ+xW1fbhgm9Z6lMis2aVg3cKlM2rpsBX/J2hqXfzQaVDO52fvsW
fmFZmqZWBkhNVgAt637PhnmqGOgZWo3FyxFxslR1d9AVFhz+PBcA8DXIeej7zFX+asj7F5C1m5Vz
g4eGombNwGMd0mzFs706zP1Opt8ROXJSD8HIv7FoXDlsXLEtpG049Jzs3AYgFTioElqcaPSRi1v6
MgpkK4nApe4Q/KpCwib4VAhiPEFiskL3quM+jQFeIW+d32dinpgeLFv6qK6ZZW1AmYV6nssvSQti
8RcVc269/N2tHTA0W0B5E6qKI+ojYC0f9EXI6ihNJjGCSl/35zyLlyT+010GB5GNLDORRiFQHTNk
rYObnqrSQnv+bTuulXkwTCR9Kke+jzZcUD5b6VFZbYfSUX2BM/zjv5jjD5eqOjnlTwVg8cc6LXwy
/+mJ5FH6utV8FMPabdd3mpNrsCq5JdDpAxPY/NJqsFJWn2ewoAIwORkseoct561X2bpf0FPFhzGL
43Uq8EOaGgCEG1vvfG3Tu0IVz7tfCEYmi5Wf3k0KO4IGipDIzDuk0KphIc9WjHQYsMF4WrTaJLe/
VvG2nQ3DrWWp1Uu48g5x+bUO6AxMLdMO9eL05YNOwVI0y87LndmeKoi/8sfK0rWswVWoboEzIa9f
qjczHU/xiAcrv8Yf80l9EJyMX3B32b0S1nzbPT+jHIAOtV9OHRMlD2TYKWf+PDcFsVMWjUk4wvcx
Q3pMgMZr0p7OSqqAyl7x1tTKs/WS3Re4AD/1CsKQjRrDAqXw0wTZBbK7oefmScQtulvby+0x/OQf
rbBvNW7QcYxcPXT/Z+/kF2RvUAs9+hUKFTHjxWC29Ojtrlyfi9lVRbqfbXGJ01F13U1f08BOoiST
vXfPv9ME18ctKOu5LpQrip+bVgfMm21UrUaN7SP0vgmG0l9U6TdNMkOSWQareIS6PVbmssBgRvs/
eqpiP9mLos+9gWmazEf6z0TJfts88A0clt3cvSUqafXFSwBzPB0RiWloEpzGqFoeXZqtIN7BuxMj
pu+pC37OlCTyRBIpZ4rBHhpcIyV17LCowGFfqLNvpowxTIPHFHRi8h8euwb1yg1s581D5MO0wvOA
tiD8UigsoVOBQmmz/YvwikGeR1AfDlB5s0jQohz+irm3Kr5v4tXlYZIrQiOEqViBJYGGt5PmztAS
yGNEYEW5DCbTX5XKBYD+XrA7Q/UeTomyNJ9epAOGIx5WkJRl7U1ge6XkiHpGDzZQtShphgbSpQ9H
rxG98zx8TtGTU78u70C8/xerqGp7fCNfJFejPzxPO7/liwQ11DnOEw+oS/vDartBW9H4z2CJV1qw
/3U+6W1FRvqXtxRi9HOAvHNjPwl3j7sb8yV3EzvR3NjuwjqLn3p0vHHRbHZ4CN5vPlDJnJj472vV
mfu/1g0JaR+Mcm9w7rlrjYMEWExJLhn492KWBoUivjhmIbokAOy5WlWAgm3Aa+FI1M7mxNE66sep
F1BLnzzhMqlrLIyy+iI6SsUPvyzbOigk5f4bTRyqvD2dPLUSwV7u+eJo5wOll6YvqqszWkcsdF7T
7YI6pj0ngkoeYBWfbs+7qkjDu9X1SmrDXfTnnQ/DLLlBaUZjpTvakE7fRIYPgDxUgXk9WuUVGA7Y
fsUngK6mk4qzZ35/SNpWr6yizb/X671AATgPMs7iBYYsxJYFjp2cxDOnHhHqTAb/u6po0lPsknr+
2AYGniDDigLNhTEo8rtY/H3d5QNKoVOs1GRjDwY8/xzXPRYtB/yMxIb6yKkCBY0Lef7JKM8CDzCD
K5Sd3wenxQbN3mY6JJtQgkuz/F901lqKxbWE5X/cCyirSqpv3xem7JooBYAPjaR/Mmj3tQr3CghR
Kg/kbHKCKJAA0k7I9NnHieLeMVf98kVf8i9OSu+nLT/UidgnehdOeEWnIQyrmzZqnZiE8M86uSgE
OzdcR1KfsDqZo1q7CtWikK71wO3Ry4TzD0lPBrN+HNAczNo+63bGAX4C0BjK3DQ/EezrdAyFbvfU
OpQQoyiAzJCS/rinAdoBuom7bNJi1Z62yPWCCD94ssb5M3hdigCxMbgn/vO3lc56rdDaoKIznZgA
6d/gz/PbNot5bHvP75B5fTpGZA/q2XUrF6GJacUm06swOsssWYGAYI3jnIIRWwmxL+Ytout3Hv8p
6Za2sDQYS0dCdZ3j0FZy9fLR/Rfj1uXti74SDCgr8vCpNNIv9r6pgNP0MHMeq77Ve20jUnl5ZZtu
ajcAydp5X2pCfjcV2JxvKCDsjoWJuAI2Sh/p4eWa+j/pz8+oora6gzCf/gLlNNELOCJtmQVvgZfo
+TaIqzppoJga/0iUOfqnXoiuFg8+YbTyC6/MiHhsceW/erG+Zn8IBSb0luYs3CkKHeqW6TA/OS8q
4tOijTB5H5q4IOooC8eMuAWo/AdFE0NOSi7Xv6A5yG7KbxkIS9dFcaPJ/X31mo9ux7wRBLmscjEq
YXyl6S+WbkV3FKiK+P/qvR1AKjEv2WzICrc02PfdLeqMCiaQyctkqf6aiRIXcfIDpLM+WuJZ/6Qo
0ksfGXmXlerJecfAmHltaX7UnQgXBtlOCf6ku7IdzFn5tGU0ka1HqFhpk1Mab4qIcs0KzDX2mD5F
EG9MZbmPCSE9+ZALPtPxRKBBIWYArT5+RWQB8FBHTdGRPYn/bONQSr4vgqnrmMAlhggpfFcG5OE6
K6Ek5puKw8YeSoiyldIlxoTa5hDBS/8wVeMZSg+52f71/9/3UEFnG/xZQL5Bz/b6+jVJJzicTeyD
jOw/Cu4vVRC/FCWcWM8pPZo6cqIckeJ+iB++fQArqPJsxsZuVGTDK5jnTQv291Bzno880YCpYr0/
XLnjVKmfhbQoQ4kWbHPKEA1y49B6A5mmqKUXEOzZd1ZdeNcBW2rfL/RiplJKNHMAxo7C+hmr+ftV
lliX3NFEZqkhl7Lk6BP0pFciBBYjfADwnDz0nWPN7+zbsm+inAPF+4rr5PTMOFekNtAAENQne+G4
lVbQqmDDrdUOs1JwI1nliV/VzhZ1IFVL6Jh1csLF8r588CAYUczZUymaMxp/my27YAql0BfnTzLG
EZ4/1lkZuvnluPreCCIPNGYn2QlJbEhzgL9ZAK0KbGyBkac3ezoAm95oZBghO4w93e+ZjzNVYzx1
uanomeM8kjq9Br+yL6ywrqGL2YEOjwQ5MegoibHgnu07NMtiM2fLn7Bb4G6aHMet6gGj6eT5vFjn
65JgF2a0Fohtpmews7vdmg/vB+7HCvto4hZlWZfzfzGsg8owj9FqAvOKX+HNyZfuMG30ZhxaHPMw
saqBJ3PoBV0Psqi73Uw5MEKXuzGhYuYubZKrc8ICP3u4/mLeezRrGK6/2DPb/ZlJFcSvEjjNpHlN
85llC8j000eMPb0jQosQG/3bju41V4O1GYq4kR4/jTw4rs9STRcu14QXVy+n5uia8m1u7cCCTlRu
SdUkxum0VLjeJUrXWwNQPdb44ZShKobWsOgv/OMUfUO+uyrxQZeIptDp3JW4L5J7xMm2OirypRAu
em4hBR7EmfL8gbrKZuF6E6ceDAnrJSsTFJGSyq4eeJHeAA3zJ0TlXT1IGA9wzajN2iLTmdhd2LU6
EVveK/MGF8Q15c+inoaAUvlOSQ7ZgM7iaYWI9uXl466D+uKRU1SCP2U+yrt9z+4JGHZUGRDXpFZg
wEzoE1S3QOtIELNxznCsf3VzJkg129rLVOQ59nuavdOpcsI3QUl5FFOeNmNPd75Vz0OMJwdUFiOa
I8fXriYgkIuxY0brI7HpHi8lDst3pNxQqo3i8fQoqsettjDmERy4ewXuCpQePCZaJyUOpB1Gmtnk
LhtAs9QkC7jBt9Dzt0i1RIyupfk8mkIC+ov4ySIgx87asQ4TQlS7tLBTr+2OIAopiYBykx1/HIJ9
gyxTBkWdMvzg5FGos8rzP8WHTf2jmV1Cb29OUBtjsJZw0LR8CFPhJuiMI3c9X6G5Filt2mKHJLz7
V+2sXVa6PoppJHPjwpxmYEBe+YWxUqiJASPpgC2ItlUIii+emmW6e6IjfqplHae4xNRVUMpe2HEm
0Pj9AeC2k8XjLye0WTuZcUzJpQvkXDXRGy6Wr/BL6Yt6WzQizDpFAGDhALOFtf/Z2E+PUu1G9ItW
2t15I6R0LlTjoibOqB+Y4Qc131M7K9z0kidX2gRMIYInV+A43zj33nIy/tnJG+9nnSUXIeRvbw3r
WF0WQaLxTWeH/1smmcSt2JIsPzzUZPxZpRuINfqw8+eLY1Az0H+Ga8tDvvzCUVZiaAQg8NbOeu0e
Wo1PyeB9LG7ukJtqfdSq7b4Pylp1pBIDaulELmaisszZnZX1csbOVTxUiHbsyZgYkIHm49DxJyxW
p09oyJwX4XwUG5Os1JjJmPvStF+EWohcBnBpyjAAA1UzBlLwbHmQ7to9sXb5AoNyxGgJj6AXnn/O
KWLrbd9tQpPGPlmfPblZ9mn8TREUz1RPAW4a4BsKIgdf5GQga3GRJEeJD6EE9FvI9CFf6sGvw7oT
34PQ2AM/Cac1TltNz0FB90yImCXqD97BDfU8rrUkD7ER3icqPWsTiImjX0mMfjY6VLAHfBgPCyLR
HFcCCSqq+I5Kv7AY8txN4KNF6DnSUTFiwD72E6ijS3gFUX15wHhe+IsgWl+cQre51Y614ZyOx4hb
yhYLfvekSs+quhMhpXD9rMDZ+ZEyg3ylVXwqKU+rZ9eSZFQ1cuo0RB+MkHT6V0txQdFoK5kIp/PS
pc6UFrE3ea2b4COcQmm9/fHygxFVa/on2szffkgYUZQ/uuprms+2RNyXfyubyEokt+CgKTezG2KH
NIQavJjacH+tq4pqLK1przjvFQlGzbVg9TWe4jjxYC+k3DuzIrt+Nv96S+pVMDu17F3Q0mp5TKjT
JlosOswLBtrqi+YgUTrHNxhW4yWS/LUOzLQW5jUbsDIxDQFMCzJ65Yiq3Eq874pHcEB+6D/5UFFu
XZtC3mAukUmJmxM7pSEJnQY+te8WtpjCmAOhYcfExzdc9sYNG4rMLC0I+Rk3ngZ5N9NFPpZFscwX
xKFqyYVXqOshIGevArwS82doXduW5OpOYud22APKt+BslDH544meWC4AAzyEaqICkm/RKneAvhbE
z3flBTvT8TdQRrfNL8HPKosOMq9ento55ybQO9ey+yDeWtBEqo39WKQ1mbEevj93aJQ0DlHlbvpD
WxGbqRvP/FCrJiX60zwcQ1goaHv/eVTPF3T4Bc1v/4Tc9rq1uNp16hPTbzaVT+LMOLTLm0Vo7zsk
vVI5CYdWnLAw5I1SCoaeKafZrc7hrSI9bZ6z6um3SfCPjTWkqJHc+nJf49wr6csZELjlSLPiPBrJ
V7BFH89XGG7+BNEpH/48h5NEnrlh7FirZcUXWOPuWgB+MCYlRKFQaelIwI0LYOsh8t2ODUugfckJ
NvwaKB75Kq8yb6PuNW8y+WmmOsSbY61Ajn/AqMWBqSQ/eWgR+gbw6cpP9EodMcI9bN7o2pfKUB4v
9rn0H6GGH1QUqIGbZita0zB/QB9l8BeZQ7gELnWmBTkncnIN8lQlNph8NPEes4Wt+8IgryfBDKKh
VN4Ku3WN+wZD2oNzlUNt2w3MA0BAMLC6MkWtLdxAeRMQkZ8lYugvn8UkYmgUEl9Csgdrn0T3PgMb
HfzMZuH+e63sHPDMXKgzXT+I1tR/XnG23EM2qR003aVnnAvBmzL1qXcXYNkDsFKeytj8EdrC61x5
UCtsPypxGS10Ie5iW9id92n5h28AGbP0Hi9e8MderIDwLYpuuIlleEfgGm1WE4alV/WKsJhxtq1K
QYUb71N8QdYU5vVN7kgVafVPaJzphbOEVKKTDOFsCUsqIs5cEZDEkGcMlVOOlIJ9QBbxJqMJxjY2
Asm9Q437Apu11esQ7Mxh0alpp3ENDEdpoD9XFqfjqi7GX0GJwRnoXVqYmzBOBN7n5o2hyxkrV6Kp
d51hMNccj+hC4jD/alf0J4QUK62XQWGOURhwj0hXYqiYwSnmHAQspmNkbfU/MCIOyvYs9U9K6XHZ
XkEjGc7+HiHcPnCHyaB/eS6g4XW2S0ebdbZsFuS+Tr9YUdu/sJ14T2ynq21/erS6xKJR5Sx5fGBI
P8U5XE4EQ8MjAi7CG6sdf6d3mAxPDD9I28S2t8KkBEyMUIIqfp7Fyblf/HoE+TgsWVdpE15/GPwx
Ml/clbXTxpsmmIY179BhL/OTW9lyYAOCmWWLPMGYTWD/YJCLZxGpW3HSuRADuoRFZcR72LobCdnA
TS+AuBtnqZ5XSXISr8UIHm2BT35zRkWmP1fKkN1nkowC8nALLU4z346WllNGaZxZHGg8CkBCo3jC
/Ztu0hY6xxk4hcVXEwtLIsw67GOtLzvYT8kKBUKaidRvA14tDQdkR1qqsJkqPTJVTY5I0Wvkgz41
iYN5R/kdh0sOKdAxKTlfelJW65R3tyyMpG3BD05v6Xm9pazyMbrni77KSMO1pmVthHy8OvuVb7di
scKa8u3DDTXkml9I7rCrujaM9IFhOXemIpPcgJ5acl90QXk/X5K4hOEAhWjuOX0Ga7dAj67BrAoa
JeKd7axj+MWrg/s8+P5FLmeMWjFZ8p4CcWaeRarIcHB6EOXHA2HDEry+Aug9BGA9/rjB2NwgDVeU
S4SLfU+u9dH8bFSighHMf1DD94Hv38FY1h6PKbyQOJBMDDVPma2HDv0dicJ/0fCbCrtSP179ZEbz
YYkBJ8Cr9o59gTo3ZnvLwLbrbSDyD3judEAnFVCeM+ZwMZn3KEQGlzY6lMKx6+ESDNoHHI8LnmDF
hR9gY9AbdSQQ1fmuZdI0h3iJ66rEV25qQeYxYRuZ6RdG/Tx+3KY/zw5FoIYRZncIxT8L3q8u5D7+
EJTPpK/1vt2llSntudHvlVxs5UTYcHS9EYbmnSZHLHJjjcuABM0K88X4adIACSAutn35FBpfNaP7
hlgt8VDpAWEHuX4MSajYVH19WRyhZNCrbezo1hpZ8rKHAmOy7Yx6/LeLT48txd0wC11p0w+zehXN
p7P2fGLIf47GVcE+ffsO+FIaSkfyZxwliF3qrASJYONw2v+iG6kX70S0TH4mY7qS4Z1lAhCNez1W
QD8dHA9be35G8AgOer5MOHmGP0cHjB8wHt2IJCZ/SPPtumwjNZjwNC+Vavzcp4huwCxD+psGVi7c
/624jEFSIhm1zJA817XL2RHA4AOo3xZ0G+34g3rQh5m4OGxWSymAvSUFRSBtnrjaQ8rche9c0rIA
GegKtLYjgxTrZ272nKWbbpLdOCEPwwtAUdzMEYtksXFmeLjkYR9JS3S0F33XV4vDcGI4e/QzS5+4
VfVm3qsYdY8KT6Uwhezel/o1DOlZ7uxTOGi0q++0FyMgPAOdNoMgtgpSSJw0xXchMGX6V8Oy+6fH
s24hgQOAkI+1t1upgx1ojCUVX7aOggrHa6oLbMbdj6LdoH8pGzIf5mndhJhOVZZvkcjcydXKJmY0
PDsXYc8maPAdw8DnR6zkbEvp5TG/UMjfgpJgOx+SbpbEl3tpJhyDrQcovDIgQt4Uk0Q54EXwtLeD
vw6hjqS2/yOKxGlO1XayzNxmKjQc9fGTY/T2mBSWJDYZfTmY8TPMYnHbh0lIAsOE+NT2kGZZDbQ6
MRtGALn8lvm4wPDaxyAG135/LmNTisb2oULjVEx0r78gafei6EJefIuO3cEgD4lJ94ol/9W3898c
pi97s5jj73IgcuULztQbZQTf3fj89YaApGaJkj2TovtwEOYFUgEjZtW12GxS5PF9YbB2+UrfRfDJ
jm2fNA9jxHDeueoBOI9LpvVGuPpy/A0e3oHNVpaNVOvLJFmNLPmfdd+nBEMhwPOR5H9clBiunr7U
OOzMeJIVRx9Nt8Rtl+DGNRnUzJKkZqmhudg7bbISMozSvnQ3PtSDpM2CN19NXyvNhEJnITyxHBUg
6rYPmfrCqF7t8OZ3W6oEYmNg1Stpxn53vppbxB1iHFowKH2A8d/jq84Kreu8Dx/qqEnVFsHm6ma4
5Qp9B+IWRaw2jXk5OxuEO4N2/oFu/yYrLse0Jm+w1i1lJmneplO/E5wA28ZqgJYhP40qPd3Dh1yc
13AJQc+KixQNEdHmlxippa9lYohxr1KXXe+pEk+UGmd/2Kw4LnDX6BPq/ayaT3xVD6r999c5AlGK
JLkB4xWkta0Wma+JnXCiNLTPG/Coc/ieSxhontEInKRnWXh1iHsaMQBlZ5FCiuvHHRH3zqEnQYnl
XHRTVyrDuRHZlAZX+qQvgyOVYhn0iOkghTTWsXCNA8C1WQUF5vs3AWxfrYlLHjK3Lkl3DV7SqIxv
SUS3Pq1vt91vKw4ujHTex7fBcQrYg6oOlmrZPt7dwJn4eTpBXjonWNTiiPpi6VocnVhGfVLn4EvV
/RrmgonjXJUE2YwsPrG2AFQpREXf6h5yuqWm/uf1FudULC3b1zSr8j3M7dljZd/AEm4Tnc7Gwwyi
kcGWFITGeUv6qPZUzRgfBI5EAdUvdMYWZVcamNlHqVENB8RWYqo+BxZSK+rz6wm6Y81wau1ENJr9
kdigdTaVj6USA2ikwuLr4n/Bax3QjizvFtKD53lDCxEWNnFZ+Z7HYyhO1bGUF/tY98Y7p3iDt41F
DQ+H1lMNBrLcsKOm24DqlPTaB+J5WXapChgA56SzI3RxJDtjPSurZ6WaYFHDDho1UX4Qd/U5ixxg
8PCbhlhN54c6gz265w7uoTlsqyib68OzD9InLuKLbtdKngfFKr3YEThcoTFBNhKh4smYgsvOQ0fH
m7+aw8c5DGbENSlnRF0S0F/aIc6g48UGglABoE9BQXpeXs+PnL2X9dV9sr3PE6sMXnb4TrcMpn6V
lgtxX0XWASnLzcT7GbvtNLSFqk+1ayqCTK3Fmq40fd4cVskuWg5wCf/do0EOw+0GZlNW8eD2Nn8y
iUtX0Y1BJrbj5lEpLrLK6oRqKnc+9bohE5C5ZX43RVvCm2HApQUWGYHeS69w47daL16p+7Nz6I1v
YgCU4NjeEUFbL0vqKGmGlL7XPvcUDIrrQRb4k49hCCJ6RhQ6sjueM6xTENb1UTnGaiXZllfbOt2x
BBRCsIMyWwjukfLRUIQktXM6gCUC4yEXW2ULXGApzhM6AvFek1dIR85ss+LHShGHxcVywaMpPIg4
A18ft302T9vGYsC+itWPC1OPer4zycExHPu/KUh9mGEoJdM07aHuqlGHyUfTiDvZNVf0KFKqNOuf
BKm6DzV0df2JY4c4WsawPJ+kG3Rze3IJhA3Te4IdZt4I1X2PAbS2s2tYWutHvlW7VsUTcQn84lLD
tAnyNtSx6I3mbwW/ry6V5YcV3XG8RnaV4vIkQ9mvt4scBh5pQzggznEzxn1MhKm8Bq/bvsqZFveU
g1jjc+7LGwhqUJ1av0lfrY8zRJJ29NDdvHlIacNEHR7HD9241UPgUBrKkXIWx5a4m2AtAhQ1Z9Vj
DHQLaeJuDSWvlarcXvU+m0FSxcv6meGq9t6trvjhB5ubEqNVdrNPTTDxrnvOOF55AwNGVuACIX2I
mZph5svsUBlcm2pdMH1oQxzD4cd/fva34/ccdtan72yB04VNL62Isj0d7n+6uP619FqjfE+v1Xb3
8WYz4BGetTiV7g6bqZjBcaiXCO0qKvlrk7fcmhU2RHMsFOOB6+89Wy9iw2IZDcmr25VSxwmgeffH
jiNo0TpCLXkuxWid4ZHrcEHtfEMQDn7uum0y1mytAOKbtIKKqP0UYNvsMzG4xqdcd6NN8T1dxUGD
ViHtYAH+irjFFR8bm5pdyPaAF05WFP8pgSADih7UlYMV2h5zwF5zbYidh91LrM5xMeb07HDkQNFV
IUSvSoPSNR8CFxuMw8UobuGs2xd/PZw7YbwCwoyj+ZCIqPisw5rAM/K/pfOFVOgtAlhaSIk0lA+R
8xbOW4sIbvkaYhXZIeuggpGxPQXbI4y0mS7IeKA0spzZmS8edDblPKuSHGsm48KjVMCxLTdNc8dz
t3MMi6FW+Z4zmEByIBnYzQr75WEsP/DbKWeX93x2LsbYigK0wBRBK58UsBS73SQZaqnT5rS+Wn01
sJ8WzQSZ9qZixCi0Z85WuXOPnHrBxGNgdnjp5PB+u6oSqUsd0X6bqQcIWbcZTHaFuMJDjYMlSf2U
hFwTCROPIkQTcagZTEAA3wyTSx7+qm0zQUUz1Q+6RQ/ar4cPNR0uTgUJ5VAntxG+6o8mXW3Plsa5
LZ5rAZNPM82feebnTWLk17ELe4Zba5jKv95QKkAS+OGa4UH6q9kV+Ykb9N2b2dLAAIr+h09+wYaX
Ayqvm2W8OHqbq46c7MR55/cuZ+WF8uDlwyZz+C8Q5jKtoDauxw/LQDxxkUgYXl/YfxMmw7QFU4b0
2+n4/Dh3Ls9o6IWwhhKw2+yV7KpWQvFXX3g6Kpp0++yw9WNtiK+DmZwpv/JC6BG6kccYc9XK9s7o
tTFTx4++rO2wrAQhIQdAd/uvEaE//tOQfyLM6eDZzOFiows2/h40HWyeK+IqoglbzFqTw/yzUVTh
RFo1EOF8Q8fTE23ikWOkvwBJpLJel9Ac1eNYPrXEB3okz8czEGH/HrJWhqwwA37zxSl4UTKSWk1l
OD1GCKUm6JBZVS0IzsKxCSghIt475djHmbalFmzmb9UJ38/I0CMFhHRbjW7fLn97lG0VHb6PMCGA
mcRezKqdor03JT39KJ+uvVmNIb9UrglwjhhUOh7J17fOFyyZM+2Dhkkuo6EI9LALQyODrqZQPEM7
zb1zI5W5xUWFRyuAcNm1xSPRq3BtLueqpICMMrgsm7QCgaqLnIT+bH3kEysNgLSpLaLefxQD2jZN
RT5R/ntWRoC6W4t76KXVLFuDBspHMVvH4jynMnu9/UaDVANQhqBe7S0g9afrTtTK3EresW74LChA
wNar1bvDbQScm19D7FJDfJoiS4WyMLtHod0cGYfHI7qwfLxbOrQQGWxHrdXyzvHRWmGkTdafumw4
TqmPuPTNCdS2oQg98Holv/GXDsS5cyOTSFEgot6L9c//zPsBuoj8seH+PDal88fWD/6VwbozBrnp
izTFjRWCMEAE+k1E4dox783Zg+fbsNUX05qLGh77NQ/SthioJ1m08XPzfNJ8w7LRZd0edb5KQTnY
uJD1GRLY8rsS29ahRYz7KBBPj2B81C46CKuBr3LOGELS1+jAzP7JWQft7zBpyvY9mgSGDkh9l1Zn
n6IcHEvFtIopJBtVolueERGG7Cjk856q+b52d2zIbGxJ72oK53nMyDXRT8WvpfXFX6TgT3YZJwx1
KbxoW++77MxnOGdnS9qBU4gpLy632BKpQwbWEFtHifZHMTWotSbYP3bB/REdFEs4wuri38vlxhXu
0WjrIOi2Y4WMZ75QhiqjmGe2IelWh2JebPdojSVaor7AWc5dHMb+jJeob9y420qAfg6fGWtc7CuD
eV0GvrejIWEkU1VJwm5UamhtT8Ff88HfaHuw+Npcdf+NJduI8d+po3ADLOn2CUQiaN6JmES5XDjh
eHEl7Yv03EDCsOZh8iyU42Q+AB3W1gNsV8Y8s0guM7pkg+FBdH9na4b03f31HlilqfoPybPlyFEG
+ZBiMAgXtJ7/55y1QCoBifTlvfwZ8kkxUsq+SQ/BfTNOTZx8S62C3qAyAaEF8vwBwze1W/lfh5OF
r4JN6IqDtVm2Rzlc2OaB2LrQM2K3UgHeGzrT9KM1ieIJuWFOcf1L9wTSqL1XtfUsenVnFT5900xq
PJPktEqu3JlLihF2cCPVyHjHM4EdoUYlfdD/dGUfF7Vc4iPVMIi5PFYzx0EcfMTl+jlZnC3BbKqb
H6TAzF4kjeEwqGLBCxoLrIukHHQx38f+Kb38dCzZXcSzJ6J4ZQd0Rw/1cjV6g/xq0DZr0J/i8ESo
A+DQrAxUE102oVWTumlfQ8QdFPQ5RiY7xbjIa6us1SjtMccwMRIbvU+l6+w5fts1K3zO1ZxEE1ur
xyg3t/Dm6MUd2vZtcOHeubQBjhZ/jhQLFYW5z3ypGKdOeTaLEXvaHgT2ljLtOhlPm+HSY+qoepSk
/R9NIc6xS5Y8AXESOiLuaC/lmWKQ3G8zXbcAG9YQ7fdMBRw/e84U9fX0PAwg/c/Mwue2Edg68rmW
/h4cBDk+cluVCsoYNJgVSqkM0rm8NhkyaUMcf9wlljnRHZcrbQWYcjnGBGzbIchadhOh7oKTQcj6
s8WhTVoqkwS6yRTAac0RlKqnbWKAZ0EsTl56JlvQfAaKRh/fut6myBk8iim2mp9tCRbu6STmVhOQ
sUgkg3OQ2kDcFCL7Jm7ci3kLLuCpIuKppFCzVnphlaat5GUcaXsM9Y605Q3PHEO33T41VhAEvoLa
MdLk4/4j8JvmudtHhZZkBuAKtnKZAS28ZJC+ue8G7vi8j62RjYshYtAsuUoLAq5QhySui4R3VVb/
xhwe2MGRt3HZsWF4diCflXqCGZtmmhJKqjgnzgkKX8kb8zZdVwhvW3X22wSZh4KqTd+PmpFO3H2/
aI8NUPrNZR3HzwKp464mE5xzo83DPzmq32+VQhMorBI/+lm5Mzg1moMex/Msw+FkyfycYzRdpcAt
oq6zMzhsiUCkRllJrTX3uYSGnOcGSghRZ/G+c2BY7dmeSi3fOux/IzhVrWhL56D6eDTiuJ/O5o1C
fELShSZ+1cbCq+6IqRN703lGmKpewWoBCqhp5WghWi6QWOh3zWNvN6syRMaqyjAbyvRbYNKpiGUB
Qw1QSsoxXmP9K6ya2rHRuf+i//yXmZSq3Em0AomVxgFONgEqVQzg9aPyMeX2iJki4ZmzNyL1ZnSi
QxsqNBpU2OY3htzjnBTvjuu/JH1kPjhcMKAw+rNYq9eOVQidumjublDEp1lUesegx5B/93uGSFvV
1T3JV1xnMmpxBGRWdg8hQx7rGQFYPLCj6NxhPyx5LrXKE8hLbCdBZwE6yjPMQiDDQ4TLspboP2U+
AcQaVV52xQnFVrEoXoaOFMUIGDLPwGS/6KiZ8tzbnIcS9qhEjNsZN28cwrsCck1YIvUj5UtTSb02
CqhddzwiyADXXVXHqdDZYX4hxDmd2QLUt5eQDn91bF06DwkJ9/RxSgg4bd1MhGKr+rj6JtfzcIDo
8zlRU+6k8uG5uZqY5jClcxM/BvzkwROACsJHdoaZKOYc08rqec6M45O+KX0C+BaVuMm3eXuBecJg
3zp3AkiJ3eiSiAJmSNruSKbO2Rgz8akcUHLEinanxQTCW8Gl9gqy5+GgX8+VKBJsHrFXWFFXSQWl
h/UafRNgdrMBsXvuDY3Zm4Nz+tnmfj4dFOxKAyr1WqdGQZrrkrOjbrUVdf8oFeZxp0NfFIOShqtC
o4dnVc1W2zr/QdvW/O/+glRRA+uYufk38d1adbMwAu5E+wDJ0DmXdUYFJ2rrdV3V6GxHRpU4X1Vn
SmmgHw9PL8badEcDHk7b2Wj/tA0rXt79GtmVgWWudKgRsLuZO6KNtTtTFPXTUpKABPy69Vnhfbig
ROBYF0i2WB9d7PIQzJ0sqbRXW2IlA9EUb/743x/UjuU9VfGH2L9JUQjwvnnz20X4eJVhKCNgg1QG
s2uID55/sFUsSX3uyYUCDP8VzV+4aXej84ySWP+RO8qpl5IAf2w7vEHDlF65gWDU03pnfqBypnvp
5/fuFty5OM/aTzm2hgm6zJD2c99R/03GmQVJReX726aQtWmWdZ28UMo600nQkCGkyCgbXE4tBL98
tbl73GBpvODbaon6awHMuX+/9n5jkRKx8H6osBkBxrWPcYnZcEMjhahYW53iFkBkrZW0fTakWsvn
tuUnX1CfQRgeKxMXwAi1DgI2+kMH0YZsmSa/A1fpnGBNQ2fuwCOXiGdI3Soetg61/w8z8mW6MXIx
0osp7OmizOYarBzHicoyzYMHvJiGeSLDLoLSsIw+O0LwO4lD5RhnZuB2JQYeNeVSqg6NN3q/We66
/Nm1tfbAP91vVDAab2BPB4JUyQCJQKJiVTedQrCubSKvm2JCvEfg1nHk/RE4in6H7zM4lh6Qod+S
1XqY+LpwmRTc1ozjPNaAJXZiHxqp2eI3ghSj6LuWnuQCnYC6ziIxWXLWsB6RE7bGXyXKfg2d/O2R
jSIIF9LF8orElFVvffuwK03GzXP4PUXWK7X/tExu4o28czYcfqdbyTcsU7XMw4MWPj0ZmP1RfRwj
352WB5i49FjkHDwQo1QSWWNE9iH00pQAisQOv6qJFJ1LnZGLy54f6ylvcTl1BoovQL+NGSYUI6JD
mg/G9xNHgWKCa68YnDhNmpn60yrWrzdtW1OiRMVrMzTZ3Jbkb2TclJMN6pOjOJsYb9icth/fCHJ5
l966URJlV2trhBTs9EW77IvzNHXyrC+88r+xyVXKgfGTrTVFDVopPAaMCwxjJZ/M88+EtQXaQlga
JXeaFu2XzjgBo32aL7Mc8+4RL41ykLGDcNXaHlZPxfzjoXsz/WwvH1f9pEMxb26CGHkxsTwLWNk7
bwvst5uPUO/2A1BuMXYyQm3EyGuoRKUpTzwfWGXAJzVLVb6s24FTdDz1CFHjXhCzy0rzGJRBIAZz
QZGUfl3CHYAWWXmGR+ILU8NhHSXcEG6m8s9T6B/9qHtJJa4dG+Nv6Uvp05AAULpVpGJ+obTDNNK3
q0ae6pS7+g0eBz/6aJa8z3mIjBkhRWlJC/tmyMlWdoEGHYWm3KdUfY36rD2TykqV8mYt6cJ7J0wt
G0aS5Aw7WhAvQPezy0YPfs9ZgM5DRC+5rkv+rsB8bKEHLND2x7P7+/X18/+B6WGr36DKmIvQ7tT8
/fenIOJqfdLfv3FXdcGigTpRRlTvk53q5aqiNLr/muOcrgwUT6iWDbbU4qWApJdnIMqJXO8DL7ri
QoWYeZNMxVu1v5pfPlT+in0jhbO2EgM1uCiseDEdKmK3oml1nNQi3r7/Qdq3nOe85QW0a6mVrOPb
72GVcaam+xk3v/Pm8nagKHHnEvlqyFIPHM6DrnDEAVZEQRNlB7607kuoVzF5OKqaV+QKJK9Nz6Hh
+0Pv00qKLcaEPg8fJMLoOJmZv5hRNlh+2rMH3UfuY9xSz8KSmbayOHGKU+ofDA95x+S3mRzeoL8v
lNBoNLrbQbd9ZqskJV/5yK1mZ5zNjs2wj/HavajvMkOvspEvGU46AFqm+mWIUtuyolNuLh2xjupP
GWc21CLO+0i2vYwvU/bSzEJM+nt/yG44cAeHNkxPhaVsI7MCfwlECP9WspGOLdSnGrS6/SiiM93n
HN76XNE0U9GgmMnPmKcqSa5Q6y1v+/tgXULhaHwzutlIUqmHc5upgSlsvFPWskq5ew3Cv7qfasOT
G+gBV2FLpKZ08p+j8nguiaK5p/0/2tUoU3e+XRvMr+sSQgcEJa9AfT97Pb2JuXZFhmzcTYnDJ9rI
M6iG2k+ryCp59RG97EJxfFrLNmvcn3d6LTqp9NW5X5ruMTKriepoOA0dX1tZ/pzmNhCERQ0sq3VT
SNJkHsHAjcToyml2sCMvbAN9lHNmay/iLSLE4dbr6VMsGLSVn9RDZlmaYLZSpM9eemv7f/PLfZpU
lwz+fZttZchx3nujFt68kLW3AynqdmmIF1jaYk16cA6CeoCFo1F5BDyRPC7FLm5plqsMNg64zwP5
UI3Oe/4UtuFw2mjrIQekp+Z4aBkeZ/LA7aYASMrI22fSN/aXBqKDjgy3lRD5qLC9w7GKTzXBsI8Z
jS7mICiHiRrfh3mNy/RXStdfQDy2BvRYSyciLlEVrXpqLEN06L7NJblw+zxMnfYiuCsBXKu3SWdk
GW//eWxLE5J74BQ7c0Q5nZS4imfpHJT+kvT80/KJPA5cBmQrzfvjDy7/u7YQxM7sERqVzCtwm5dH
aSVl+cnYTNYZwXfitl7veo1mQdHk50NtoOMz29DCBhA1S4lq/XI0jg7cwYektZkPF9ye+h34mVny
3x0XuFJSUpEnblKGeCsTVPGAqw4xQ9pLMofWskn70/YUT3BATgBTFHuPYn9E8/qSFSSRG43ZawsL
0NsByqK8KaxvTpZ6FfJ7D8YAl2f6+0VUlr2ECm5j6eMvB77WbhMimcoTGhqWirXtiNiLDyTfCysF
3an5x/y5wiqAShbc+eK05+0q9GwJ/k0riMRc/CYo2voPBMxotzRQPZjBjLaUQasM/S2J5klocNqQ
xD2upauPTigHfOhLJ8dR5oO9Wf+cGF3p88SDzbVkRPMnBoJjIs4cn7ehMOqgt41TdY7x1HXsa+bn
uHjS7FMXQOAqIBn1o4lq+o+26a2o9bBGCc2KyNB15SCHw3GzliyorDPLNMQuZw0/H0UzhCrhjXI2
f7RhTAdEDSb0HCjaWIgMEvw6PbR5YjZb47FydSScy3JT+vYPZ3UU9hoOsrunlh8vg+qNDP5ewFap
l0pfII05rmrx5EJXcv1+qQAZJBJGM577ms1c8WXd9x3jIRqWFOwsno/fZJBpUp/uP22Weh2hMDXh
5rdNwc+BWOP/xYZdvytWgC0rkLe8x+E+BEOfUr3mSpcgPhobF8DUScFrD/PvjpwaODl26yP6OtH6
2LAkzZtzsboBDxQIjS/8fcSr8tchBnc41Rer+VW2ffHcBtKeNzS/mLTh15zBN9Ffk5LkPJ4ym3+E
Jfr5BVTm3CB1nWphwGFTb7yWwhrZ5yyIyo1VU5woP/rmiDpPj7vouDUQPIRr8iP37do5GG1YOqOx
ojir85kBc6Ur9KrFhfoSEC9gHcCb0UL8WfOIrbfZgq1BvtDRyXW3YWyjcr4B21ds8l7hL6LC7ktt
nx+W5WSDkiF3xbr1MdsxIIkHVqgRgVDrQCXdg1CXmpN19JUP+UEMIFOOsULC04+lo60EaA5XI1DE
GXNcIYEmHQ+OfVy9v+6JetUGXeMhOk7ae5oxeehMNsn4oQJP3yF5AkEJHPXbxcq/8lFAJTTvO8Bo
WboIb7hQ84p9snOlZDOSGiVx46s9gTGp6beFm0AIeuV6jYKnxCuXSJl0cgNXSZALZvjVSRPVIQti
U9oeIad/fArl7ovjKT8exNs+j3kZbcQjE7ly1M1gZOGCPZbUvNBLAWnZqS2z2PAl4ltgaQyscaMN
92ds9V1VeGX+44E5r4Wzl7EpFWSQ2AG0qteR85FdM2/S+98pC3Y3gfYg6O9rE00fWvetvOycJIya
I+WbvHgXtD/2/G8Of05M8qRlQGdXibNNv4PGkcvxDBo19WceIbljy0TBkW4XZScBILAQxQ5fS8Cd
OlRPxY0M6SPPxIG1JzLF95kS0rluskzkApojqveamhdCCxoR16kbXJjgQFclEc2pdSDvxK0B5qc9
U1rUDzhC8GaiVBcQFDIyN2jMfDsIOGzFR7kAbJh6u06msS0LrlMqPSEoSiyLIZF6Clv3IH5XCII2
y80ww+6RdfsfAd9xkjsw1NnBfb1tpWEneu8IwDbVte8/WtVm9SMXP/19UFNDVgjvZy6I1krcBvD5
8IaFhgcm6Wz9Hb39E3840HWsjoU4wDLkdo+I/9dT1V1FUd4ssWz3h0MnA466QWphBOa4ON/1sSzQ
peWCK1sNO1d+fP/QMAr2N4vK7Ovnb5Y2No222dtLbtLvnosamOf590qrYcugj1PAvYhBYbH5E/14
5lO+5Muxioh1knxRshBMxIirKlz+ITUBfXw3sE40zJAEdrssthl+aPXt52eyQl3ygim4EagQGbpk
cI1okrqLIL/0RfLUDYgHquPiTePETfTPeZQWWVQ/uF2tb/Gs5qsDJNA/c3rt+Mdzv8+X/D4lk5JK
NNHQUubWfkVBE1zeR58VaNQFcAIKrdKSWhNzEoqSxjQ1XkptAaaPW+/h49Z70ExkBwzDOOM+IRFa
/Eh7X5eqENxFqNCs2160rSGgaFCih86bD0KxNgkl4ZZhqvrVubJk14Mxop2+qFFFsBC1KJjXTSuM
gMXHpeX7BWfdDrkrPfuL/QGgkDPQbaylFkp1Ztl143LjnXMDtXTGR49EeghF3ZEB38Vfhble+0sv
4CKEqCcs4P1D4i+LkJC+keejMfh+JRimuUa2a5p4qgQjkZsaMrEeNS+sMdU5K/qNle/Arg2JBWDe
+//JYC9l6VtVdCj7kT1KixZ3VjyFfjJ0LhQlNiQTKN1dwtObByb0p7VmKWcwQmSUsgVdTb7M7ZsH
IdOT60yy+fhgiCfxQCBXwgvRAslsRE+cTNmev00p+qD1F7XZAG+gk4+x32k0Ejc+PV1glX449YVi
yBpMeTDKDjVyqPIH6Eo9+TSXVaeHryIg4FIjhsduFhHp2NRdVGnV7A92r222MZTaawsaRNYvw99W
fLzyJxIYlzyqJ3RYlSyScqAD4gV0Syfl9h74ZfWqCerq3ZAq7qJREUNCK8JGso3zhXmPCzMOI5n3
eWleLj0AHmClZIAx5521Uzz6/dw0Jhx8vC1Mub/bnkpbqtEqvj9hFR7V+EkfNcLN4VSQWRmVlXek
tdf0cC8PTgpX+UT/O6hBlUlZ3nIDMYlRLotabwvTLIEf3iWE5BSrjTjtc7mPbE4up49PiTLTyuaI
jBfrCBxdMfQ+aDZmBJUx+aGYPtw6wU+WmRRiAWPIeOI+IIir/RxurikNJ6aKJOYIrFKfzF2OhvES
vaba2ntxlNW4wXyvCUOYADL7kv8MnSfus5weWOEJcqJ/W9v4fH8ta8r6+qOLfeGOxkwQfbeidT6g
1rQVg+MfsywNEpYV7V6B/rK11gxI1BwGCJatKrkzlrfgtcwq8EIfOZIEh8CtKKufLZqz+tWRBtYq
cIpXLYxbZ8HjZWZQ7sYJZJNnBi2GVUv0UrkMZUwZZ+lEs6UC6n1uLqkwlpLIka+epJhy/MQObDwW
G4xk4pk4S5cIgMOyKgXQDTSV0cKIfomdUL3upJ3BpIEzsW/DAma+ghoIgT1Bl+sW0uL1wjlBTsmH
QTIVagBeFqdf1dT5O9j02M9PECH64wTulxqQJoD68jJyCQoFK+OOV8paxxl/TLnnLys15QpazkEa
ceNp5J60da413L30mj4N0Y7Ayfj5SFcdC/ySdEf8u/+c+VA6IcyNo6dU1Qy8iAcYgnFfoEWjnOzD
R3F1nQU1caCfI2vcBsQ4Hfi70Q1tUXBoxMiFIOQh4000Bp10lLXMzYtI6qqaCNM20qPoihewJYYC
h47uDFPiYXMC7JUzoVbfOTXNz5hA8L9FcN000/OF0YuyTQjNFYL4N6K+/GI66yF0FBzdTfxC6Zf/
SxvV78Nw9I3bq9JuGfLEcAzyJ9YznyNDYHMMQjqE+kOwxIpIR8ChR0beDRYbMC31G1nUV9s/268Y
CQTPhJVE7ipdnBuTkLMwYcg6q8HumEf6whbVNAB6YOx3GLuvQFeswXa+NizUVoDkXqoMwkeSpaxZ
0vvLRZ0gCu7tk3TWhGTx6uPXZrsizArIyZRhDYQShYCchDagzWRsrguw80x/ltxqhozz35gsrGwJ
+zlm9nqblBhi/8rFTdpfG9NOutfS4ofKqQvbvDOeCQQuj5JloDGxt2jmtuguL4S3iG0OkEDVY9LI
uhlskIidC58TNhSDYCTDaVkjriCZxvl9SQiJnrHpc+/Mt/vc3l+pP1mPwz3MVBX3+ebVYl6ggYsd
WkJiLetotlhnUQwkKwUpbP+Dy+Y7m6kq4WovnWtb4ZMNSPkXelgSAgK15r6UHDaivKX8MakMkp/L
luQZPWQjj0MsHvOivxtwa5hIxZV81hVka6A+aNGwxZFOkbLYJSM6Y+Zn1r7mF3LLxWB6Pwb4rOiu
YIuU8qM8jPvJsbljYmHzjvk/Bzjqb3EnGfdwS+y3CbvZVKrth1O4mAfgaxCQQQOr7uC+1hyV+XZN
TrMRXIfYxhc3V9eRiCzW6GJUzbysNyNhKvmuc27a4SmfSY06R3Yd+3M8GYakg1irWKNXF3Msw00S
jCNABqPLmjyN9omva87rW3kpPbbbqQkuBNXqIsS7H9e+aLlGlItkarK6uKNnHpOtSzfOaOsoEz85
9m6SJ0Opz6hEmk6iRse5+JCp/JlbZzB1snEXJndyxk+QQ0HBnHvJZWRPEv2qm7eLvwUj+Uq2Us+m
hY1dd+PL9mYZ6ZoFtMtC5anJvzUqN2+3Ib7XEG9ZMdlvRNHcZDHb+6DM6jN8mMKoz/kS3QQkwl/H
6QbyOccEBMEA5i919N9p7a1mJ2l7aEQAgECrevVu7z2m7LHssXxnssJJ/++LPZ93tYMyubw3UG4u
0bZPbotDktS1mzQ7N6mrUnVwNSmZQtXmcGGD260zK0qoU3LCUuC5wffalJYdsVhxqhSi2EfY3P1e
XDf/UiunCSOw+hgVUXEt4lmyzD2ARIK8d7bi2BNsm4wCIM3GfpsDO14mR6N0JjD2z7gDKWCglEc0
yjplLyTpFczTss66MCvTYa9qmPY385GK7F+Kmf3qzbQxNdaNlRguCvqVMfUgtvVuBJgLWUVfGwiq
0YBdwcsXVv1XD1tXK5il32vwZ36z64WHFAUkEEtSXljpKvTh4Kz14YOGYTdv8molPT3w8rib7owp
3JNYJ7s+VJpRDjeP43ULk2mFvZ/PiDWOxzqiKbzo2+VBIYU2ko7ZgPP7QnbtUO1bqJDL8Hg/qSLX
F0kQYP4iWBfQHApMdSdTuL5FViluYFgaZ7ApsKZS8JKas5m5s1iNlyJR2Wz2jQ8YKTDH+kF05f+Y
CkdYZKK/231s+Ri4pBZlAQqXgUKYDOzZz00tS9DEvV51pL6qxn/AdYgr8o7gbGwgo/Rl33VyX4BU
F1fmJCgTNJeShMiIkwuMRrMWU8EblXVYeI0EHl9WlEY8/keQwztHpirZ5GIXoZrhQZKpn4BHLb7H
pR8A+7wDePImq+AHSrcj+4dqWjOpd4qoLVpQ8gwH8jY5jHiEZv8TCMbWubA3hstcS8IDXdR3jB46
5bN2AjMq9XUBrczEE247MSbSd18+bg3mAqeAfAw0tEvm8xTo1VwrTxNVCAiA0O5WqRKI9MCQP0kd
x5ilYQLkDGpDoAef5KIijwdbNqL2eE8hhZ0Kl9mW/ydBKBOxFZ0s9b59HYQTxwb+sxSESb37jasm
NUV7huhPKgcgMBAU1B9Gs7fCGaoTVGkch+Go+AlsTJELLqYx0Nx+Icle3Yyv6Nx87t5sBG4XDsLJ
DSUJPr0QPkm2qZyM/qsZotj0MZRErvu0D978j+J6hAnx/on+yZCnT8wSo3b1KfJDyMxZZ+sEU3LK
9rgtHU6OYTnF3PHxpR48cQoyZn0u8cqk9bNnLHd0c5hLMVmxEROERsO2WSvm9f2D237Cz+3ukL7r
x/F/1JhjiZCqvV026PpC09vmfduQqcp0xgDeAAx2mzx2m+TxTcvD10mwC6Ko+XN1wPlKjUoWl8Lu
Ci7EyUNepLrdPPbf9gdAT9WS3xhj1C2B+6y7GK9UdgMqaztAj6ONloWNqrxycUAar8tvyXYpzelm
HeWvrkVWcgkI6yBEo8M2z0eVK7ylkVjU4P0feM9aCTP20jFwnaqq/8C9zFXEL9MX82nRjzKT+6cO
K0Ev1zFlG77hcQGpaatNZvu9PMzZd0UExHcZUBcJeo2EEbzTSZ1wK5GnBP9nlyQDKdXaAIQB196V
bKFr6n0sGpKUGFtGsR/j1WHrF85/jNhSgQgxd50coAhUR2bIt4RuYcrJn/6iSFG2MGwjMt7ziLKB
dU1yFguk50IuVgmQfMw2aVxFmZTMUQXB/hj/ZpeVx1iviI0Bwbl79YYhDIW9v8M3C3Rb1cLm2CzJ
zzYvMGB8tAoYj91umU3nwQgdMlAmcQtgpNhfZFdj7+vXrSzC8uWtXjk6hnlTRZBkDkmp47Rowp7/
lvZdFmiSaPzZMD+zeGlLscuGjOz+NazUJ/K4+mErJSvsekKeQDw8EvTRH6/hPVfTLzqSrYQLKzfv
ex3WQnJWGxeb2Q1O8zQrdZA39gLbmPPyVszF8nNCBEeFMmVpuWpAtOBPrKP9XphSSsG0NKepYqaa
k3lpvkJ7uGDv86sDMRG9EGqaGSl0Smz0FbfjG0pECLHzkGzpjgViSmeRiCTlRZFGiqHwXb++gb7j
5cNXxhFkCzJdlj5qUoLSKcibNzcrQH94xBunHxkkJ2pSIx0U1fbdDHcZrxMQIDve/Sw+rZz0YZvu
72Qa8zADbPWWMDWs/IRg5mzHbmNocAFaK0Gr7yVhJOGMkIO+21FsLRwvAOknPstupGv1VBHDBCJb
dxB6tc6G7lsqVkuhMcks5X1VdRrq4fmxCTmYB9TV5WFaHNgqXLx8hghwBKvr2qtjE2Z+IXXKNAuZ
Oqj33S0ioZfuYlX6cAsHZn118v+jriaAd6Z4A9HsUFf6WZnZxn2055jFL/DJhG3iQQQMr9bAmKAH
d3s8Zru3826AIEcatI+mcjvURX3QNZXV75UjuWFPziNBUeq2Omt+xrLtUq+ZOeNcrcJcApyD+Idw
/gaQwSkFK+QTMfs+Ih3wSgtqxZE/J9CKJDkiPZO2L4pARlXEHRP4OBN5f7fW9wquQvO1vhuKNOBt
v1wc/ySB/B/GHT/WHJmYAWfvUtSTwS6tCRoX15l7G5r8PBjLt67YCWQzmzOr+SyGuoukapbRT1p9
pg9WBj3u8koRpni2ySdJx/tcJe7LgDQFw3fdCQDuxZebvusO2tm938n97zSN7e9L96COdhy1ApdE
Uv0mtz3nH5Z8csjJ+3Ph9pWuRHitblO4mCogaUcrSoyj8SKmQeLZZOpGtRlJD1GQ5TC+8Rb7QTx/
YBv8T/6edP4BARXY0xE7IXQ0vYV0HPhmZPR1INq3mlWALHdjp+IVPpMmJuihqPJ4xrClQeyVsUVK
PRktmcbm8KP91Ot35l9O8yCe7jkJ2RciXmLXP5TYhGe9OjRQDX5blm3C5kdLoMdbTH0ddh2YTa3X
XocvETx0pbbpFM4McrrtaEOnboWyV1xDop6Z/mUjqppBZ4ig7xfTWxKkC90shFsT1fhjQy5hmTtc
pa2cq/5ofpJiC2VRf9BsmFNZrmgoPzE3hj3FxYM2yMct9ng7x3EITlSdqIKkL5hEGDKsiFxffBmI
e5x/rDYcmecZYd+py4BjNwMcm5YTMBEUb/D1zLJblnL3GeJRhMbEWD0pmp5/xqDwAQSEsCtNw/xW
mEU2oiKxEpg5ypUViW0bDdXdzZhaobIw+Ld9q5uRckvkslqcjNbpYk633AaFZp3n06+Ea7dIxaFP
Gn1lmtT5xSrDb0Td6aT9eQim/E1aXCTpTGUMEx1Pnt0mN2Vuw2LFUat4sgHxRQ34tVfyiX7lqrTF
+PGqCyW3GbNZXoounhxHNwMP5jdMWRhjHPc7ZmUg75b9sB8UPJQAuQ1aW0/N9Wqyj5Nx69GHR09y
UoMpO1MNtODV79jIVeCeM+hUj6E4izTf6rz+vWp7Gt1YWspxJXHCGA6nNCaraWsXFPEeiuNtDRq0
Tsu7dxluQkQb/st1P8aCcKlqr1pFlOoGW2JK6Us/3HslgRG1ePa2ejZxIs60jtvASpHhPbSmG1Fm
5KRp+hXBlZTwgsdnNEMrbc/Ml+SpsvQJK96h4tbqVpamfM/yTL8QrwinISJVV8hAfnedKrNEO0K3
5qi8gzqzGup3VstrZ6EQCAyqk3C+8XY0NXyptGDvqwxRjIOMdglyxugEJeqEuHdQqqqg4zDsqieT
VPKmBwzB+8nybTERBLBq6zL/DIIxBwFf7VAhD1o/1koGhh0hShJcVsARh/5acg1hDAjRcnItd5xM
+rDyWVD3rGCJYv3lcBGOw7v61TlqstcTKTdVQ1jXfvCG7F5Y8yZqgAQb5rO54EtkHpn9VmRwA5Mx
vDrWYD7pbyvYNdd6CN1kvdM72/v9Y6ziV1S4f0mV09sJkZTfGpYDcVLiyJg8pGVs9wuJdY6lpTlf
DAVrBA3kRZabMobvo0UVmFxXRwaRdZKN7mMkvZxh0pr3byzlEa3noNZLU44mWQ9yCMwwLE+pklCA
KrMpJt75ePIW9EO+3ZBtyt/5/C8Dp1+0cnzC9DEvjct0vpwVxEqb8LII7Vd5O54aKA0gd3dvZBWP
c+Gkwxdr6IPHJox8XsPakydnIKXhj3HNOrMxgSVn3TlpL/ZfASkEZAYKj8gVszNQSBXJoGzcF7zl
7gQSg3LUCbT/DjQDyqTc0bX8JaAQEVxgj6HcXQN9GtbVU5F2hPcPCPmsUpaSSQA36GKtWczi4YIG
ps8hD2XpsLF2sS5uCJoEHfIyAQ+vN29jkKBhB0htBgYyc/U0OPeLcZJqR4MKc/IZnzW/CjbMv8pq
c9QtQVvaMmn14pI+MR8bsg5eh+u/wGE7r6gQFkdKxLr3rKLwtOhv3qpSQ0lCU5dsgQqj8+OjBtI7
e/B+/yefWuqkeKMZwAeC9wiyTM8HJbrNA814qHfXGYroOZhJHIFBVIXHW0pK32+8y8hyUaGNVLzv
Us424+pH/HJFw4Yq3tcpB9XikiiOmVJrcor6d0/bAe7PFm7zawgSirUUtyOqi2ZOkhKNtQE+JD/w
V3svIzyKCwNznAshTaSsc86ASA3n46pDsScxfA7+Gsw9Os9rKFjsD2pryCHS+7b1WFNlHYgJPSar
C58owDBnwJaDB4vfH6+zshqO4QTU6rt6gdbp8VU4rep+m0+AmZ2eJ4UhCCTEfOkV90GeuJpdjIdW
5GWWwsBHE5dDnavUDbobAxonn4Mda+CY/QU1WufFevqmDclso6/yEx9YA7JSIXsqHjVnDInbbyjf
vJGjV54wXKKWAymRKF+BghGG5UT4M8p6S67yijrgQbggkZqz2FXDcQ6gWEmlhnVsWNbfXFjm6Orb
RLE3DH3y3j4BsdiMC/tMs2Sewdqb7te/aG845rwcbFCeNrescPOtJB3Xm4ZYReZ/h7qALsoqeDIh
MmB26/tvhKlLhFWRa+4JjLOgw8ZT3ok2b36loJNJJ8PT5J9enVrnPQm8sDNbVNoi6BPSZcz1eA+E
NM1OCTZ5EbnqKaFd2gIcy43jDXYNwB7V8R7bi6CWVQrL638BUKZCzAOyuRUVSqM9XFVbbhudFyn9
nEK4pUUs1TvQ56HEWgpHkbfBcJ31nRRCF6umSuoydtphUL5uJMnr29/7Xsfl00eHU/QTsNe2sXeJ
i62Fb+a9PaqsgXPXQxxij+o7AwbleV+IjqF0qb4q0dGHB+WcMgcp+ziT5t26hWrB4yxsO6ZQNPoA
ORh0Gn2idAi1Nn9P44j18m+EufvoY7iEtRwqj85sKdc++V/rE+qb89nap/C5KOM/dntL58kJ7T1u
EJyKPqLXAj6Ovh3wjzAG7XpxPt+7AWYxb5pQLnPYBvTB7xJ9BVybD4iwfOLTq/+RKI4yayvBZ1PK
we0YMIrfsJ6UmeJ0POFiuzFS49onn/FgiecfvSU0QqdM8ylx8dR3j4iP+UTVVPXbb+vl3402bIcy
3RlEig6cVNgE+sGrqcAGuUYLLWoZCQGAwPo16FOTt4+nM+ghOeYUfO56pTACwIz+U48d2OyE9n5e
0JdyC1kdpOxMxKwP8qfii7soMUQ8bFl32Z2q0WjsoDahdo2Gd+9hLH4+29BdDCXkQPh8cA1invvo
1MIBbGHyu2eWDZhU+z4pHK/HSLgfnM8FdxwzkYwGJUcWYwANSgtLoENuSTddCFUEgED3zKgUEiia
9hI62bQFbq+lwNUaTQdtraj78odQ7sxmLFlvto6AsaBsTXjJ7hTkdj5aLNvVQtlfuJ0MGZKYzX2e
Dj/55BaMxyXmuQ/eRRrwvD1qg455OmY1RjZlw9UzdiLSbUb01yecD9T5u3HTC3oZEEF6CthM7nvd
EmgokW3ONC/0PPZKkXzwKYZBg4GPAHN5gAHAiHcaAsebxzo+OiK4YQuKMvSQy6smoIzZ0zXJbPXI
KG7cyIglsJnyPwuJqf3kSceO7rupqJjnkLznmTPLXuTuU0owfY6PDBT8vykpo+gLhVb5GjhaCMEp
J3Dra/Wlf4dlnfBDJczqvqJCxPf1305dMlqs1p9IWzNaXBQFtb7IISkHcVxU2E412pGq6G3+kZTj
6LqXDkBaY8ADVxZjz3ji7mZgaLRf5r+rUtFtV2tULKuRscoE0aI5KoxxAIHBwoCtoTHsxR0VFAqQ
3GKKm3ZmKgEgu+5WyoC8SoyA8OBanIclKVR1LMaINpyMQ3+C85zj2YgICapzKmu9T0u/nyTsAd82
MKZ2BOrqd7Z/SAPCItRGkLHj0u1w4dhPH+LppX/u5RSZfEcA4bJobyrmslf+j5zUoib/wV5p3jlc
45I0BmjrK/OV5Qws0U/5ogNO4DtIDN9aXaVlIpvWSJCcwEDRvmHxDFCxrx2DXfgU1lfsfs9Vcy69
5LN7ZpfK5tnSTK7kH2CjGVNgTVP/FZV79BVmOXWqIIBfZf7YrB1ICPms5e91rIecve0owCSyWUUx
vBDLqDItiOuiRpiZbEMRQfY4u8zH9GlR1WGnryoGlbyRVjg8pT7IUEUsCUx8ZrI+53NNhO+7Kygq
CGITiNMPz+SbsUkLAfZoGBAzxzwkYA6M/gjUA/vTQCd6URFnhZ/p3mnqdjOd75ZkZ4vUncQQXTOa
BtolgYltRjHEFtMBzOhUH11zvRdCYABum7idV9uAQiUz8zdbF+bVigxKKIY+dXmqAaerDvyecUtT
dQdnlGJJggfUI4PuJGUoOard4vcg8+uM602Og5qUeBfAoXaCYi1GsMLMRU0FtLDoHgYW+cvixjzh
6qN7E26zEnBNzIRvFH59HSAQ1R3oVaWAwyzOwGDSCDJUSruX/r31fCnC2/2zQDj4ceZSKvq17tFP
sfObPG/489g3hbccflJbFxHZX7OqYnDtC+YamD+95jzJLnEA4lSYuVEvHU9c+28RkV1WeqtAb9So
Io/xq+uUkKmvqVUpdjT0CFSltRe4wMwFseKT6Zgr6Bh7cX68hfP4VtoYjNxRuyE8J+x35dCmXTts
ctsO0xpzcX8wwGLvkJPxg0fV85vaXoXhkpADpOtNpvLjHCMbCQ1Yt6kB9tbSNFgjw/kZIXwam3c0
5886ZToy8cft7QJQEuQePQ7+OnYmeNfmwe+uaeKYDhURjS9WGkx/G367QVXJ50R/5+28H3fMMrmq
W0PBBaB5hrPUN+SstiVdUXEnBA5CSKwYZWlQOGe9SqQDkgfbDjhOdTc93bBpMCIPuTQdS4K9XyOr
R/IKfKcYWC4sDlgIv3uE7BV+j1vbZNFHHPxDGWCgb9KLWuo5n8BRDknK4dHGPqBoxiKuF2nBXA1S
4BpvCAaXXZ8DOi4Ds0rr+Cp+vNYNnpEhmJPaQ2J3q5cpMWJmDNGzL530yxflZC4Emv6vs7syUart
TBuky8M2/WL2hQ+YxrHnoQqSyjEMhDFejpRexbXvtF516hpVIunR6xLQRt1hYJ/0aXKCQgodlzj1
FHyve2Sg+oY6ZZ35HkYk3BEeAV5k19UJWy5fJU0kIKUYT0doaaZjo4KuRcokUiAm6Qadku5XW9MC
+DYA5VynWN8x3rtb3Yo/+P5lXT++rxOu5+R57S/sX/ZtI4yXhRQ2AlvjaPjycIxZRxRAEUkLg9JH
Q7qHHiswK0koKEgEvBweXRD0a/RAf+bA9l2+9vK2pIAW4QKfNnq4U4YYPumshZHpOb6svwFdlI9b
NIAwCH+hckLF77F2w8COPXmQAFVteq+vjgmIFX0c9CO5Wd/g25byYtZI4yQMol0U8Knv0IZetNee
c4LWO96drumAePkz8vHXBsbjK88GXt9fjS/5KuDZ2EFfqN9VQRbKJnc/pm6vr9wa0M/2x2zdQvZD
5tthMhSOrveJnnrb2wR5F9FJxmUXU1uHJo5q/Q7AwLeqenXbRZufGWHzlMFiOUPisxBm036Tkcl5
C/wFWOpU5QlrNbH5uKX3ciqPDD+AihM5DCZhX2cHHCT0wVhYrlxGLUPNWrARrItiK/xyzb/vt6KE
IK4Yq+1zPha28nLuWrPyoIc2sutiwtsiQu2fcsEcFW+/7yWeUlXgZXw0Skz+hS39oGSEcJbIC5Ud
1cPI6ek5spYDX53Bhu1g+pu55gx1IOz0G4WyEy1PxALbu1+nfOe692ThHL7oZsbVAxI+CzSvGfrJ
vyMtudwBit3+N/uduTEhYb23toz2tGBivNXOQKPJcnEq6GKvwvalxhlLQWYlQ86X9al/ZaIl1QEh
uifvzr4FMN4ax77365dpEeTrwknaOJzX45aStEbnvQrauASB0Z+D9MsaMaKcvmZWiUZ7t2dCWUOl
9yIhkTzcd2QEJbtf157LKd+VDqqlOITsZXcQKPrJcW+DZk2PfF2av9c2wcACaLSn7ofEbOyPp+Qx
Z4oWBmOlIbZhUryiajq5cc01SUP2FWiq1QK5b/3VYWUuoq7gYEQXEnpatlR7xoXg+Bd2Wb/b2Cyh
0RAfvozEC/nEgbp7T+7TWWJiDOoQW+aq/FIcJtP87im6qFy/IrXWjxF7NV/VACM15kf8WHzctXqB
8s/evRgcu/UJIbewvgjFsIifb/MFPvTszpTbT9GUEUkYSRrZiscNPxC9UQqdBX6XMydSwUUPyllA
YtIplBtI9pAXOnS/ziaMFpn+sCdyH/QR3pHQmYcUHRJ/K0Q8ADKSOCh33j/Q7MTo8fj8h7utmMBg
+bS2AvrHEL+4SdR9hLk+cvk45W8rhR9loiv5g/cWfFfhOYoUVkVmr1lsaMlEBEIZNSRGwcK4Za4E
FKxGv3Oh67mLDL9uBGVWvEuaFnDdtQYezmnGtWdfIqrgCgk0lJvkimW+i+maTCadWi7DTqBhrZUv
CUUScamOjFTJ1vvvWlSk6sCse7CGr1fKjYLDOwIH+HC3C3V1IJ/UH7wWVPsMW38WTYSCWq3vlZAK
FCFYVxPZ/zSMQLChWpA4HXOMn9QIIVgqaEMVam3RkZ5JeRv86DKIMjTiYnal6qjPuqHaVZ+lNBcb
C425DtNE6qWmvbVgKNKDfCW7xlskMAq9eWrLMgpDUoLF2Ec+bCdgeSSOO+qf1SaO5eYGy0bPoa2p
In6Pb+j+FOQapHxCf2r+t08/xlhBQOhYH/wF6SKmnnxo0AyMkY/I1RA0L9jIEzZ61HViS6CACylp
Caq4F/JVazCyXy55rko7fKEMhn308AvfUUdIYWqv6pTRJHCBxRiGo3AiCEZbAVohpTSBgm2JkdtH
WNR5Rw+NfGHmHAeVLirmUIEqe4NTIPyQQOppWM3RxETsXnpDQZWh5JoXUzBg9MevOEi8QHK9Y8l0
oL04923QIirD+Q5DIQ2U69WiGxi4SlYeGua/R7QKXyGN54xWfM1bSujza6kKvO9FLpAO6SaIjmLt
cxYIAq9leQUyiOH4YXkDV11coXwNNl58MoJDrm9AwqVTRwbNuvlKaWMterH2hHtXQjzzey73Caiz
HOe6DPFYsxsq270AgOn+YMSaJX2UgsQIGYe0KaqSHTfayTVls7UJELfPk6wQNBUvUf7iD2gP8tQC
Iw4MToa9pgi5Az2rqz9V5kI5dI+fAndTF3B6oxz80rzgbk2PhZJCCDJ8IwlesqanVGvtQyguPenc
z6ZvGQOy2pgD8Zn97Dn3VMkTFmqkJDQzj94/ZEv+cQgbnIFxoexIjAAizcajnAjBo9JPJRTMqpEc
28QfQVf35H519kw0Uz6lpQbKw+zr240Jll+7zxgnmZu6ZQu6lRmiEqDe0LKpzWc2oU6gAH0/em6T
SWxtjibfQfb5Zpm3e4DvofGwMsvUUKvDGgwAKVXdpg89fGLFdCwUB/vyUBGXXnqbMZN1wJdTlbue
fU/Ew5xeFiTsWd2xr/cH6Q6LgpO+IFJQSjix24OZMcXlTe04OZh36aXzIu5K/cgn3ZicV0E3iXYH
zk2qdSUEksSIbQmkM4GLKYkvrd20A7mz4TeCHHH2FSJiN9To2AhydfBITmqsxsxkkeUvTKbtqtzb
PsqHZ3rrd/CpDUJomimEAWpOOPA/ib8ZnzRoP3oy7Tq6r9oubvLcjO2cXAUWYcqTINLl8ViM81Wg
dJ1lUgu8LoRppX3RETzLb4Qv0i0MK7fgYshIy/ALauqbMQ1Qoee537htN7KAWxxVHlG6EEsnI1/I
AbPy6NcWo6H0BXDLZ5d3Gf/6tM4VuRTvqqDKrh9IU2Yfi39lk0w5KSjIC397xOTcpohTTZ/C6By4
sElOqndQUGYyFV6PkYQPMAUxzOYoem+t+Vzthm/eldKt2ETxqxO4xkQjpY2dHjr1BaMvXhUuCRlc
CFxexPfNigutrymINcllEMe46Pg/bO4dexuug+2ikWWRwlLpbfJO8+sI30LublTND81qdf2kw8eQ
jRATjb6ZHJEA7gKXFsLlMvc9+NBulfwzdnWV+9+bsEIR/EQjiHDaXMnw4Vna8vpd9JYZ2q/2UkQH
4DJFK64ZYiGpe8YIU3gqoDF8dsVrRqmECJvhNTfMCf7Azg0ztsSwD2x8o0Syal9IAwHvqfq23KiT
9et4LsvGybRP2EE3lXyVdMeGUzYylzxKJVKM0ocwMJu+W0ti2r1t1hwItmDcS5lE2JveQjZeDZFR
TNqOm6D/v/3nB/FVj74dAdHVp9ENXVmHnE/KgTWWtT82HIBiHr1Znbd8xyTFnC6Lzm31HPrSTV+2
ISUgwWeMnXnjfkDDPXe3xcE67XxbGg7L8COI7qRPzsN67fQlaVgO0PIYAQDwMe5SgJYcrMu8uqR9
RhyYUr79MLIfxwaWQe+2ZOw6BBlRT05oZ1wzBkjaLo/27nEx8tYKDqDrEyj9Du8dCDTO74mMAdx1
XZmDw1Q0OBUj/eCycogAaGV/qmGfuCG4jbb7Rkl6Y1Lwe0KGssZ87qON93XhpWervowVj8g9hfhw
bCDuGRHPEUxK30uPEkRURSu6FhxEioCQFRqekBYYEeeETD9+KD2cMSbyonakUjLxBqxe9q+JtAhU
+M++XAicraIwYwAxp3WdkzlIRZbHywk83+oAyFVWbdMcB+anBsOuVXPjMY3koS2dYJ3IiCJth1uG
+mbo5PYJZW0lePnAXlyeeHoLG2PfkmJUF0LKh+NVC5KAdNT9XgEYz0CtbJ4xNCBHE/WvcpUuDZPD
a3cDfP4YxC0EJxRU7hEotLv5jyqcacgscKaYU9nLhbu2HvoG/Ab0UDTqzo0ygr3MVhdbABa6E+0e
9SW7lf8jFaTfNO2J3QEdXm/cT/1mzIImFpxx6W7QVGgyWxab6a7zCSgCy9zTFeGprF5rbRf31HhY
0TQHAGGgCP4BPdTwXiUP5GM21xafqgXxo7rfTeQnWa0nVxq/tEC7EiPmAbUVBG9rBHtuiaebVZC3
aXdy86OZEJJA8RFRHBVkpl75tWNVRb2ygLAebQTZqGYSv5DPzC+myIHpLTp1/Vwk0XWR2bUn89o+
y7kAtaNnQdWnBwvb3zR7WXQMfxsl3uZ44gyHs2N0qEfPQEoFljtVhVhthaTrhBP2/531ozIUNJuh
8tja2jFllpI6/V9rqEEiVCOfJhxP/vx34jfp9b+TTAxnpvLWiXchqRyeOWtnhoF9Dd7ksLtRnm/N
ehLMgcZFhMsLJZ74eyx68oJyVidNdjoClYVrN+mrEXJU0DPXj4H86DAjaLnH2goSyuuD8d+ruQy2
i/REBw4kzpO5cytlyErgAXaItzmxoV3F2KUlJR4JtTS+sKKwQr0hzzPk4mPyYMTwsb10yvvbbDzm
LZOfy7XvUb0SgVrsXcW/81bLiD9NnAFBeKKTiDQHQ6pSbJDhQfRUqMeN28n1yNs9pmt6QFGK2ioC
2TMjMHXZn06mVh2GM+/YkI1oAJh5hfQkSiU1N+rOL6k3+jpAYIuO6OihGbLxKzdDLg9qmI3XVWFn
EUJqd0Hp5Py97WDNCX/er84VZx9//4kt3FvKhtI+YeA1FAxslYsx7sijkpKKNHUuJ80FieOewQ18
BcC/4J5Siihvf+Nr7qYE3nEZTIeHro4WSr9noYuYPW/VGDZQ1AiG4KKYZ3Qww2ryobykOA/y2og3
2eRtBAPCfDX702mhSfdo62IazYKzJGWW2u8Z3p5A+JymiD8G/ZESlO3nAc/SvwTq/yFe1XwVFcSX
1ShoA+hctXTXDM12TdC2l1S/jM0mdOl2loL6mDXql0YnTdbo6eFG6PSIZfOqZMDmmDF6ul7vGyVU
Ju8+dkK3TWGFCgRzwtqS3N1a5rureUP2Ypiva8Gt6VjJfylijcOa296jeGO8EGj8jLp2em5eOAWT
0Ason8da2F2WqUPgMXeg42ThLJMqm6hnolmdnbRs9xyuk2mib48k1KozXUkFMOAroEvznnlZXAMY
4f9ehql4NsFJ25xqL7MmEcRxUvnUjyxyHuymDdH3KUssXuhzd/n3G+IJXtgaj/Oxqm6qD47/Ex9f
MMk6qz4i3j4urdcZt/ubqN+GcHi5O8Vnj1La21BTSTgnmnTIfdaur2ggb6ns0kV5Jgw2ty+BMn3V
vDI/Zwyxm/a5mYJrRE1sghcXAoXTaA/90ZKRVT7sKCjhSUB0MvsK/6jDe2wD/z6/sMhwQHTDVJcu
S0+y0T9qHbhcMD9KpkWHCqOEQ7CNzwgmmIA5njRWYp7olnx2iz762pu36yxia7fhys8SP3uRn20T
tfKLSDllNFfby0izB045/L5tu4io/T5zN6Fu0+1SY6oEd7GuKS5NqIohDb//s5RLIKFC7Cp9e9we
RUyknwMkJ+xrL3ccP4rfQYS41iat/uxB91SGczwdJS9ulzv8j89wQ3jkVlgDhvSsCbzF8vY/kALj
TAdi2pWtpkshdA/mS1msfhdw2e/6/iLBQe/PHhGWsJG7FA8fhcr23Sm98PDIvYOyW5atvtYLv76T
Y6lKCTvMyRyU6OPOtMT3xPLKeO8MEwsGPOj/LQMU3mX6dQso8xZllKVI8ATOchURtTyD/0RbYj7S
wITcSGMvDzjAc0ozrv/zJ4MN2LTRtgwRqPIcSpSaJkRbOg1oxne0s9tGj62gG17vLwY+hyMxFdPj
rRefj+CT4PCEa/EaFYiFyaZ8JFvnSvGa7vf0tYC0j9u+TIxteESqqzO5ncS4UyvvETYuZaH8XPy6
YU96JtSqfrZKUkgGsTSCdbqXUOrWOvNPqnu5D/wtvnegGPSpRfeEVFLrfj+eb/6fCMjoT89aCscC
UOOTBP+ildrPAxVuundqmOqDxveSd2mozDvHTu2MDn+g+fiOD1GIxcnTsyHwGIiH+enxyWfW8RRN
XJlI4cuKQNZxxXDFxhkfndatJLCj6/NJegeESY6wuQk55XIU4pRqCKPcyD3zQIrzHsayNlnYud+Q
UwSAgOOEEylkjPI5OpikZqgNCH/CI8v93KBigtbl+bA6ByuWybyEL91X4Mry069QBI1Zm598gnd2
FJBZ1IsWUH3bGULAeROX4HffDprZslppqHzpT02JKCJ+kgIuanJEItrwC47YCTT623E6Er9XKZr/
yMMhc6bq3+xFfU2ddf5fVMJJ6Ruojf3Sp1Qj3o8w5w9T1mWfC/xMKvGgeqpp4F5Nt3F+41jIUPNN
d8L2B0Qv3o/BVMLNGx5fYr5VZJQKdlsYtabapd/4+2UnWs8qDSSp4nCr0/nzAQ4gc46kzGSzDcMk
tyAdnkkTb/YIlzpwTQLisfdwQf5oLDDeFVev1NOONcmnsO7XW1hISLqlLVVTY2YQ96BBJ4+RG/eH
d+N2cCWvmuiWa/G5YZTTzWQkRU8nT93Gju2rgF+J0cKqp35WS9L2ZDJ0z14ajamM1jD1BK6bVTD1
mV84BUBUpeayYnJih12k7JFergS5DHVtWIUID1XMD9dO2Ni4fiTGnGkJL7O3ZTM3ZtR7AXTcB+EX
pojvSKDAa3t3nSnNJSGv5jPbegyrbrTYKcKfiesS/V5yG/MlXW5ogxUokay4xfAXqTEVd1PZXenz
eaYCl4Eb1c9YRfOnuo405fLnFSBBNykkGeHtu8gZ9z8JuK02RKr07JK/iJSh30V0EdndOqWtmTEE
PWZ8M6o3u5Mzs0W0AR8VOwq5rz7m2ppoSxjPnadOQ9/Vk3STZEdEzzOMoTSIJIJ6CHduhCY3yIBa
6FNWQZIoD9tEmM6wjK5751RONoEcLk+5OxaOdMg4rfpI1BJY1bX3NFFFT8OzDt7nut2mk3pKjQrB
r1WTfPT/DBv7JZWozCal28dMRTghZIg7nYZ6sDPDn2+zstBmpj6J0fIcefUeaTHLOLFC6T/TIRxd
yXWd5m4z2rf4yuCmoGaBCNI1j/h7z9oTXcC4SJkKk/zoFz5tIjB7kQlw2Fl1Qk4q6I83zU/KgHIq
3O9IY5OeMmsdAF5QOZyEu7fnZ3+fXzAFbCgJihHfyrvuM+yUKiZjQBCOrDJdXBNuxQhJ1fzFBxg/
q5xpHaxe2MOJYY6WeCxXg8LY1UElAvoLTmesErRslIbKpXUKyply+kJ4tSOQmE6hnFLyCCI3qR+r
YQdU0DE3Zf018My/OrL1bqp6Cfj0zKV5K8RvCFUubK7BNehqgk14Rp7l8sHCcoR0G7WRND+/Qf/B
cQaA1dNkGQ/Hj7dMvrFTv2oEY3GpmFENvQakBrZAu6SYis1cTdWXe21hQjOnLMWg9lT25qlEVVFb
yRlGh4hrWac0E+05OnBS6IknZGj6mfDmK2MNI5N4GiHdoAtnmJzjEMgEkJBo+g+hBJRwH+Y1bSBa
H7514CcZuerhjDFyOOWyxeaDKQdVDTbCmHYua1z2lQp0DWtOmvfJRCxFZ7pi35X8SLsuTX5yiM0Z
rigALi0fjPmM+irYMrxv4YB6qVl5VpBxGoSh20NvsTJQ5EjoFUCjKmzeXw4hzedG/qIAcPe5tQuI
NXiiLPh8rS1OODIDK0HLfH/9qBS1Ly9nTk8yKKp/q+e+E4FHz/05pQ8IA5EATnPyO9mjlMsBuewQ
CuUlGRqoVlyaWMUgDjOAZINm1VgEVtcg+V3dWZOh9CMdrmde6/ADlMXEpPIAvda02aIpJbzsgC/E
h7hR6plXspt/06uEG4Qi/02n4uPBU/mKzCT3VGI9MhgMaOdtcCIRTtkjemcH8Iehwpq5zVRu0iGv
k4jJgqznaYdcY1i78HvWWtJe/MrOs9GxDhoIj4HXgsUZF4tlKncQSVinWbMey3P9hiUuU2A4tyn2
u3QcxriXr1pUCunfWoYQ2QuTgZC4G+pBfSiHwvHr4og5Ip/p2miqjhA/4iBMB+F4Zf+hbiWxF9YE
6rxm2+Lc6guch4uFMD/tRXy6ToFIy7Uv5Mk9kwFliP+C8GTYu+Rozn+SOEDpZPpb8gv5SCaJBwYV
nZ5qPiSzoEPLkB0nCdsJa5UfF+rP6v3sKVncmyGbrYuy/OvJkC7OCPQKFeLKZ290g7Y5v+5OF1UX
CBEjeuzOjKFchrf65cbJxgacMQqvsV4B3tigJuzdId/kBtyC+bpHbyFHHt/7cyw0iohBo081bMY/
UNTVUoKySSrJPbO70kS4CLDh2MjcS0tpR5x2EIi9NqjMKVJp0eKrNxUuXiWhceXac1Qe2/f4+wq6
9Pl+Px6QebkG4NeTO4Qy+56Ep+qduv53rwHrvmQf8ODbWNWwZBNqpzvTruMjXxqSFzvGfXeP8fKC
b5dj6L9HyO/w37IOe0hKjyeizwqLIThA5BiS/TTN1Diq6q4cqQIZZfcS/gFoPGrmess1B/rKqxMM
EdhtT1sE0ru0OvniqIgideuEEfoHspc2xj8YF51YGIZa20T+Y32C5c3sTn9kco42fZcPh4og0ZAc
OhdDaeG+AEcluJ26V8FXkCndM1baS2mXFMSl3M/srHdsz3fZf8MTTIN89FueNnlhJXPY9VpoWF9n
0vljgBt2qkUv1BqWxYtKH8qPmzQGsSgHXbGH3UvahcQq2+QxAE+JGR1HwOljrbzzeF4JcCRx2bvn
tttJfOkBMRBMbaKPUFD2CGwua0yPeL+uMbI6qnWCe7JgYwofYQcCdlvnOawzZmfYktgwBEulnpe7
0Pw0c9zncet7xsQgmf+a4ArRmrTzWxR8lC4K+fJm/rPT8x+lCsyQsoXlrXrb9CCrWrdJIfjIlx6o
EWQUUxal0AK+UaueEz2JrRQRLNj9JaZJvKJsgC1QmsYy7jr+b8mEUPpKrGPPrxMwbxLT07PBGrbU
tqbTIkfWSryMf9WIgciTvu2ds5rpu0JMBa+JLNBZH+YPzQCOeZTpQFz/rOWVNuyl/YzYdMNfm8sZ
oNOQ1TBKRXdFFPPyLI/V3RuAyXe6fkzW5urT38hkvFQF3T4AhI8OmAV79C35gdgmgxcCB/aEiEbI
V8yj6FEGhZGOFsI50MP0id/BeM85aOQs0QnauTjugrtIXxGSqzCevvnv/gL7Ejn67z3ah4nQFFhA
g5qLBs69x0tuH5xvtaIIIpWwFt5BqXEdyeOHlxzSDCs3BLydasHDClLLWQ35j9Shg5sv9Inrb3yv
7kCGFh9LkpkKC7b6eCRm8eeBNjXgkeasm7Nkbq/k9Ld3Y2Oip/OsGxPjHxcJ1jF0huHxjp/zRARv
8538e23ZgybDMc9uykgEiebFJ1iMVrF3ho3tzkPAKmyRfG2JcE7A8PyyXf9k7Gp+EylzpZKdMu2t
yxUuKkEIMhtTy0I3WsCx1vPsEE2OoP7yUlgLzoknxNcRDXZ31R0Q6cIsNzcK8Ld2aiEzHuiDAO1i
RBjIpj4ET2xlyw+EBFhVSb5kJVsAz+g1i4J+RIunPazckrqwizWNok77HJihHXlTMxFr6EiKwdhS
Eetq9l0QYuB0KkJdd7T5pKyNwtjRR3WoncIaz8tsXyWC6IeNapySIi8mjmDi4Jf7j/bz9ps4s8lg
VcIQ4tmDXnrktYz/T8SxKTTbgUovfnzqt1jV9W6zs30TZQJUqsog+vAMBDa2KWmqgsWRYVakO2+J
tvwouLOU4X8u/3gBrZOsLNwg0VXNoMEi0Py+VF0w2bwlSgYkOaUw6WJfQM85KZtPGkfr5mFcU1wE
zciA7+Wk7ofClGJfJCicDomJ5S4SumGDtgo08KOklaTgiYZpNGA30YnBmCLg3anxlnHgaX7CnH5I
W77+flYxYG2XG+4CwAyCHAOa07bAbNsyv94Sc5Qm/nyQwetMLLlz13v6a8T2OvyUf9IXW/fXXEFj
szaWr30tjGm2PoWBToMPz/onCuBqW0XjWMZZtroYUIrjR/le0kl4bFAjfAkOmMxWz0+09Zg2pMWP
7DLRvRO7zZT/b2VmArs+ULpTJFLwkrQRQJ6ORpRdfVbXcH4LauCJc9CTsouKR1jYv+5mbNpGb2yF
SpS79z+lBkp3k3q6NaAC73p5D/G13/JbwweUZ10g0j5+Fp91RRGL/a8+oHffCILJe80u6WJUxagr
yndKkidqA97Gj5ndRW35rCgXLIsjpJalVCFQuNOnHRzo6pxHyzyUpNlyA7obymp2BEYlbmi8nJ5z
pdj+Z92HCq/c5P0njeq4vg+1D/i1WgDegWb0yfyoUNX/dkQCsE4E7xA5gZcFs6g/0D+k0WlrgyO+
f71B/sa8DC37aWwvrFSyTzJhuv3A1wkeaXNo9WE+MclKixV+5PcmAfjqEvjgHviQyVehZpXIygcp
nrj+ZHYqQJEWmy/UodN8ijaWgTxW9wNyVYtq279lwkzM7VmTcDotPtIcTOPtCOxrBmX1m30KCXD/
6GlGr09rvyQuh226jCQ7WxITBEXyqp0fzYjAEDn4ryE2HWgEa2FNAHGO8+bNd7H8I0YE7csoRZ+w
cIUvR4OqGXefYGN87BacvzNbHjYOwCIsF8HHgj3vZInzWHYhXkUdQgSLMknxM5agU7icl6DttsrQ
c3t3WrjCfYJp3osqxjYDcS5bf1pb2zgCJ28TBmGVg+TXU/IWR+nPuMgygdhPlrpG0vqwA4Cw3ZoN
Wq2Pt/saa5Kkujif3EzMFJHDpiui5rrwJTYNRCNThwexY/Ia+rD5H/kAvdFnPrh/AcWSfQ4gc2sm
a4CFIJLb4wGB1VAONobB4ZbepwrwW+Wh6UpHKf0s1u5P26D3W8IGjbLNWk691GqrFgaNytpv78aJ
lTHJdwsISqOf0soui89IFbOUTI3yHCC9M0n0w24xS4ga1GHDVpPxPGtfzFk0et6hokJaEC6jfjnT
nGwFwHLMiQChKGqhnWtSvONi0AnKcPI53tF2PlyuIv1dIG54rmJYCfmrFvp+t/SQeHFFVqo8yy8g
05eLsm7IPMhAmN6kVuY0rWZBiZcbUfblBf6eTzOsiN2pdPKjzFRo80jJWUvZOtMzFyh0VFbhuXXd
oQe8F/jcT3+3QkZHPyLJXgvlYSZgjJHSojiOrLqhLtTlCAzbLXI7aiuJjNRjGkLDoDKbG761iG2Z
IA8OGwDpg/QH6yIO9sR4lkHxK7AZg9Qr7x6T/fBl8z9rtpocmdvo8V0MV2ULplB/al2okSR3g5qE
w2SHYc4OMYAp840cIL20NZtlmgZY7medDU1WQ12a+3TGn8KHXceE7RKZTmCuJvhhA4aW+EnEaktN
PHT7xXE6c6koBdC6E4RppiUymZi4+9658NECt7l+BmA9e7pEYQgtS2T7eCfTZtQTyHdZoDz28f2B
X5CtAyWrlHsPyKuJz+6qzWnnPUIV0YcBlmvGwZki/NV/ez6mTVBqThZ547vSsPvMsYgJRrP7qSWQ
FgAx154OvhKVNkPfx0ggNUEHqd3ve1XD4SlCDUP8sHyIDQk/URY6pbhwaPO3IEdZ3fEN/hBMdtes
qe4rs6/WOwNRGsDHVLd1LpS3h3vJE1mXOyFMsnmnmQAXpG86juhCjIjg4fkOciLkkQ2rZMErWFWK
K5wUKY6vuWwkRoul2FsaK8D7nrWq3G7q5TEVMdV5zl0S/eA1aqxRk7plo/BW9A5SYhFm2Byj26Ht
TL//XydIF/zfc8tExoqVdR+z4dQouq2lHqpYyE9qCO6/RmvaC1hEAqm343CEjCF/oXlfMO0SNsC9
nJOvEWxsBd6P4b6uIx+4Y0SXNPMxo8ezGXg0DpLdnSw7Hac3GrjRTFGyncLu49GSXcWzJu/S89Nd
7hhwWeYPOLn91KgPaRhz2Pk1TX/RElvSulTEwWekcMdqCoUSTYbCX+iinD47cKEBrTcLLbhaPArX
9qRXUaHo2zOckZQpeis9Cst6QUewHu6AeqWxwCI7KPWNkFjXAVDXrzfT+J0nFyF6ir0ZGuiOhN0x
bmuMFCBrUCO2hnJRsPDlSachEk/VMOGEjb+UfSkI0g3Xb9839Tnr0E4UVklgkpMZgO4psZB8Zyqt
b9fFt5bz3K7jR6/jkRLYlcbF1RmctQvyZs1OpyfBl4LDNBcJGtCDo/xt4WHh8IOGupSsU8ZeP9XD
BDnsZKX1N5sme207pVhrl2tdtoesXJxb4E8joVO5R5TIgWdUXXfN1OD10SIssWOJab7Pr/yeyPgu
WfVnOdA/KMAD9GviaXJmL/3oqJrv6cwSlWaPTvNnA++qt7vxSV4sAlVmjVmiD8MLehbsv6JIm4Ka
TNyC7qeJZUeJPkigWbhzeiGJw3sEP5e33hUFY/M+ommwC1dquQL6+y4VXksJrUt9AjkGQDTlxmuN
eO6qafbvjmNQ76FBqN8aBDJDQK9EV220wFoLVpLL3Rc4WHO32gZDJm7XmjwWFaYD707vmSGQaL/j
teAWxA+wZWh/fzjZOnR+1zE8UCy7RtIcy7N4IJ4IF30yIv70lBf4ZMjgaxiQBtXXZ8js9KD+TuXT
F2gOJ4StzlQbPvOtVO6GOwZvqxJZa+aq9irJbdK+QvYhID6Zz0EWDHzn5i+qIts3gdZXHhziOO8n
v86g06mMt8KyEbTmH6KiNZmqesNb9SyiaW+rknj+FwNpRhK+t3qnN6wTOid98e0/3WFSNycJqRKr
+O8c2lO0vUm7Ws5GmVk5Yt8D8ZrlUwdgI85UkZstuya4NCugEpSnZYSIVOTI9SZTVrJe3YO5qg+j
hsdx3Mu9vRFU5bJlvB6gBp9uKzT+GA/6RScntlbijVNrgwpbbO1v8g61i4ileXViuDGpcPpjE+LE
cUD+v8WanbYONzl2jEclai1JIIOoKeETELHPDCxMJecmkF19ef5AGPLoJSY+VhPCzq3EDTBRcQcc
CZk8P09SR+iRDnXLtqEqT9b0/3UN0joVxrjZlniFmauEjd6ey8WWXttNcBbxtB4DNCvHjBB+tDkU
GurnVtGzMXysO3QINvh3VaTu2jO803pQllADa/ZDXKVevRDmiSJRYgTRV5UBRmsQvG0UNuLkepfg
VPA4A2Eropta3vM9K1c4yh5zXIR8dmG94dROyvJFekya+JZbn95c4ka8Ubl83QuURlE+P/xT1r0Q
0OTh9mP1WOGd3lkj4gxXUGVpoCwzHMRcOGxV8zHpSi6oDjky5WveGJ/nhynUgD6v4SJpJ9W+Zz8i
HL+BTlFO/lDQYRPH59OytEml+0I/DyDWw1s+G4lGpg1xa0yYL+KifdP0YcxL24Z2QYSpzzYCCBel
aES4RqdXvp2VTDyteD/6r6jQtOYkX/FVoCzNRn+F0nmgdemYM4FCZZ96jKxKVqKpcCuTALsS1zZC
WlhFd5ogIqjdRJzgo9jrs4OPCN3sRg+OYZKdsqY+EHBy3oGRaYi01fRZpy/lcdpXwNQQXgFQjCyr
rX6Ii95/kIQc5jTPHba0BbENeR90XoLG5WhpjGgsKb5IraqrPUAUzH8e3ZaMfwji9jRka3Skmvio
gCTrDAk9bRtgqrRc5gLakpbI2ejDcoZGQqX9lK+IQ3o6gi+jLWy8ZC9azky04/wo92g8a2RpF6et
Rfk4Q1fvSKohVY3j4x4HwCb8eG/k26WjPwnjvXFOMkIO7evG51TsZTeOilN2V4edZuOI/4Sj2EMy
aRW1gykJjTgVOHrcUpyy24FXPN3fZr944XlydAg4hs3H0LJAQ8LRc98kcT7XaR+9hL3SdI4zQzIV
DGIdXZWR7viXtLmP/kiR6Zdez8UywUlH8N4WcK9upinyRtIb9khYSDSmUDEKHgimbekdAmJNNxT7
IypEQPwFDUVDu/iAlSuaCEzOq7Zn2dgEbV6tXph2WrhJ2C+YpvJRnBdTdRHcyCuV646HoKaQFaUl
hNqF2Gv/Uvr8/RyDy3h9xG/XD0bEXqSSB5Ut+SlIOwN+KiDfyeywcfQDnYnMvoSmVR4GJNGyiJwh
o5X2aUDNZGiphswjfHooukrt6mK7rNF4y+GudklEBxiCQCroru5RYL4oW+GkkmEs9claSao9BqNI
hwlhZKabCt1AZQEZnRwMMhGO292oLL7s0dPZoO/G+LhCR7lqlTntJ/r5e0WPIdX8HT9bk3mSVFDq
GMET2cfq9uuQZnCaAbrduTF8ohFAjSApTOlrWy9a44C4+uXHsV6XkuYiC+EmluyaZOeg2nX81Ogg
VWOmyRR33iLFYQjQrNmBO3p3zbGfBISs3jhFUvuqsVI+Pawi/MulqlhE2DAzQCIsb06BmoLPdcmj
Lw69IJp6u5gykmNS+G54b+R+SsqfPKnEQFMElU+VUcsG4jIOQekn2UotN4XPCnuLU7OE3RnQxk07
SBizTwTqn3qjyxUQspIJxPHyWy/B5B3/PNdbEYbcEge6OSn//7thOps4RtI1cF1WsoyyNj6qvRL0
tjnTLSAIdUry7yRXT3Xn2B3HqE6SttGB0/thnMJN8HIDqHe16PQwz3N1ddKZ3+Jiq3keIctFHeIF
yn1ZmA91LGKnl4V+3tdk554ZOy2tv+TrueaAovQeGxxJqp3Ee+fVI9mpUatUY5/hJGGNKaPU6ZNq
VqMOaK5tlaNn6q8Dp2CQ2pmfBdlOiiFEnPaFodoOIXyKygSZ2Oxja5uBBprURTxXJk8pbqGq8+G1
u1ew7Bl9O3nzLbDFfn6tgVvhwf+R3EMC/U+qcoIsWb9RUmbLTxcCH8Kb9Jlbf4GIiLJ9FbBjz1x5
whYTr1Frsss08+L0RJ5E+R2XMskTffNk07kL3xany3lMItmuV07WcHM7XWMN/o35MVoFjJrZAa1L
mVBINriUcZ7+OqwZUzS4mWAYH19IUh2AYvyLzjbQbh17OVktp9rfzbM175Gyt1uNgCSZVMHV5bvM
DEm9PEAGcB5xKgtHwkJ1IXGxgRKbimSOed5TEijjLsklykIXqMLBz5Urd7QXz25wQAuiaq36K0mC
J0h2d6AnAF4ezWlGEkP5RHoEZ9rLqGRVDIcflTNzEtddKE1QIiYf+U8iiUL5bT7RN3Zx/hVv3nn1
iZbhd0uU3gHyaovPWvPt/cX6T1t6OOzvRhXa0jDMwllv7iTyavMmGel+ARRu9i969WCUa6S7cRNN
z7NEb34n2ikMbpugjdDQM+EAMaXDRN74avSH2T/hGyhirceI8maq/aIAL+y/SCZMps20VyIEl5Lg
hI8hCuZO5TU+OO9iOoXvmSAT2DMc/UELK7jBHA+28nDtqVzlUVft2mPM2UTGrtK0lUQGJVUNOcs1
JjhF9Cn6SCrzwMJg6KYrlWSVIRiBKBFF5v7Vf2Q66W4f2nPo97Hew7S8wM+CAOyWJN9+MbLOWyu4
02aAZtkWM/uKBDPtGTmMG4Fb5N9lOB6nCYcjNNfV2OYc52iLLLN9wRLPzhq7rLJbEGYxUhiZd87V
5+92XZykY9YCiwzEyKgindzpNdjIxSKj199OrV5btH6FRLTFM8T8gamwXB02IvwHZUPT4Ih1ZM7d
7F8kU55OggX5NjP1rR14SCPbTqGVMKP1Z70M/8QMEMbXQqaOvxT4VwLPvFPwDvHaw7lwxkCvWIWf
ttEth9M2gsoL6RCXlnjLlWQce02NiOnGgtstBehCe04WfvMBceTddy5W4CPtKd4iQXBZU5tHdDaX
88bQEOdNwFw+KZZxR0v1CNfmt8Pz2zyih/CgL5ubMbQ1b809AzCN9aFz394AjPvB0iJ6QHyYg3/Z
rZKLkU6j3+A4vxMbJbJpuLiPz4M5EF1KGFXLuzNGJx3gVETYRF6gKgT88D05HblsLMksMg99noRt
1x1vjuhKaDylnSILe6TfdYx1LVQ97yGfk0gZtHYW2/e9S+zlfXQK6uLbQru/brNZlxpSXf+cO0Em
6ehXUCAa0xzv8DMMue6qZjGgXPZiYZzJs8cQ0rcof1cWAZFrXi2DA9TEnQ33ZXPiA/0AjzfyTPXL
LmC+C56icDC1XQp6NOTp0rJCettpGbkQFXopRLab+kK/4MBO3uCeNJ86K8sRKOqK3YBc/jUnHSQN
oAb0Q06wp3/OdczgYdnRtXKJ2MidkxsdFOL4eKYS/9bwAU9DglPuox6L9j/VjHc8sAbk6A72j7Al
nh4o46zCTbHoV44HBRm6Yqy+wmxEwKBO6rIyy59TCRgz75NW595Mek34gWNzEOapdPfvK99vyW9j
zisk12kfZsh6EdDX860Suba+Q9U8y3MEHkqKMLDonFgh13UraJgm8F9NlGbgH3KQ9I3IvZ0rG5BV
cKEikg9yqqOB88qSsE8j4+SsIxHtZqvQz0+rrh5J5eJuufZ3eavc08N8rlE31MDob+JoUhTRzdIW
7H9Njf+3dMkzCbTcaIlpfj5TEcAUNX1Yp5Jima9h4+lxl8M0/3XC8RCWdlt2YDgfkF/TiVdwjuWW
cV09W3QbXHa4So8EKv2X90FXLgAwdM2ucfSZkjIajGZFI+uLXsXx79kWtXfkD97ba68o5hqV2iPq
b7Hzl8Ph6z1mOoZWwgnb6VmOtM3lOx5WJ6XY7l/8OdMLF+kMZ0lZ163grzCNQkTredfaAHfkyYeo
FHpP1QyL7wnmOCFXM1mfDjLPUwhXSG2dzFC/2X0UWwuLR7ZJiBLfMq7j66bZIfopnxc9+0mw+GkC
Z/Fwg7D59ZHmx6cXDvI2CeKSNsJ/bdz4DgJNW9+Lbr9XI0mTPViwYha9QfoZ0Z/sEecC4QRf7mcJ
z7H/lWKmMWsKPrq0m2bl5dAQvmdTc8+gInGCBRUpIgtOfUNeUkYnfVzXfPOtOHbJ99Gi3FwKsDOl
YfBJq18Ggindn0BI1ce55cOQIFshnJAwrOv56MzdvAsKa8E4EePnRkTiHR0d8WHCYgfgeaNOvDVM
qL6S6JjwPdYUEVfOYH6MOUJ/vR/EtzQtXvN/JZC1uI3CPXxnlopwRBy5peQphu+mX4oiYtguN1ga
b/n2uZfxp+tqYnyBYaSxXy5IzEDYWhl1WUldleFJ688l++KB0RRTI2mueF05ndbk8cLEQOSjLSZg
4Zkq9MCsKXgr70IAY68SWcq8ndMMuhOfAeKfwRUr2MVpuZ3sgpbXGveF7wIWxj2XgMEH/NUZif/a
IloQ1mTPOkQG4Jd90lHERwBQ11p6SNyKJ49ysfx0R4zoGET5jsA7zu9IzMJh+6lsZlzEU3Q1a21T
Izv8juHr9oBu3KUyBtu/8Szk4dPU9oWQtsXXRkMSvsOP0Sp02jnLgVAAmRsCUPcBvvYq6qX33lgQ
IrRyHPhyOKfQnSxlcmFfvyZnYFzFTXL8VjNLmXwTkTwXIlATHRhgdKvpUGkxkaWo6LQr6eYDJCKy
MEmY/sSeFs0Z+zZ0kn7/Y6zAVDtK7ET7nnzTUZ7EaDQ9lWDkHUWKEOWZOWSdjOpVP+78HG3BimZF
90QehZ1e58SQxhIL43HKkxKO9mtZf12nYZelLfnBNWUK0PuHbFICAy2NyBSUayqhmuDx2rXnXHYM
gXaay57qU91GrGwyrKDCTQ4Q2PzXLqkPm8ZtE8FiKUOOOHakjIgDa5yJnDn8kKWvSYWLfXhhHHAo
yeFwdbvOTUjILGnok+XS1qvyZoTGfRP4vm4ZbNRJei3FQCb/rPBZvnlN5HxbvwXrSV7Y1/qL36xA
g483LQv9+C0soIY1aDIn/M6/lubjkeQIEI7krB0E/gX22gm5WqZPw5Hv3KegSpQ/jbpARV9ciqJo
yszEAMFyYwLq0oUEpkVzLgVzNb6ZikXg5LYRa/sEUjgX4gHr59u0LCYbqUQ+lPUzcydKY6Qla7D9
2RozlHF/RtnK3LybSbrf+7dyHfHUaA8L0FG0vh8kzYTtVLFJBgtZ8a/F+qCXlpz2JOYarplEe7xq
ZFHhAa/qikLA2NhtJIANOCuHqEOEgYQzhQ83hbsT+AK8MNGe2T8j88iZ+P2CC3tbFKTX1Yp9Gz7H
zuvoozT1bY6BxNZAaqqN9wFnNPKNUhJBG9MPoe/ID6sbXMOZD6oEdd0tCDBvyyvPclxzqD6lbPoR
xBB/5CMPyJIc1eyMmMgPLS+hDTkJXncV0Wliwa4PNVL6YfsgdK9ul21rsvvQiMZ3BWNhXfMR8pn/
0sci8wjqPpyHZeTMRDxTPoYAEgZ1D9Q1f9oNs7a0Q6FvfZGu0JueWlYssnSgUaEb+ofrdwP7SRww
r6tOtLklf6CXbimK3Ib4f2XdeXB+g3t79ycPfwLr7KV5O4PBYi84pgskpahEgGo5Vb6XYqIX814W
1q+UvOZvC924gQKMLWIkTQMH9o9EPvo4oQ4XhawnuSHQKPXbytRvLwzBK1VPyqRP1/XZXkXCpD2Z
2fzFB+yy24XbwipGVgfjqO31+y4rsL2k9yjl2vyzXzWkT29ANyqrbcd/Musohsu/ImujyRZ0R1qm
Dm1gEHRWlvlLlcrG+Px7g03pdLx8TmFlH83rhxJuZRLgdDbXBSEzX2Y3AYQEkFh38hThQIj+DOfk
+h/wajBzn9OPws5lH1wql14RnJNLj5o+NBq0SOkqaEFLpAWkXDangOobBL1TkGY/SfNy4uCa9I8i
6cqVOdKaq48cM5DzcVQhFflS+m6MibGliwVuLdw5KpZRJDHl84hvjWKhSbc7zpQ2J59dcnoq/4HC
a0qVFRiE0UveganUCvba/f838ivzhaUfmXQSbzrJ3FNLTdfnllkEmuQoBys7ANAskSrVKkd345k3
uN/+c/7QcgwUvb+Ztso+V2GcMQi8mdjhRSGyfAYidBsvAY8owYGlruPnrkBsuOxlHEPEKRpjlcbw
iNw9GpdZkw8ZEdffMF6zJ1x+HM1MJ1S3RLfo/XPTtGYEcpNOH2kAsO62Cd2Ul9xwJBtUQSJ+xqKy
A8W0bvm/Iwk7+Jk92tmaCXvzMzA1Xcr5d0Y29chFH22bZugCjkAdRTY+RD6M3DG9P6x2o5QK8OiC
rW745dKvrCtwjSweb5zMUbQwlKFR8hGxi9mWXtJnqGp7a4j01yQ6SUhvpBbLXm1IR7jFj1YWnPet
lTXX+/mvE61wyFFFv7N9tVu8DxCU/2mKA3g+ozqo87EZbifZd5b/1Iki17pI5craWPa9GehV/Fkn
slvsNSbG9WOuuMlPCEglZI+kednmQJUQ+/B4fTn8iVlmhvIrDMYvn7bnSj+pJnaliv8dFUkrswMp
ybX2o7A1PiMxctDqbUypUmXzoivQiefCrY/cCrVBah+m/UeWehgiQKu9Lop0XQgd3WpL+VGEMewt
MIBOask7CHK0fDARs+Z2kulRkzct7g9N/K3t6z4LagSNp9mSbMtRuD0BGOfqopGut0KAEeOXSLW6
YhAsLuGty72d19ba+YMDEqFHsHQbmow6AaN4iTgAUOfa916jCxWgTtfJI9bvsqQKX7HTwT3kyFjq
XvSotJXozsXb2I2DMBA1KD2LfE9yCDutH6F8C5pul56wv7PV2qctZgHsBBrilTcl88DcdHWpviaJ
B96YHBLa115p+FRn1LhQCaa5wpSlvS9suwOvHjUfDsVp4xGWp4Nwtlymz2xQzhFHatCQQarV+kRi
1/Nj5bHOSR5+yF/LprjsGm05irwhEO70cRbw/JFync1gPq0LKtFkhgk5JqJqKuiVJik5OBHIxbQH
Js04sJpaZdHotiTN87kIVAOWx6Rq02sWdCZY6EAJWPt6HIZ614/CFK3or/iPD95wzWhsj4ivvG4d
yo7u03Wvk6w/uN08eSu1Du09ukX575XmeMwy1DxAeU2Xjis6TxFdak/oWGckddJNMeIIFJrppUkF
13jQAoOqKql3X2BoIQQ/hnZI0anmKijU4jlG4675/ni4QCoHVaxpoNSZlNCgsxHkZrFl8XUtq9HV
+y1nwVIfsT94/RrpCTt8YFJJ7QXAyTzuyeihjHcPSCqSGRks97CUiQVpRuIbMs/5oithwXcrhkP/
EEwHUCEYVqVyKTI4cb98gSAMtHLrAjyHyKIJ7050Loq66l/JGaVEFBArtF/i0sKbRXZEDBgYTf4e
llHNMhHnSvAjjXQP7Ug6898oCfCPHr2wuCgPJaWLxEmNFloztRi328zyIezZ9vxr2ib7oUCMNhLx
qHT5Z6pML1eyFxBF1VszggRNAu4R1Gl/VlJn79/vtPOnndLofgQf4HXSUqtnpY8M77TCCdJmnHSs
Hs56C+Dll1glioESHf2XpJ+cBnj6acY+NKSboL1OrqtKgjMXK3KmnpQ/JK3Irrd8yjY1TgNjaQsE
iyCguIRE0Qy9QBR/zSZdgNGblCLUK4dQGaNvKx5ocLdV8xvjHmRkLKUJvmFDXdcscyWQBEGc5E9/
jrze/UR4RNYBhRclzXNRaFTE3CwmrvPfZzgVrX5PgXzyUoPifDJXAdGQ+19tFxhUtxSP9YotIZ1E
HWf+9DKhwQedFhIDS4QL90o6ky/VIe+qux7b/0ZNLuNrtpINrUFeg2GGT2wk/Ow6VMCedIRr1ml0
1tWnaQ+gn+JoVPpM4ZOJnhJpGvulGYaKQYQ5qu4qXHvjl2NeskDVJB3r6p2IQYiE1eQSuejadT/D
YRQR/aCiZIZBRMTEL/Kw8edpfToXDtXj2vF12cwVQ6L96wOQEf03KdDg5HzJHgM/VRiruLoOSB4Z
DeNMzQIVeOALpZxZSxqU92IuZWGg79xhn+ME4HJFaoeq9fgYSUMrj8hJPFVW0F3CZ8PK/MJqDTGw
0q1jHPvnqz5vGoKtu9KkoEmW7AKAlQ9zwQk3dpNSzDZMm6E/9EFPSgQqn4yFn2mqVm0hSy2KQGrd
vKqlh1A1zXSb6jD2iF6lRwq2hy9bBD6hQD+yQ2kTQEFcOcW4JhI9ZThSeBfIldMor9oK1L46eeP3
5/LDAMVswyuQOmO/8mRQrk3KGWAGhIVXRujDqyC9ICAQGNdlWoyDq+/4JRxU0ORwnzE1L45ybbr4
4Mz2xntjhBpK0L+7Zeeh8GrJnhk9KNflEy7e6JdwspW7O/rfecDUj+Ic+EQLSvOPnz6kC1ErdF6l
d9NcJsAoO9jLzNVK+Sc4BHplMphDNq7AvIp5LkCvTr/mtqjFruEifcObvbxLYHGqi7AjXsXMQCML
RGtmuSFh+xkjoVjHbTsSjy4LbQTOAkOTmfNmJZe49KFBrqYSshW/ZTY6KTZAOXeIQ+EfitUbA4wY
Z33fM2oUx3AxeHRQxJFc/myqdF9p6nLZkgBbRSqbJLIJO3o5oHfDRQWKRchQizfzuvn1VHGbY/kV
+F+onD9lQ2dGspzwXwEDQNc576KT12OVOhWPmeP1bZNkB/GfhCJojuF0E2j0Bh7kA4MtYmytleYL
QSGVI7l/XfoRSTMVetDWJVbxssQ5Y/a2Q4ihR4ReVueuzZkQhsuKjN/atarDsxxbeywhK/l4QbnH
ma+CWI3un9BxfZ4XVW0kXm5Dev4yDmjEZOhGIxMm0+00M/mijhpaDl3jsybr1EnIeXUCJT0eH0Ko
UTW+f9U0pcV2J8lfXtWSewJ3DTEcQPKAUoqpFARJgY4m4KI68EkoCUtUaGQfIaz6gPrAhA8Numr0
zDB83TSyG/613GmNfAiYjZTz40qmR2P8dO+UHgHny+yvbc4hpyyfcssEUYGjuEluWrlY9eiK5i6W
9R7CdCW2frnsjoSKJXZExlmy31Cj5WxzlNT3oAFVUX7UVAlaVxDV04JAvD56ZiSuitmajWf7t4Sz
5ZTyGr11mJgUiBRSANYsQw8xrV3cf3zuj4OLQycezYCN+y4XsYAGBFwDuCSYc4eA4pJWasrUEtQ1
7dWh6+OriXKsdZvcmcQiTLWDu/gcpV8l3hKk9V0y3ud6XwujpuuSf/Sux/09HoxbS1/Wq0camzCJ
wmFZiw23QwnZ/Ydu9wnhVZRUtcn8y5XSLU/Zf83JVj9j/8CESwLo8XenCVbgsSJtifZkVXruyvXK
lF9VY04IGs7MHOcuADLO2D/Fo2oG/aY/VWDBq7jhmflMiFTbX8keARfHy3WzqoKYa5hU1DbnvBAY
tuiirXTZqpPu2T2kghHKN/YclBJ3mELGN7NTgswunsDp1Cb1M9Ky2GlVcKWzwO9VEKfjyUz+FwJZ
bX+tRcAlxBeljAEZl521UibQ36CW7nCNFRE4pVvQfJUuCP+jmxYhK5KpZ1tBY8y3FaK5N4YYSBM9
pV/dymWKwWNCRg7GHprCGTHmKzHmuq88+SoMFJE83DigBNTnssQpQT4JUA9QY7QUbR97PKXJzKQ5
2EAA0RddGlYyb7S9Mqd0vKEQ0Vr/e2rVdw+DTojN1mh0QP9mpvvd1a5xsgxwkXAzjXJvJH0Kqct2
8c8gwEyzhhaW6uo1UyT6oAoijQmy88Ln8BwFt3NsTACezGWMpwLmeakDxu2QoXG2GBRgemfZZSMX
Ot7LWNuprbhMdtPGmFyf8Sp7UEJgPE2iJIqX/vhv+407jl9ujTlqiDyqGAvhXadSzYr84TSPQqu3
HDPQGtTuWnLy1gHW1vS8I0fuHFNMs3KlmATWKYP3rgeokKLLytreffFugkEq9d5cZTu+IzCle2ii
yvGujY3TT+OOKe4GlSS3RuZxtP7jDOWHE93F9+AejWgUKU7l6Nq7SFRaDw6NcWokUjrS3ixacTj/
lbJ5xiNCWTbCcyKqfeNUHUJQTe7iOHKUVWIsxY1E0SZtG6ZJ/QbufzzFXoOqKkZl2GG5hKjA5u7A
RXCKEPCmAt6ylHLbJsXG7v0lD95jkFlKDelbf9isf+h3AKNS4lzCSqeQn0QYUmiK1LJ4O/qMEZdB
p+SLyQpz3CmjuRtV0f8CEPoH3y8yv7zjrmPvB9aCepNGod2nRasxjz0H7Mv8kCB6zD0cqpTzyK57
v04RYrUX+YcuPpMq+e/lQBmHs8qLX57WjQzm98EjrDRdP/IfDD4VzCgU9zxx8H+Kgq0npOcA6ydc
HML3e1R47nRVSk2AgdaIqnyc05acmLMNdx3VB7B8rqCKCoCR+8H6dBBRcDq2XsNv1RCNcPUp+CY9
lFMJkYcudr4QwXG1OVXY6Lg7xJSZUIXMtESF5D8+in1qL01aC6E0EGVhFVIWY5ggj8ekS/GbcQlm
9XSdM+NlnVwNze+5kdYJ75uEbm4dqcayET2TgkSt4mo9i/K3aavdOjbiwI77PbON293cVOPA3DTS
TFit0yNJ5lQ+ADg4PHIeqVxaScS1JuVo/E+wt4mFAXt2pEfhkulhoQDg0rwbET03gvA8nhhZBZO9
7jQTV0HbBx2y7L3ywtfJtApKB9BUyM5Dir6M6KB2vZT78o3bkyRtlJp+0yiheodRvLfYjCABP504
8SKC3O3Bz9t9/V52p4w0DSValSbQIsQIopg4gglJ6KlxBoxMHf+Dsha/YhrVy/GHgaOtH0NYPSfz
Yityu3Qju+FVxK0ltLOk3Q2uz6+chHOBdvV8n++8kAQeUadAuuibS5bkfwBS1Upx5B6w4MoaDsdV
Epm/yCDOLf2zEfIzMpPHoLLHLDzkxSeFNDn6Hkqmv3cXRnXFs1YYrdLwEQXrHkjiVT9NfI/iNVO7
MyOtIyua4wuTtTMYqXy35nemUOe3PAAdXmaHSEmXts/TbIA0q0l6JEvrrBVe7f4DZxO3NdbLmZKm
kLI31/YGOhxaZGj2k1QWp3+V+R5BCxZZNxRakDFHZyOkpUaAru7fa90wYvYntHp579brEgegvHer
duvlUjzcNX5OHVRQ2c/o9qlcAcE1dmbRp29zvBzsFMErayXgRTKvAmYsMTlTXnkhGuJfJb9d8hNQ
KtS8eKDi2m90eCQC5nvPIm7OdbNOqXwqdZ7maOupfPC5LbdPriKPnbIRQbdPa83bZ98cc/jJX1Y4
juou0FVbWpelrOrekyBG/XLj2tuQ6V/kESOd0l0e2odi5X361nUhs93SWaZWrP0HZ628ZO4tDQOx
B8KU/khcSrnS3rS/vMu7Zvi4oYLFoLIGnejTJQdnoAfVfcK9TkkiBXovcJJYQ1K+3qzf0/+AC3bd
s1orblx25o9wGWQ1ZFCG/Cfd12fqEqdDEOvJpnJzvzIsxYXvQhYiYmRpk1porr8LBXpE3O8MTbxx
apQaxUjixEKZ2x3D82AcBNNeJ6ZPHTZp3nEk66A4SSk+RJPi0q5gttbhMjslXqHcrE0FDkPzxKjV
+GA575Gaq2dFH1OlgU17jyWHdBa4HWoZlQ1Qo9QdvMtdbRJCVAPNHCwAsEK/a4ySfcUrvaEtxpKA
A9JQ2g2TkmE6LfkDim6T+4iMY1PHXZcd7gaAVvyMja5kumsnOcx+1eMdDlywINk8E6T0YVfv2qJ0
g+3Eq77OKGDtyjXhRVX8Kb9PFr/UIegtoQR6PnOT0uxlQXFm5tuciM80wF+bnun5uKncM9d6nu3i
Od1v8so1O2s/0Q0cQnK3CY6i7IqYvl+8PwFOirwiMoSLv57q8v3bZ9pHnc+/G7F9WPlaoSa6+Uzx
H+leheQEr6BY82r+CMPd1JrJZBnh19FVhh4R1sBpGS03RjWuLBDT73XWJwZk8tc+w31umduxolsa
cud1Lxrflzln3j96mn8I/S2XoEtEWaNwXk9bN+EPqvoctuUBCmxw8K9h8DE8Pn8kapkVDgxkJ+M8
3G0JY9+BkRfUMBVdl3OiCwrsRxz/mIDqegp7/s5dGOQsy8FW76je05IJZ3NDTm1Hj+eUpX1EQVyT
EpqZzC6HGGE4KHl2ISAxXjdE1Zv1ViqBJ57FMCMN2BVuuQPwv/7oFnlOHWiR6D4Z0U7HgwxFo6u5
o3hXxjAsYBYDy0aZC+YBGMLQPTGIVht2iokKcdz5uo4+pnKqZj9QCkXkLwb75QIgOy+vHKH/joca
KUxUmncicEH/CDbVtit8Q7PnIoej6CD/CZJWYjGRSIjLoMybBMtwrA4jPrSLH4qN85Qoj44S4dFY
wsRQHiSOUELv/4nGWSjUr1hUqHOxWuH2mtLfIMkY0vL+KyQXerSQrtBeyI5QI3nmQKZw1sEGyIc3
Mx+MoiHXwAYm9oOQQbI5cUoTi8au9BOYMuwydbWbtG2ATId7C62uXwFGr9kcI7UElYLSPzeVC1Oz
Z78n5MoNn98T/Hpcu4UhUncjTMhAJ+0uhNwEvSjVwYfkkbqaoQ+KcRYI2+ZidVohuNcN/M50OhIX
Y1xFNcUfRM+/iV/eBvR2nSO/3K40C9eanjZeuXNBI6PrbcAIY+OPt+W7hfuB8S82bxCwJieHxK/v
kFYSQ0SJwEeZXnGT22utesla2/ZX/LIdrd7EzMAYh39q84+koLEmw+sq0FxdQjR2F7kw5Xy9BU4F
/7Yom4qLNF0UcjyvLh8R5b3C1560xMcWlP8hqt7fp0iUDd8OSMWVkUPGGU4hXYQBGyy5vWVu6Uct
D4IBwh3qL0G68nD/ICVusHcWe7MlRr+pU5IDextsd2fmmwGZgfbxCTGfJL8ov6eYtLhQ+wS979lL
zQJfdEgVeedWaqz+OKc9mkbXSU9N6XMKqGqmPyJTZxIh7GrB+SZsRSPF40tyZ4MoiF/AVlQDy06C
sZUfD4mioSJq8rtoS8fR9LgctGojYY0I6YpAcr/h9ZEOb9cQXh9YQ5VUP6TM/yRxyw1fAJAFOi81
HJMxi9dNhlEm9cA3VXTdD0l7ZMc5hL9wLZzKOGFKKOC1U9KqERNqBqn00x3RjOj4y2hs1AQ12yAu
H75dQIrnephyU5yoCQfyFGPDe1hC4aNAahaKd4EeNI6Dc/47cytMHa0R6Ibc69w1gb/SbROViOYE
h3vwYsOk9V3KHRkh0raWft/j94EfxkCzKa0hwOFKcqaeRd+/TDzahrvZDfh0G5NFoFmY2XHfmWZO
8xvghBiMIGnmb1lPbHKmqJAwFiI176OFOgjgMsICMKGlloGFeMSQtfqOEC4qvQlF0yb8fesjc/TP
kUX55hPt+2yq0zdXzIOjp6MM1m5F17IEQUuVJvtNFppiNMEEqvGLhwXTTQxRjqW0jYuDK3p8FJ7N
4pvwLWXppkFiBA7v661LXwoXOJNe6mG+3CFhDw8s6fKOZMklSWAuTRPrAu8KpsBB2arAyR/PuU+G
KVH/3dmGfC3lZcrCMZGrfkcEstcFsa84CFv+2FZayZYh82IKvCL2BbJ/LKLTEZAh+CXVE6lWGr8d
+GIH3NZbmkM0zufz6fxrI8HAyDYhC/9d1393KhSdILAJ0gZ4svuqlv/ve4Y+cfz1w413Mc3T1bA/
tPOo6UGVLbCAbE6OBBJOYIrkwZTY8B5beJUWzPv9Y0ohSzPus09XC1ggdamnD97nPEBrt7iey1Mn
GopYnTLJIptXQ8x2MwBwL73bZBk7/SHQQyeHcCZxCsFtWsTJRgIFphflQWLhzsWEBB5AT0xrHjr4
VSV6dbBylpQM1rszMdfQutSayvinHFfDTCZ8H6Prxy4XoAunhzZsm8+T9zXYviNuoKaUAKWM0Vhr
6KCltLnUhOOQZ+sTvuOy81uISOimgGgeIy8DDak8Im7fzkCMvOsaoJ4q4OxqzST+I3v7bGDHsf4d
xuzKItgjci0Sin3Lur5cEZmfgg+I7Rt7N0s4dzpv5Zz7ovSop3uxd14T4SLJ7AJttuFPA+UUqjrL
h0cxA2bCiFW7ugNpV/belp16GMwrx6sWLKRRu57BMBJRG+AIO1arXW9BivBNyzL3TYmwkB9+08Yx
xu3vYLAjqRiEip6DH+YwsgLNr486slJB0kP6MuB+BnqPLPhxZbrMjg4VFXyQoGwzaH4gRXO0zww9
AJSq2R6n6rTwgOud2N4RgOCE22EJaW/1sYrl2YTEvxCvyaEUv/xo+BY9cP8JLrKZ+i/m9fj3rvQ9
TxyC6qpYgtO7Rrzro01PenCWPm+jeDmVnBM2p/uLeOcfcsPkKidWi1cA7JPk4a377IOgEOfhAIEi
c9kDNsmxcuvSA/q/CwNsmWNgXsvhOAdMWbTzpt3I/nrTsu2YTNGzTX3beXJg0Ea85ZwZS/z0nZQP
tayEERfz/t2hP/NJGFQwB4hKXGkItj4mnZnhFmdWcSL8DULHJ1Zc5V4Opuhv8+RcYPO/Zhrf6BBT
2AjZOiNFaVKuu2AGdZfe8GQ+QL/fPkD+OIfPuuiK8v4q++sIJKZEMUHfLqVjCSuRbssSMQMSudKp
xgIsPQABIAMB4abliPe7CaK4L0v1egfZu0Mh2lEs8k4TRf7l30F0REYR31lv2kUTlv/MKRBTy61Y
wo2eN30U1o+sTh306hslIUihGOglq02ixOX629S+k6x6Z790GWcklNh51zBCOCAvnYEaQHs2QfTD
L6XVjyS1eiosoFvgQalnUWt3ItRyHDwJYc/aWauQQfpkC5ApTPEfolRUc7dAnD1+MxF2dkI2SrUP
vxScwATX875v+q3ELbFE2J2KOrKzpdOXQvo88u89nC1OTjhN788pUo6CU9ZJmaNPXZVQBGu18RAz
DW5pkR/5cJj7KDD0PXxpo17kToRuRQWQuvI64bqmRm/2hMEE09cg5JOvbQ1+/2L7uxu0tm4aVqr3
hVIFWelGyY9pHqNPA6iPK59CHZHZEhgibmhFyMMGmC0OoHdWLElKY/ft/2XdYx0/qyDmqS30hgXr
41hhJDK+iqpgYJSJUDlsXgc1QBo01R8hWHhu85YbVa0HoyHQOWCUf3GztreMjIlCQdf7PqXSSPqP
ykN9NPKKxgcL6YDJA5oeHACuU8EPqKjd9JyiBIS3QOV4wOjI8O9DFsUn9almB2/0LyfNV8lpxy4e
rhmDCbqt+NjAMvXE6u1j/hY56lj1qA5I+2M4q6kmZVMNsU9RmhdpVcKy8J+xJ4KUMn7SGOVRtN4D
VhtFKXi672WMCQYPVKOEoPirojWcucNVeScmzFAbD3Z1vGStTX78gnnNpGDqapu2YN4VRBTz8Dgf
flI/NPZIVjLW6U6Duy9dSH43lL+ZRfQz4eqNj10T6vlJnd6jv/OQ75l8CXjSvqRrQ+j69/n0PpQe
HuOvoCZ+rztqPUdogl5ffF8eIAQiPkE+KCygwVoTnBEYFImTAGZjLfAhkWh8OxgyzgOWTyxrc2uF
5XQQsie3XFUYfZUmhUzWBqxPvnZufvXYmKcgzTIxRsOHnA5zS5Ddz67IH7XK5RXz3YyLJSJf7yPl
sF2XUANjaQhS7zUhM9A9eL9nMLRh4yBiIAn+PffvAVz8qGJx/DtEgpCDZBs944WyykYy5RIVCu+I
KzdNdAeebNCZYKrGpVUrxO44r4iKJnyI7fJIDex1/ANgCK8UOGbeWpYZcKHUUlaBsyzEOIm9/e9b
M4mABUIw3MDHlGXZZoyr3CLodGO1B/k5+wes2FCfXieAeUDU8BXby2LGYqq+nqxUm6b6NPcqAqFs
m/Ti1pyJ1pdgypnaWJmcY07EeAfY2uPVVBdoOCBQFSzJiFGuDSq4tfxZ301Cs5GjoshCyDnN4cK6
vCCoznlJSos7BjkUrMQtnYY7dTIZiW9A1rIbZJgvktJZtRUbIpBhP5Kx/Y7OP7PUAgx1YCof2uHm
DzqSg/q5mj2EMTGDFyOrxHFuhQxI0f0RXFAhq6JozF9POStb4Rr1K5flcU26bdNt/FxAuWRuy+kR
G76Z7b2Lj+/0iRrHeWJk5nE9miP4ManIeriSn2BdCsJjFr+XCsi2z+P6OvsGpxHZgLFMxq5NNyPs
E3kOG4+3dVYxAPZG4p/pl5s8BAMuXblAIqz6Yi/aH3Y/D/8o6C3fFAiRKMzBzrvx0Lcj+M0OYaNK
wklyC9QQBHuWsOeTMKfSGQYY1h7QDmFdHCvKKDV+pnuRHVQKHRs0v2NOJfxrg1t/FOfk58vgXou/
K9IdOvhslK532+/IvVuQMFwtWp0o738P1BbCxwP2iygclCc4aC4emOs9OhLqc9KbIf2Q6pB3x5OU
Zh5cbgBcY9GfAsLmud19if/4JT/Yx/O+88lACrKPUpwZu34NN6qTna7HzprRrjx793qAXkcpSkIh
/AU6u2/ttg9FHkDm/XmskmoUkqtYWJBvkSac3eoroaAoTbkJFOQX1EXA5Ke2z7CluGXhROVDOfud
wi4s1qdGllxaw8ppbfuUQbfLtCYpQgZVYZKKv6Nwf5LUfI6tb3wHNDC0MZ90wwR+xhQ4ZokjN27s
qUZx968uK8QCqUFKgRhda+9BRE1Y6VVdknVgv27FzKyDp6Rmo6MKmlvx5ocYPqse5C3YtAVD5e0g
y6qs1gVXzcjiCcmBdQLJzs2z8w0c7zGH9oOTbyYNi2U45buzxUps51hCJMOUFKv3lUEstVK6r4BE
W/lY63KROAgpvZJ+slewxHd+dNANd52CMfJQ0eNyknpqHD648N6I2ASlVM0bPpm91Rv/62p2+k4x
I3ba3yLthq9dRiete1CQ1+fC7/NnAQ+Y2TPG4kHplOXxGMcMDAiBo4ZH0G0Xgj9DQaLHQCgx9Enx
wOY0se0gxqIWIBY5e+3/67V0eKFGNgY5dmvhZfFOKnh07yCBa29tkyQz1Kb4pcok87h642/JI7JH
aKAV5EI8FaJw9r2NZ7AtBOYC8chTNkHz9U+/UI4MXXMaKFOcVbFfgMb+ACjOzHUPVj46QTABtrtG
pHlZv+Zf1gEO3MXbvF+Q1CZHwXELKU8DRqUbSBI63mDFrzyDYYCBn6ICqNaMDY9lx494NboSMeRx
y2FvuHqPUe+Ic+65aFpxvuWeId3WyZGjcafm3z+z1EtvE3y1dagKHP/WIfbi0ruW4Hp550lSN6qH
Y3dZDNiTgOc1h0kY2/4l0JUriSBo0joKciF6xDnh7/BvEzJFwsxBujzqFclIAsYPU4DR1mLcET8S
DNNqCIfuMv7vjTuAau94u2vAoHVXtRagFbzXVJsA1V6fHDNuOmo0tNBWDo/kgNJNEOnn05ukCzS2
oce1w6y8aVXRbG9Nb/BF0DFfpib7J2ygPs+ab9BeJhmJn0lqZ/PvPJ13Dz1VYnhevzPsc33CvkJr
HKqaQnMgCMu71WHBX2tdkfWGTwS3NhcBOVXai37ec/8DJGQFhnaEPK0z9G2QnWyIXYGP9hi79Nbi
Q8BsAQV1hNFZUzToQ6iPkrLPx1qdwbFRa87YMnmCEtHRccsBl464nyPbcOo4n8y0QUc5G28lv+LI
MoZO8BKcBdPACOKK3mWzLv4gjeZYGCS2WkmZKfdM/s1QssG+i+DGM/fI9S65mAitEoAeKr/Mk8pI
aQMcp8kkEpdaA/8zNbEefyJQO8vbIzoZ625TcJq5KAE+gXO1rKndcNpLtzO4msNkIr2gsEdtJi/7
cAKq2EfQCykIiu3OcEfbE48QdT2OlakCoV3ZStyyxzppD282CTKAxZxqiAly+033US66VYMThDJg
gCsP6jHBOQeF2mKuCGZPs39f7ghOi/laO9lHGz2zmsxxlHHUNBS4oCaWM82V04d6zHY96rKbUD7A
WyiuFBE2GpnerDmkjsLhyqkOzPFGimT7CWGc73FkNBEW7b9AGVGJ9q4Lz7x3PpuYlcrQR+mFhFvl
Q4MgQ1HxlZisHWbTZhGUTGLxxW7KKM50oZd+LW57FBDMq+ynCPEVTD3eez0kkAH01gV45TYQj0Qp
I5dUFKv6Dx291vnEau76alRWwtvDaksVGLdLMe/nSK88KbCkMEM3PbjTCsV2j6d6bFwB4NiwB38N
zEud8GXzTi8STvMFNM6faIgLncNL1erC8uJaODqvsRtW++DuYptfarneuWAUDOX21kOjOBWDZmAh
pfVKH/e/WJSFfy8qyu8q/yZVqSRW+k41ESZ4SgVTq6J8+TxPmOpYGimUW1YZ/qHachw/N6lqjo0Y
iuPmycq8pR7Io0UcgChikujTz4mOMTNNr0pgElArH+BcST/FlrzIv35x9+cDsbjZHjNXveNl8F8v
tGCyvAm9xFk/rdk6i9SsyriOrl/jElnoRaRTuQ12SHLvwpkkZ/2fVvqEBua092KFek/Ymz3hEjFJ
bqwpUDZlIQhxulPWuMyeV3EzlqnlCOiYkB49OycVerPpcBDjHGpg5TVYrZx+iSfRSHuJOwf3wdn+
QAY0Lk0iIKIyQbikBkB88plXl5232SSzT9lF8yywEjltih34OcZ20g3jGNByNwMnVwwEwfbUvYwP
6NwJVvGh+H4yMzwQaTTtwNQP+gwKhUDNwv7diGlpqNMAPlyYBMXYIMOgyayzCuiski7ZQWYj/BN/
BuBqrDufpwF3ZeYtylFSMDwA7AtLkyXq9T2fo+dneul/YyExDI1k3nPzlID8T/cufn2wAbC2e7gq
nsLk3DHJdaRXGv8Hl6qIlTbaif/XsJ9eCxzMvVV7JVIcaDCo5/DsM3VqcgHUIoYrAt6y61GqEDD3
F8OvQ09gsSJ/iIdEBcGvufvUbADuIPORuQNVuVcB5SLl3MROejkVyibx0NQhO/sUuWKustsUg9Q6
jciX+4iKNER/wUjvO56fSVt5wjlpjkByIg2GJnAcaZ9B4bxv7BDijXASW1et2V8tQkVOj7xV1oFI
hW4SPMLV2lwxoEYV/cVoeItNJExWr320zio4XYnElrOL4I7NO12z/VWFye78E6AaDKmyXQ4qSe2H
ycUEvoPVp/q2y9gLLY0QuMSxaOtDilLe8mp/pp9hxa7JUlu0YKYsEpFSHQ5YJCVPdOkR9E7aw1Fv
AGx+m/zm3daryfgh2Z4BBLuqbQp5lsh6hbz5ZNE0+n/gOdpfSTObWH1oEaCQIUCwYWUO2E+8pfb+
zFSisPW0sIwCCthNEH+BLpJr849/bqemYCzvC3HPg9TNHqWYtZUsJSOXa1QRAacKMFKFFtLPp/JL
YLfcy7ujCbfspYhzCuTlMTlaubhJrSZNDMNo5htyfB3i0RC+gqqR27noHIfQd1OHxQ1W3IyOu0zx
7WbyIKBVwLMrnoMjq+DuLax5b4YbbbAy0vYx9URA6TuiggL+xWup+Gi10jM5W7x0dWJUTxt4tIvq
c07vLGI/xG32wcyByKm/+ojDVoARujma/YDhPM04uv2skMA/uWSjthaMSiFX677TTyZnpQgMmmHt
g/gbo5oUhLTwNXLMBkmifTBFPOuHfi32Y1zjQ3wJe3SUnSuoo6SrCzUDd49QAbLabx9x66Bu/FhJ
I9PmztsFrTe36Ng5CktkmYBQuUL+bRpGflYyjbQL/Mp2kWlBXprz7jwfYd0K+vX+IOa5FPIyWeQh
j36X8Rn3hDbFuh0HPRYwVyBNpjNCoyNNVyO9E7L8UG2OZP5IrJQ80DlVRtB+nFqPGVgSFgm/Pi1V
RN1sWI+yxj7f++mbHggwRLcKmFMEMTuxYzE3WHfW38bMvuAFjph7eD5k5TFXMaDmOHrSW1Kghcgk
1SfuMPFpJcU1mS6SD3cHjIj3g3jd4DO67WK+0/wadXiuCN1VTUCLm46SKvJSBMJyo9GZZ9b5kvn9
QXCRmV89VZIZWmNEYljpZEBBOCyyJ7gP6klqcn5stokpOw3n/teTp6oR8uD25mgvjKByEU3IbewI
0Txe+Bey7VpwaEiMJEgjFWlZgMbwMR22X+gk2mddl8Zy9ihjNjoIkhWxxA/HIHaT41XxkzcQVBu2
51fGs+KGDxMaNAFjxnglzI55TYlzMni1DF1rBpCZ/F/8DlTJ8LBA0n179e5S6FY6Kay9CF9lW5A+
a9d2EFMdOIzt+14tXiROmcn6AqAuoQq1o7zcLSqunwRgkVbopAwPIPKkgt7EkrLvl8OLTO+SUZgJ
0b8uuVfI4GWh3vTmTNs0w8lOPrCflwzHFDWAhfCfCgnws6hq0TLVVveOQqzfgIRX4ShvJGSLF8Aq
ZYTQf3NKzxCsRVxO0S6Qkoxb6nEWEIjBdlBEfVOmWH3LKuNIqLPaKUi1pbL2kxR0oi3Jid0g8Xdf
kzA+NIw/EY++85hQN92z0BMeL4sR5iiagtloNHoIrX61QxgTa+rklQKdSYL/V3ZgVNOMCRIfK/8h
k0SGsrU/HzJAWnhbPps7cJw0DzA3wOQTy1DiF03S/D5/4oSjbBSOQS0HYR+pbyRs4xe84op+TbrO
zCIM+4mEtW3/dSXPb8oNEkjXR7O3rlgT5otm5ObT3+mQBNaxZpH5vfMKD2hp/MFDuL1hF0+8hE2v
XSFG8GvjDa1/i3cWJDBQZEF2/ghmxxfswqgZuEJs3JpePJ85ikdY8Car3yOb6PJ9s182cCkO+h9f
B86U+xe/ekADTyeK8n1id3hcXnkuQ982wiYQ0JYDJRCAcZd4H0vtcY6lZRjCzQQGVnYKXSrZ8qJx
4fKVL6ujbgmrE7WxeN43hnVqr71tV1SR4Lqxt+C9+ODQkZeS2W0jZxFOIs9lNlPAmxjn97lw4TjC
U3YA3/2f1zIL3napweEJ2+8Wgbsm+aAK8JT2BVCgegWWJ7DaExwx/uksD6cz4tSpRW6V4Y+nt3cR
qGSJBCtsjc5l1b1Y3vopv7ywgY+9PrWTJ3DO4xsYL+NXNJGuRBrP48anAQWkIFCAh1BPF8qgvybf
4y5nVs1cbIwjUiLEbrcBv6x6QpLXCAfJtReyoiI31qWdzX28PtwS9UojnnTjvdfX2oOurXaKYWRf
MxdmpXCA8Km6+WAS7X6ghS968SdAXkMyHN37wzzOn9FVLTp6f9vEDtJ2XVoODKbWZiXyTHoLu1o8
C8NcNczbUfkBIDgq2CybuvDW1PbpSkPswHaLT2fXuuZEI8ADFxQTXRmATFVFd9kJPXs/tXANLlFw
/SidNS785iY121/NeIdfFTNe2qOJngygOnSdt1EZ+4UtudXJhuJSfoeOOxGjlRCItXXII5TkuA0J
++sYgg5Fed76U1tD2RrSt5SOp5Vlio4t/3E7s7x+E/CN0VtBvtJyttSGnzeB+GFK7KaZ2fBKajwk
qdC/bXImyoNkfZNOHEvV/7esiqPpXmN2Vi9IvfFIoctBBdzPGy5esjY1vXLMKVrdSRTCy3UCZfZF
Ill1BjUO6WQ/cp7a9LEMpNWBLc2yEz6FlD5ME+TZD98kwXhy0QdiHS1+haTxu3n8mIVNjK3lH96h
wx+Y9924ff/cwHZ22wZu340VDxEdumOO/Pc2UrjFFP7Cl5gvqTTDj52CnfJAbn3Al6Jmjn9pRLyB
yPTyxlGwcJWaY1/2UIvqUpjQchI3KzFFE3deDIVbTt3iA3E30EzuyMPOHdOogxjl8m+xPRIm0nl9
PCvDCwNQtkRiri+S8/UiElFWT8Vz2q4+Esd22jy1E7Y5Cs9eMV62I4af5T4EvcH7p4bPM19YLhVg
eAucwEaiQRRyPDeK+9BkogNoAd9k35/4XQkdcSUbfLsgTDgYohJDrRC4qjoAZPLomaOM+toLBCsp
Rp/7nE7fwL450fI187l45+mKCZNxElevxg5qvPdeh3LFltCVBdMsXNyfpb6iO0Xd1ZFD2N0CyzPR
dsAIpYkGJSxLKveU+a5odeZNbyQT4L2bJXwdgxSiPWgsDIqM1KWLbnPSUM7rVfOTM1Fjpn43yaD3
ezzod9OJW1QmwZBScSr6TKbm7FXh+ydscK2uhwoHjjw8bJKcy7AF5GUpT9QnscRJMwZnRXDUa6SY
XAWaqv7pCnyxAALFlBrafDUJ+o4ciZ17VW00wciP+aKjsSkqqpo1R5qAlWLNh2NdBGU+DUy+HNbQ
b7jsp3HP+ElVlkBztb2NTNIqsnwYQWZOev5Hv59vzdR6OHXOzrPZkOqLO/L1m8ajpFxf4fLARMw0
T6+c+vSOYYD3BLS0S16tMUae78RKykDr2JR+UYxgxqrwFgJ/JrBEPeA7UKyjjvg0VKYo2s6ZqEu3
5zLMGPQPmNW4nP2pf9Gtu3Zte5GPI8pWM+U/5KK/L7A4kiu7XGFinx/8UqKryKly6T7WUHX9dDWW
qCooomTn45y3GjwURXo7IFFQeEZTYDqh9QkOkDP8ZE3K6l5FFyWd0c7+WLE0n5NbBixYVRRPzX8b
DSCzeOzpVNQUDhv5fTIn1hxehh9b+JHEr6l8UruZAdctwLFz5t6Bx7WixUU0aRyMG0r4Ie0wJoG9
pQhEK7piWtqci5DaQ8QZovjxYbUcHFwOeTF/8R35umWU9uPhvUVkuox0leufmnaAA4Y6AGXsQ/iQ
NcUb+nnQtHSHbdlf8A755zIkI8BBSNx+FpZGmfVUg+bOHCeEs9mehCR70RsO4maIWAvRC1SDfsmL
SWw39c0dM4v/zLxM0c6kX3tE6JskF8JbSrkND5xjpi0Ef0tRqb/6UrdUVSZTKvNUAGwtrRAARpvB
w9CB7c2gLSBhkA0taDlfWNLfMQrJxeVZNFoY3OtnORhXD0CuW7tucAPz2fRxS63wpGuI/MpkYd8h
sCA6dszlsT8SVWbBRnTkLIfWiZG14jmCGtltvfdxdH5hJ9LzISkm9yF+T5UCbWzGNKgs5pIce0BL
PF/vADiLkn0OySXfqjGbHcXguhUipk7k267TFM3I2Cp/zz3RgZ1rJ7xHtrp1ypij6qKzOWfBE0Ir
XHLnjRJWv5rxsWIsUDzJlSl5UAhOQhhaPZ6DGbnJghzx13R/lO3H9Naj5wb/q3ZkCTI1MDvwEv5C
2PJNN/j6isC3BP7SOSnPA3QwjopCp8mHOr8PDhcY8BOgfnq2DMIn2e5BlY44XKcil8ZzG7qz8bao
qLtuY8rnbUINvstRVL9n7ZuzP9VnlgKTeJE6KMdX8RXU5B9MXx/lXopbYp/hDl9dl2DtYc6bIeVs
1QhukdLqcNPDqeBt9MWy7eU204KR3SFrAwQmnYKuD4oC7//d+LEJMgutJmxla2inFol/Gmw9TsT8
XwpNd7jWinv1o3wqxcdfqh8giRSBVlc2ZdLyC4zz/qK7S7vPoasffq1FuIsqtzMV82HBO/jh+AtY
NnjsPKqwOcObhZhxMYv/AgQ4AEgy2Cb+OOavqlCcS5oLIpylKzD1pShIcn4xhL5hDBibjUK75RkW
CGAV7M214UCdWDi91iN4t5lmbjwUzUaTWOgLw04LlALZek0BnZhj7c9mBt3mWXlkH+udrRfhYNIq
UxUHCuE7iFeOWXr9raxkGogQOIvbnYNUDDPjfh8JPX+XvPrfsLgMexM8XXn+F0nes1xt2W1oOm43
CBrsRghuD2oteVhSgGFfNjfavAuaIwLp+2E08tj1cgzmAbREEjdSYzCVtgQqymtg29i+izIuhCQU
lXl8Qz0gEhl148FA4K1Ofi/SNMy4uwEVO9p4Mt5mqEwv4bS4oB7bVpVJUZWS8aHo8dpjDft8xn0e
s0ON+O1JNeuEiYLQ0NCjvdVgb6MeYGcX0cTsdCfrwBeuTXQjD65r9n1qgKjO2gJTdXjiwLqeZ3SH
XTN4S4ZvjmE1z7+tnjgrP+yo8UZKMEaeQqiPqtVx0qUdODNBLRq2qSOwYxZ6UbufeDCLRkqqlmNz
E15Vm0eYnXLZN2hHcnJNHUfj+hcre+f0ZmOmRN5uzXWH4vgFe0q/yPupBPs8zS/wjStVK1WCSwF9
T4FOacf+fd+XlVUfMnXbfeO3oTeSlsHrCroT7rLNx5z3jT0PjNf4x4YdPDAnb5G0WiZQdbo6DemJ
nXF+FTIk6XEyokpWRRKaSjEXIkgs+3uA52mN21vo+nRkeTBsd+2cgDx2IewIbtMelA9WVP8sBjY4
b9F6Lwpdt9ARpzkvCcgsUwRsqYwBuHDJsKpiVX2UtNT9gS1j+10nmTxXmM0+/usxGDZVZKF2DzrP
FWv1abol/VcAKaqUQn6UGwfFweeyV6EYRVtrYcsn1xHAQJL8nZynnN4TJS9qyLongE446z+ko1Lt
SE8p9DyBa5t80qioc/i1gBI/JBCzrxtI3/KUEOBd+kavwyhjgv0X4aQJ86fs5cqu+dlaPO3jstso
rRQDS3fuyHMB5RTpaacQCiqqWpTIG/jw6mlNrulDJL1Eu1V0vJ3PLvk6ROTY1RRxR2DmdyA8dcY4
L2ylEw5tU+BxEGpuIzjiUibMLPigo/jb1iUVZ2Lz7rN+/cvL/eOdxA7nn28AbRCTEvlevJRU6DKh
+mN0KNtYVFwT8j74EVWxkbH6UHd4TlAlZ0320HofeZYS1yVf+l0Zx/3sLEjRncHtpczzAdO+xlPQ
5GWYsYrKKmVdG+mkdRxkTIzL1o00hgKSxgw+ATFPILctBFx6DJij8kcGCvudji41hs4r9zkoj2aT
0NPyS5Qhppv3/1edMYDvZ2TViHar+q57t5ecBfpYK229GToqiPq0SdNH45Rbg13x0vV3S5gDrb07
tn4bNp+bnu41tV0GWuUbZK61l5bMVVrzQ0SvOvedPnB1oYGcGTtgRxEsmEO//eDVFfKXdUPBjQH6
cv91NJDOksl5oSrz6Bz2U1FUmOdFmOGdTw9uEpMYmbjsF84JAMl4ZfnMJjTJLFCdrPwFInoVPUnO
IdHMNJA7BMeB/x6pxzYWBpaOSyRYVZVKvERGl8VyGb8PQJTyd2JKkPrirlfVRdLbvoMBcWRGXKkI
uPuyjEXCo70NtBwbW7mIBItG79CGqXzFS6qvbsX3J7/RyqvPzzfif+3Ds5hChXHLWW4Vbx+q18O6
RQ0ivIMUqS+txRHK1JH3eB0A2ADRHJk9NkyEtd315rbuog4nT2KnqXY2AVHIOfI6oVgiESLZGLSR
b2WaZr8ZWLxQRLbV739QYDu+K4V9myn+W1hIXp17NrIxOccaQkZgRRwFwhg2+yJK9XWAn8R1wSXi
/giU/6k2jD7N/+irTmr4VxOdvXlJUB+xtxAsRl9KgmwjsZ+ZxbpZWH6k3C2Id8HmnTYjCf9UXUrz
ixbpPc80t1fI6Eczo4xeRzoTUyg0++ydHyHHo0vUHo4jc8N/7XTWySTNP1y0Gh+jCISErolW2B9J
yT0gVRc3pobrm1L6JHM9O+HVZIQ7D8y5ot1Rxop/TiOnsiyCbX35z2iHKzk7C3Vssec2nN0GqUJe
CU4Ov1JhMGf3lzgxzGo2slhIOxNLZembgus8PjJnGFUZnoWD0bT8LsDz6Uw8NrdCr/7vr/d+6E6T
QpXSSO6zeMtCwJ/3GVZJ9AKTMEme7QCd195FjfrCF0V5nHuRt3CEUTlFObF5mnUY87zKrq0xehSl
lu7x7cgma4HIc6f9ho/IEBw9WlCkgYaoKhMA5s8ZtLiNlfBbwiXMAWaUQ4OIknqL3pLoDGmk/djg
WDC4IkAdz6TaNOD6aEjWL4seREE2I3IjCS+lrRUc0oejr/KdR64xyT8hOTQRxvN8iKz0T36RmSMh
owlIIfZ1qh86QG6LTKuMI8eu4FtY1qficXcgEoIzcmKhcPCYIeFup9SKKBZQimMObFmTHacKg3AZ
UYzu1YFJ86m61Wm7UpgZ2gwkit3F8k5lA1GcHK58H882Rf5MydAD/cvrj6BZQxx4gAc8SdAWnTar
9lybUk9IS3wxC5DGYa09W+l40Xu28eRoYL5aGEZlf8+T4bsRn+3FehA3SVtil6Ly5JhbvQb3KRMZ
rmjLSZLUR3rj9xsa6sfZF7E+kvVKpGcwGD6T0IYhR6lpb9J++sn3XVy+EAq/4tpCWKXbrRQAH2uF
Ix2jiKzPK/SCaA+R01wmBW8UqP9JVS48SYpdjoXQkXxOGvaMc1OqtTGCcdcxqPCZJNVHVzVAddk5
mDCB4J9a01pwq7gNURsKuJYPaqqE3PWySvw+ZX/3ykJp1x5dbVQOAZ97FJjhdhF3KCdYvqDL6Eh6
2GpUhIGr3z+F3KUF3J9uVrPJfXBd3m49+fK+DuQT0ydo5mtOqNx4eh9cTzLdyUtcO8nTx+iQV/Kr
myfiU8CEr5YX3vyC3qxlg2BL+5DfjIn8RxzlEvDy55bDvs7DKCcgdGrmYA9lXQLxFshigD7y9Hu7
4HRX6b1o/Ozy5dcQtlvEhZ45MXB0dZ3ZdJlPryHy7tuoFq5ZxVMa9+0mZ9QIEv5rkNi1gAncpumr
1a+VyTE6RWY9jrdOxGcjirq7scRVUqJ836WeORZ8x4h9YSL7owh4Z3drr0yPy2asukz8n7gstBg+
0LLCadKn2EKSrcHP0scgQBMwIdY+rwDINjJLSdIk9CbZ72eHua4bn5O0Lr/hz6HUOeLR5HtBkHQY
b8y/C0DMWKvl37UuV0dJC/XClvQInKr4n7hS6YbPNYojZJ3k57rHxiT2o9Fjp7WIHcgCrEmtI8a0
DdwyG6/sbC9BZSnG0xRs8oJLHfjCiQV6G10rJgcEJpAj0dYiRww9reWfwMpW/ao3yV8i++UbyW01
9Q+ry+8yMgUPWHmnTOTWGkI6QIB87sYbgELuyxYvZPt8lk2NriXYrYQCm/aFn0utysfioIRq66N0
u3EhhYT9nDVDIbokqpNAr6y6mpVCk/PoVlxY7oYSscSfIxwiTaZ8BSSsEjgGBljvnIHKcfWOE7Zi
cayAAJC0I5OTsjIU1B9fzZ5TEZCHzYz4ewGT/BGJWcTwR3sXrzLhTyh+e+TSxhl7IuIu8+daCbr7
yKUPP7Fh7aW1szVFjJm5jBYEHFiL+LEvQgwzewAfVkpmZHa1XTR7f+bdgWWouQFz78rBkjjiAomx
TW7B/m+Tisa7f10DOaE3sTRxkbNArczR1E1lpKdghVfq1drEqWa8P8xzTJgjEnYzgLRNeqlupIGF
jH+UK4eOzYhxa1vOSn3n6gP2/6+GyoWiG8OqhdfwVpjaVNL+tbbLbkdku97ITPwr1ITvkR3LtHcS
5X37VMWwAFMnQ/6YktmYvcjaO+m8D0MpWCQqIoGKz1EZRA/tQ8Q54txXh7OXyGsBA3H1V/sYcx3w
embX4ZgmRZIo6HhGA5Iufg7vKTsJ1FqVD/TYSk8ACNDJqqQlvHkratghf2aToyCCCB4jCVf/q6M7
T1CJsmlUagoB6VtnfeegcpXfV0MEjISYjSNTQrDe6kf3YLQiuIBBPBq+uoZYJfYRG5jUvsOkiSUp
ZkKGYHRWVu6epQQ8pMv8mfHT3qiCM/Lt8R0REmmPP6SRADciKDiXyDyRl7o1HaJixfoN8kiRVO17
hL2b7RY6uLo/1dOWRF9vRu2QELoVmSGc0bBg4bs+FoUpuNuRKLIJZA8FprdsE4iWyYc7HsTFa69S
p3BfKVHYk9aGbALoYj1EgH2aNY6f/oCOewjS5qMPM6YaHI1O/8+5G2OFmqmfj8PDsn0kGuyzR57o
wx3zBckmmHJP/omIe0MpGiA4RgyhEEcW2/S9ndBEOba1k07xQ0sAOqUOAaOA+fRemdb19IGOcX0t
l80F62VssO+HpTTJbuGsMvgTWph/ZTercuV45ufSeE18Gw1lUhEQ6M3lMi0HjFz34EN4tFZ/y1yZ
GA1jCHm2352nJc22z4SOTGkWEuI1q8oT42NKUqjxxzdq6/6P28mhuspZ/6Z4bOVCTAV/RjzjH9Il
62G6bEYIf9NDrh7Ze/iIpuylqFaEukYv/wGVAW5S/tx+diiBhS5tmHV9z9OIu4FNcrjlQ58IusNd
/dQsrdeMew0UnJgvZ6+wDoO28thMG9rYLJLkveDiE731BJ0Rp56YfnpxCACZQYy3f6o/Of+VPMV6
Y77KCUY3MVbD948h2AXU9D08U0eCCrr3Miif/tae9DbDWliuIu5xOIoMU8S4OhTw+dLVQ5WRIW7i
z1jf2zJIWMp01Ksfw9aQDE/AoLlK0JMCjQ3I/1AOThjHBQ/eQAhpAYGL0OG/5+aA/sRaU2FKvPiz
+FiQunerLBarkUUN2V1Xwrh0hdccOf54F8iEq6hPMydow4eai5UmAkr4uJPqsMCqakvEMYY/MeKK
VNo9Y86p464XM2aG/A9PpoMKdxIx6TvOLPaIcZbUVvTLY6/Z86AaM8gL+JfgAWYU/zGGsjb6MV9W
ZFTE1bGZnpC9wp8iJnw3QKly8Kpzbq/3FzHGOWHXWr9EvwCojGrW97P1e5mgHF4YEk3+ThvRla1I
0OXmwDGGYIU2LieCNQUcgpYzufP7aohdhyvLHODcLrMtgeeeGLe0D6uqvOPcFM5zSEZOpLmC0+G8
Yi/2/UZWJHn5wwoKxderK3qtn4imRGdSHenG6FyBHm9/C/utaoFDHPbJFvquoDnW3r809XVOoHrP
JavF3KLylcVyjiGLfM4a+g+6LUz197qBINuGOJ9y8SiX/T1UThfkfk2/ReLMFolXS97AMrzSPhG5
Y9rxRscciMHnl00FPzpULamBYay8pK84VHU50oL/CDLVPfT7MTa58Om6olOBdQ/HKA9wW8AwphGi
h8/491Rb80HKiZMYh0cHiVxuAqNegpXFI/z+3pK+33n+kOStzhGt/OzPmrD5RdqH54i6qvp27wLx
f064aDUOUXF1a4BvXZReAfa9ZNgaudO+EJKNu+JoI8eGHbNJ2K79b/1tzKJxWB5Hlop45n5ijlFz
ofET6k4lLqntou1R7hPukS+9Wl8oNawoOUMSEpJoNlQfLGyKmARcxcYCUKNjxhpuATj6xNzjtV56
aSpbk57AlCaTYFuMF29GQGGsUGZ+TPVOq8gKlSZCr/R6yr9qPgR66ZzKqA4sVwwf5Jka5DOKxaIH
daVP4XEoAJCs+SoKC1izWoYZLht1tnZZIGB65RkHYDXNOYxsQXmlWuJEerRCsKh/pDgj0SWa1tNR
3Yt+J0u8WdD6MIBfwTXWKc+3yLPoDEHF8sIMkYf2Rp7d3A6JA1EJb9vHRUPL5WRfFaIXikdTDjry
4Yjb5Nz6zuN8zSqDFZPy3m6QYnM2k0/Ke2VMR5JZwEbx+PRwgocf3Q+LRmvsGgxtAXahWUzeu36U
/iQBVCiZ7Gra9qmLExYmckVrNKlJnv6WNTaqrHOw17lUkPHLVFeNpDUQHGQd5RLegZ+yG5eTTcFw
T8aeCKorlfiIzktnZWtGtljNCwTwByYuA2WWBNShM9bWYU1jgF19d9SyOR8tH+3UXrFzr+cL3p+y
2gD5FhIwjBYuxOGa1JjUUwLeKPH/217dQ+vF8ubY/2zTEMLl7NrafhQOd1UN4nlTVnteK/cfVwD8
4ss75DY9PRgg9cw/uOI7plh8fnfmqfu8Pu4JLthE5Y9g59CJcsPZ1fCIqi4XNIJ06Z1M9hduCScw
3BjESj7oQnYwF93SjUHB916pGmtFYlQE6uWAXI2Y/FfsdtA0fdG1U/sX5UOt+oYF2wCcDtQvhmNX
4NFa5mb2iVCl2VbuSHYvkuXSS3Tc2Y5lbvSLXQ7m22pOf9GtqPMVC+LHcLctSkyXl91wYpqyG/WS
L8pomBKJm0UYfYG5EtjSWGIQw7aK6ogPH22G2VsvK1trzterrAZWhSTJeObHYegAGA2AXVz8k/bP
SUgY5Ea8RJOERj5hlrX0rSF1PUHyKvcgzEDiFrolaFNn4Ps40/uhMVHGIj4f6AO7yD/TltynYAz3
gdzp3GwPoQtGiy5g4cvfQQYcskOdQH7NTjWz+kwnQ7n8Pm1JlmM1L2Z0qgrKTgPNrO7apPXuS1hv
FKXzu+VMbgAld0dRvCAIA0+cN4XSw56vy5xsYL+RatKjtL4U13IGKZtzAQnYDFrb7ykBEmDXSkfj
I04FBNoBZL6UnqA7WrhUZJeXwQfdYYIwBd0FIIOBcj30aftoBiQ33WKoVpFUQuRYRzfXQyLip59z
Na8txayyJhX4GCxhr5TJC03hYY1JJLf9FaBsRc5gl4Gjg+RNQ6kWGuEfg+7dZgsV+3xOythXWCBM
4zaTXwm5o3yoRmLU7wtqX/YEFkpHSiN5cmLTZeKsslH1pOD22PK/yVMWDkmU9yGqV5JKsei7KwGO
7/7METf08mdZf0dBgETXc9ceqTiGAYhbNy0NylSUiSEXAqWzQR5CTYhncJ+hI2SBwscNfYtRGKS2
uN2SRILPsgYkYvN4Ha4Bsr2uD4RtGhffvdUQmX28nYqEl3B9bTEAAIya549zlbNHuARv5iORvB/B
AJjptKyaa1Eu4rso16DLvcJPQEK7nuYKeHD/qaCW/hpKqHM/M2a4vlQnWqfYATAy20rvHY5geB2z
EJM+TmcMQFy28xBbyCGKSQs03KKa3fWnF/rbS56W1cUndqkQLcrV2HsiWbzUTEB2GZpKtPDIoqTS
qXw4tG7V2B6fJNzX0j3eJfd5tPz0l8ku67lbS2m5/8mRQNOoQSNF6nDvp683eTsRbbZsBMLnkBw8
nfyiUIWPWmTIRY7u8x/mpnpHDgPWZQr3L1ck0SjOWwHcmKBu2fDOIV2Vs3HzKxqt2ToYAaCyTRbE
82BmV0j+sOdtWE6og6Lrb/tr1ZU0un/ToYZWGQrF+ShUyRb3w3gTNGPLKj3tR+zVfjDlEzxx2zXG
nIlTexPx1t7n4jUnUXEDDknYAjdN4uOJ+m1VX18Ci7buEtlRlrLaShABEN1LB/kGwAroKnYClKvn
+5Z32PFFHl2RVNn9AAxpKDE2EQorqe0GZkJ9t2HuTbHDAh1t898o0Fb4h8BbcFnFnnIFcaaYKG6l
1GZKHzlpwIK1Awes7a17JRxk3/KoK2sqF8qtn1lQqHM3PjUenMYsxEU2g32+/o5arfgE17o8LGVX
CXv/oFx3DquPsQBHz179VH5LydeheuRTBs+fZtpNW+aNzWNSgfx9gj8a+2TXsEOki0yMd/roYUrZ
WRM0fsGGcs/39I90+K/+BvIuWzQ1RCcWAZQGuo6coBFqLZhMD/Hx4SHf41Y//zDYQ9D7F7znugQJ
Qn1LNyJwklKjxAkjLju27/pgndh0mHF+BjJBoaxqIj5J/iKo3nMjLZHN0F1okuYEsI4LZlJ32+5K
ohz3VA0zP2kLz4Z3mr42s4n8xSOvLs/cMvDJTOHq6u0IxtaC+yLJvKXTDIAO0uNoGCY0XRrVMxOY
u4tWIx/AaPJUCJ0TopfVAMIIfxmayKNr+QpCGlnPuPpnygfgnhN863o0J8kf/QZcKkN2fuLBCTLM
peLbGxgm9hbdXjqa5MVrQkhH7HaPJUVAJEUrAsrRYd/a1rkgJljGjXboQbpZJiBGGLau8zt4QSEf
j7rdCiM0OM1spAeT2n/ogGCpxK9929T5QzkaTXAW1+7BS3TY48Jd035DRMrMzT1Dkkxbwg9ONriv
tPVjDgs19C9cL6ttpfJeFCMTnvXWhRG1czj2mAXJ+tMydYcN21aPeMps8Hqqk1LX4Ahx4kAd8hJx
gIy3ftqbZdy25RZfo9d8hHkBE9YMVQZQB8ZSTl1xaPixFXOma0GUffcPvjdnUgofaX2XfrkCu4n2
A62IOWzjgxWxqDA9RJTpVC5j35XIgrqWyaZLS7QfkxMfSumWQiLEjj0iALR7peDJcdTBPO88LXxg
5Lj8QEVISL1ygZyYV4Winz9ebJs2sE/NbpWYS5EhXFBtL1ZcVrhZE6CUze6CD1MFuya8StfLAHWQ
9JztvSVtISBkHeq5OpdQP+wDicnXGM0v60CY4g9gvQMNnkR3gRGj3XTN3aU0CM+lxG4MHG04YW+i
ciIIMOhRuT+tSrvNci/Hiswl6T9hP1ULAh4lPp5jip1C+aToXEyJf+hgmfyepqwxgDLeDNq/P2qa
5nSNnTyUPyRV4/lfeBOxavIAmeMbFmS0YMOOQwkddFteZnAsn2vxOeN+tOcV6E2cF1yEXzxpaf/m
eDszaYaVDsgt1AaWx4dr5TeIUpEi/aZdvmZVgaXxTDs4jAtQPrpSEndEYhNd+7pUmpy9fVC+WWzS
TUbwl4nwuHP0/gHRUAo5/OhLs+HCkaMJbxh2DmArUUFsk5n/2FHInX9xLhnPH5PWs1NnXWXm/dhW
erv8LR+HTni2TddSjgLwCOzWy4dvHUOU71WdHZalDESrpXJxKMzQuwVwu/3gTMV7+2ACJw4cAjIn
/VULKPX6oj7w6pnI07NSie+o2WKMeDyi95J2mQG5Z304FAzNOlNEEH1ZBYdONz6M6H3ald8DNVXl
Ig51q4iguoY4PEHvwvTUrCBYvflHVQE+0tpYWZSDxT8RYPRKa28A/rW86+W2EyTJZIvG1DvPfRBo
k9IRN7Z3sMgiagojqIxo3tNuEO00HbJTt/2D69OHIIOjK6hvhObRG7fXmh/gx3s8Rgg8+LeYxtby
s2hr+ILEsd+d2oOLViuvV6H4mMQTFymEEvpepNXbyQG47KZAfODF+nQZoPtovvLIV1t6q6mgc7XH
gLx4z90wFuqWlEBkP3Z0zTuoAXLEqKh24CzPu+NU7NtHf+LzQ25YsRvv8dM0f7l7cO+Z/oaimams
MJJZJ7pW5CJFfzO0hHL2vytEqSutBRdybDWfZh5z3c8N15NcQL+rk743JVxVUWcsUtWDOsQKs13K
wCjlgvG4SyjeJrWmVk3HlB1aD0cWEJ/00OkbpjK6KD/utUlc4f/HEPIcTyJU1RK7/zwr611WS/IP
doB50HpOVxz4UITKYNEwzfHoPnRwm7Gh3jGjmJTaactzENZZband0dVj4QG8ovGpUbUUD8eP8ZBk
g6yKJOSMQmaSYszc46pk2aprTsF2AzFDbnwQqlS6JG+LX2NFmqf2YigujTX78f9pY+0RyaZE/KTH
q7WJawMccPWBTo2VHGrHj6J5B8PzmDMfgzKBoRmyvCYWqIQ3Yt8gWel6BxfZbDoYerbedoXT2f7K
Uo9Fc53/5AUAvZZGhP9s6IexYsl38k65As0HTWZfw0b/EGushCp+geNMtnW0nCjpDRHwBDqPln3T
efYy2H2RV4hZUKS7HQ04ql+LQgJEUvLFyVpLD8oPLZtOejowmtIsGvnT+LdTJ2+vXQvozdWxvGz1
YZe5OL7ZnWdMnc0KnTFnwL+mJUsuRrcd7YlhR3OfSQf4lt9MPZuRlV+l8/i8AGl7Xv5YephWaspK
Ih0o136DCGd4ABAR77kx9vsRBLN8lAeX/zQ/9lfaugPLLgGszrKvsOIzfPGRut6LEpBvr970ytWs
vRSvkmV8URl33svO4I1x8PWAYSiamMJQCJww4YbE/CzWiXLqxPVmQR4V+J01OBbr0dPcX78epKZk
NHWtJLjnl3C+cx4dWsgqikUmI8/sXQG1ztnO+PWC5H0e4qN67BOACIf6Yd/gCzl+spTQhVLYs/qU
0XEzqETdTrJvrCCl5v2qYLxVLalAI9KoUukEgsMl/oNTRsmQYb95mMM+xr3gFixvKcbmvr63nH1Y
TRJujx519N+hpFZr4nw6FuVObd35NgLEWaACmjxjtGFaykUzlITwIm+yZVuzb2gmoWl0e+uCoNXU
CjyjI8fh/JuAIbT059VkX1rCXeqUXlX/O28r/vwUki4DotAOY1gwVbKE6tFFe82LocrvwDMTZlUS
cD+6fcTby9EokauJsmgUpbMeR8o5onD02mImsFjRG4Bd2IOzHZ9B8qpPiRfwzmuoeJS0XlpFymOG
Irv6d49JfUB+q4iHCDTpc8IavCNFBby6rZr4Vnbh8rEayJH+D/QmBeA7hQ3UblRqvuPjBAkpem4c
ECL3LvYlxXWPPKMWhVXDPIVv0sNmtLTfom27qDcTRd2A23e7RmYIEt0zeALnMiX/7A/oPFVk3fLJ
a7B2gc382IndoibB+57azr0I5OiEF+d1MG0Ao+2oUTDKXEy9JWlxDawfVXUdDRrvKYcNPxV/Ysw1
6BZQrq1n2FmLx+Tze36FrRq+hr7cMnxa2KNUIPl/Z+VBb/7HNUThwql2y/BwQRjgatBTAp2NasM0
A+RsNgv2cGVvGcPKDcgkuI0WFdaNTIMu0/1MU19RBIfMw+fnyU51RploEteLfN8uCDGI0rLicoIh
sTpnN8/udc4zlkC8LUDOMFFA+jEVvhbK8mgAhGbnhif1D7gJcQ/gUDjJEHqtdogizHn9Q5h6wfHC
GE52kLKVi1R03Ess6Q/97KPsxUQ11f1DyJf6kLEEP/xcf6tdstzCBlKISW7vNMpp1h2j9hPDkNJ3
SZDHo4nRAobhXkiSCrL5R+/NyyX+ulh4Oyc8FNAbh8PP7u0F/1tEnHvn1N6em0mBduvARPvZ0vvd
uquIFnztgYaqkEk7JXEC3RXE2k4+IWu2+A4wsq6LN+VU4qoDJunI0PnU1HdShI/18glKQOfR4mNd
jI9goZZ49dIw9UhrQgCDzxdyd6sk6CLTktuTyLkpVw9nxUYF8O5uA7oaro734ErWvdjf8eehWVZo
ALvCjRKK2UeDmukDhznkw7MVuaMcQ3GfOBxnawq/BR3AfxSHazOoKNVsIsfGEoC2s1RJYBn94+Lw
sE+8NP6juvcvBnbqTrGslpkFQ7NvcIkVVCRa/HHhEbd5MWvV16UlKas1ldpORiiKOtTRCD+w+LP/
FP7CFCd/s/fRMjr3vVmQUX2FSxn02S39dr5VLX/i+i82rAXqJZsntuvFua8PYs8IhBQ2oe0wNMJ0
ye55Qbrv7X3TiXKtqFrfoSE0SA8bjNIIJZJq9PRqZgHUJOoDLOyCLWKOdkDSLsGjOa7fRfe7sjd3
nvwLGlWzEX5rhXvjhAygeLIBs4Ov+zfwn9GP8U3YiU6d29mZ/qjSt6FDQUnOPDoKDn+QY3ws+gn/
3QYTV55mv6HxjcqvgnfSDYlrWe1uSYwXhho2VSpQE6zNHnCLRad26PeQ4hwDHdOEEJ95RBjeDhoH
HvASCOftPxH58L3zvj07RSq5XYDakYORsS399cScnzPE/RUNxx3X1ZXpp9FHK7i+EnCUCzpO4COY
Kgd9rjC+cF+0DQWt1uUIHa8M4R8XRhfoepkI8R7IPOO/KkAsyyiV9dvO9JMXyub4SiCQkJAKVx8I
wfkcAKGRXC5iGOEB/aVnEktvlZmUcH5EIgmqdDpZT6+ppGm52qGWs0PYDv8Hz3Mf1UHfC6uiXW+Y
SyjqDz2ZTaEY6r5KL3aPAlYEeZItQGtV5dhI5QnfGO95Ej0x9bG0aZTfODxOETWCAGz602o0wMkR
rR4IZklphgi+bCg/A50m6qnC8MrWlJClvSw/CZSLyrd8Kw1QnUjfAeXj2GTTR2Y5WR3jePKEe1nA
T+YtEMCNiws0p75bWzZAYdbwK5+cOXKfXSVkA+tx56/qIkUmkH9C9sFfq93sF7myqxDtSzUNz2Hw
LA75IlGmIA2GCgmgWZ4gq61o7njArs9fydDfvQ070EbgJwjpXb2VZR4J2rweTUMNTkBsGbTIApnJ
EaH8B8F+neEFw9qVGolzCOQ/P/S6XmFsAyj8uSB8wxF25Zdm+Ci+32RS3jskq6ypwBjP8frxQBbR
pGDGFVWyC6ElXadtZ+wNjVVzdMdMTuy3lBh6tIq1+CHCrPKNdjvBAfxW3muABj9evgvgvGkTXx3Z
jH4RADOI+NkUmt7CVAskTLULRPFiOo4OjKK/97dNR877i7bU57pvS0gqjOPEYgw1pBPkLJsuwmB7
QoWhfJzsAW5jX9rG5UY0jwUGq/Xe5XtOdNWjT1SR9IWHHn5JIfQZtMce+3zrNwYSMwR0UGLptJ6l
CNUu72syQ11F2QTh/eEppuu9wQGj5ZihUKav5riSJaxg3nG3HDFgCStEgvJiSbVGAulmq62YG6ME
RkMiIaqpW02uVKZY1yir2rBCiodfQr8p8yk5spgty9uxwc2DammTVOKHyp+Xn7QU1NpVckIDwujR
CgviVrrq4grAMwYZbYJ2gcqxEdOSyZyCeMeJi0kjVOQd7g17m5AX+HHjpS/UNYYcue4OjkpjES1Z
sZik3HdL6IL2WG8+vaH/liWL1ykzl8fX+omEYWh3jWYc1sX03Opr6T8IGWhY2oDq0qB0uzKUpDPY
3A0AC+85e0riAlR9mdLXp19Dc1bD97ToyymB10LrS61iMSbvOUXd/PhMvkLwAr2hxseI6A7EhypF
oY43G9ZrliWvbqAanI3WXR0/+iZ6JsNw2RyuugFtm8DMT5ih/dCH26wFlkLSmUCdSyUeQsuXTo3C
1rApD4NO3Sqfje7VDohNbqm+15Ber6/xaqDECCDN/OBCh3NaMu8Og5oMnCbN9Lt/HejDxoaNkfk2
ZQrGOca2E8nkFBLMejESbTFhTli/LbGt7fOMhrtLRZY+K/Tws10Qy/g0IuC87Blw9DjRrn+cnSsa
w6gU3CHtL1mJ8aDTNM1Buil34ghiQhlkv0FtKoWB7RdfdpNKKnbFtsFLN4rTh4Pt2opd0r6iVNbi
5GRDYEg0TxABF72g2s2v/FsVJthlk1zSJrKwHCc6qHs0Xg/Hm6L9U+yDAtvipozEwt57Zfb6F3MN
uA/CMh4kkcwhc41x1x1YkLZne9HHu2U7w+OQpzqvMKjIfvHt3xK+b3C/VwosmCGI8ViVW+low5th
SF8zgxYyWARyfO2cI6moQTecR+7FT6u22801u9H3Z60rREqAHcVmrtwyDIiILIKSrC/Z5dDB+WW0
uzNdSFDG6WdFMq1X6d3Otd5q6pr8dUtBD3DIbMJOxBWL7Xqr61ZX9OsOGBvZJVo63AVMemIDujA+
JMDKFvzCBtLchsxgBSAt/FbT8yG+ws+uLH0yyKAKvAIDGczJ3O/N6PvHK7ig+aXvEa1GeYa6yO2H
SrElU30uOs88K5L0ofajHprnKsMHH6WWp2V/S7FKpNnwZTeRmoSUGCvinCZ961owzkpng+HyxFpN
FQcGyPCC5dhsVsSYm/Gb0XWjKFVA3GLWiYSU8zAzpyYEHlBm5nWHblYLb1Z7dJZwSmf6PSNtKNd+
f+4b0g6QcgGkILRhmJ5uDsNhrUcd6llid2MGlJTFnNEOMZVTuQOmKjhWiGEZsiP8SSyPDsGVYi2o
i+VEOTmnpdOLgNtMnRjw0auuazT6E6sAC+zFnGSsgutM5zh/51SFfwL0GrjQziyZwqoZ+/bQC/5Q
Xwq1K9njj20moZnx1H4QJKrRnN144zv7YDEDPoANxISCKlh8chpQISJx/4OtDglt4okvm9fhvMhz
JWvgb9no0eDh7xUaWbVrvHH/zWhNszgSJkjIZzcEYe1E+DVfrO7acloNZFVuwbSqtzRGuFgxaKAs
tiPfyrZFjgyb2V51V2vATtr+Un15bB7RYBBE5es+xMS1BV9H8BgdE0JSsubyBd+CWtRVrTQ/HJF3
P114HuneKcw1vX5olrl6lOrWcvgOL2rJqXOPHU7m724TJVEL2/i3sYcSH/8Ays8Chr+UASrnB7DI
HD5oeGtEYo8i2uzTgfrHT11HHXGSZU+LMwe645v22w6l9AyfNZpWUAi9iX38+9uBIIAoRKQ4mtAr
zfrptXTFeXfH11ffu9+83/N/dI+yBUc823cNnYTL9rNq0uJwW+DDdqoa8USqHROw8ufMtpKZXeyk
0cqFjuNuFyAM0LNtHTGPwOqJ4sW3GCp754A0R9XNxtyIpkPkV0tVrA3VcJ/0ctZf00uX39XMQAj5
qV52pkaoV2OKVlOgGFZ4O3y9FdOErMzaspnx85u9JEN1Sxb+EfstCELyH9W3UZKWLsPWDu4To969
LvPujMfbEdtVRmoJah83ruPcTNcfwuJAK8PLdtKfNf6Qbu9gS0pTnAg65c2R+V37dgtzBvqb89pB
exrZUFxkl1xtojZ6ssKBdogHo8C7Hq8bNRP6ZoDh40lgq/xExRpH5jb4HwEPfO/hGgwW4rR894bg
qdHaix4T1e4wtV3kpzeJQ2RZQ26Ouq+3NqWCnaSBCsS7iAULz5oez40x021NPzVnIQB8L3XSgGwX
JUDEfm9P9LlkSGWidWdNT/+iAwPsPRaXu7jI6EuysEswrXYMcOiLmqrNljNqf6FhXIqSnVU9pg82
G1fM202o5sQMUy+KaSFR73bYeckQSdqMu2mS2Jb/8kXvI8Amu9psPbbaigNa7fVIxeNBCU2I4IvG
pqCfxSLeUutEIT1FwLHe7yUOKYuymGEo5j9v9Rz3RK54any5qsw3+6/aohh01bX/VcZS6bCztbpP
P11BtoOU9DILLhHHzbqsYdW6M08sLaSDYRQHuCmTDMbVJj0ZpC+jLpydiKLi+GqHhkOE0iFvAxoz
lZAq/J+FukCDyxiT70EXsdB9iRHiQI4GFBBCRndA08RrjN3/k2R/5cdR+0VI2HeEphLwKW2fy1i3
sdB+HsEmeWcm09L6k4dxkG67/8bDk8PZp22/qnoZVpNnuWtqTOJq49R5698smFJlRFPHK74c9xbr
WEPP9UHPdBWxQX/uH7cB4bgoA88+ufZb4g48cwT8MidgiQTIWbJx/dVslZCjLpjL7EX2avZzK/hV
P/TiJtCqn5ZqLoDVp1j1Nka8s2xfSVXpWnRC/iGhjGi8Ne9i5UEp8bCHm5D9nv/hNHT2qzF048ls
6ed9vYAraVcQyfC77Sjevbx5zikOBd1sF5Z0KMiV3SGOTfUO6fD6WWs37gd6O8tixbVexCxmhNLN
Je1PHj1JOaQpTRxkyT9ESh1ZK37dwc+O9BvUJQp+8L/2dluN7Imk03DHNpI3AoCqdt3PZdLIgOKe
BgnpV9CvsBT30Tcl2+OyrrK0eqPpwIw6PcaHVYz1kQcrhMfqdqoQlyvrml6bvulHvsT7/sevS8D6
eK1pvzTA6jOwoP8ohhlN8cEVQDMYXLld1b34r3WFVD/OXeeM5IZLl3HtCcgn//hnVqPpYIp3pA/c
PIFYLf8SDMZIkyKLTFhioNrjI+qCax7OsWWMkGHFHEapMz3/iqe/u4e4en635HtBFsPN3gqGrzrr
+WcW/Psg9Ga1kCGvoTHq8qV9Q4bgUt9rHTr38Ry1P7zpi7rvDQ2fnB/cv9P8tzMzTpCBeQpY/UEi
3G53DgsQnZDwJrPI5v+CujjhDmAvCzTqqGBtXrpS0iLF4Zrt0NmKfzsT5oM1rf2/D+7nNd7GMV6A
qNfZi5xpWeHTcMEDgKoTV+WPSp0y4BgHMvJENGP5dd4Gukzx/CvK77wUVhuahtHanQEimgTe4TK4
PjFspAdT0w8TVxkDY0qxkfucOsTmZpX4SVVY8+zs5V7HpZwBHySRcDtHmAXrcI4P68Kh6Ne0kqvP
a54G4+EhnuUWUoFl6XegggDjA97KI9OBYLoCfAxcMLAXqzaP4RIOmjOkxW0dKWi6ymhxJuJJooek
kN2U9e7Kk+MQ/22Kp0GIfPKDmLJDJvihfStEQajMQMl0sboJcLLQoXRAwwA3eVVMyVH1QB3Mogt4
StGHnoZeI+0ao78jSs8dqAWJ6y4Cgh0uEarNeSQk4mGLbybFB2BtWjzJdHZNQDxrW+c2Jd9m8sa5
gOeC4UY8QnufZk6zRFUGZXu2JSTjjq4CH0p3CW9QIyXH1XboXM0tlh7r1mB9oHPYAeKqdi3nDCwm
dkzFKNCp1PVaVa3PAxIeOhJJQIUr49ZTgSBfUj7/XQKEaZSdE+IeLJDgv+ysL5WXl9W9NnEjIb9P
McgsrABE+acNeyLNJYGg+BeK6F3b4B0AhtbkIVb+gatR79WKnynvvRfiNsjkKN0T8QZb62gbQpm8
nP4L2CrqLhjMdMQNBmnRDEhP0oi+XGvc5m/UlSqODtNDEzs1g14xVTWg1z3/AC62qymBcw6kwbfP
RilYyf/HMK++/FY5QRHmBesIVLsExkpa4yjgYUBmQt1toB6fu+7S+edkjgv7bneRG4p100+dq2tx
RqMrAcFmm6D6Z8Xd2y90oc57NoFLmPmKltusjOnu5sBOEicalUon8hcbWNRnpzRJlXDdTSdUJuc+
TfwL6AM4e5K+N47OUHtl7f6IsZx5IRl3/4dUQG+Lcw3HZ9iEMm0dmup+Ru3IvdAo19UQ1Q1OthZO
HlFAAwv3ZP12C+6pWsu33gPJetFCQKUeTlc3OawlEWK+wey0OHD8k9wfQbAXSpg2zP9uYqe0dqp3
vPz33Qkal1Zn3ZvOrFI3cwMUeVOTb8XrCIj9TjhWwSg5Pw6ECJ8q/iKXVc62luBa2k9TMOy0CG96
nbm3LAihuabZCOv6iPMyZWz7McckWsiWQIuybm5IGZN3+xtF5uUxb73PTMa7RHob5JZy6s9RZWj1
DMFeNFwapOS6CFs/U78VoNIyxUA2D1mqzDz8Y6k1aXh9jOxE8n7Ltuxh/B+YKher0gyzHU/+tzSg
aoxhCL2PIbLEx/QMStLXMHZ5Rvy7j/fdM2cYo9/j0TpY863x8SMniCh0SnXDXiWjs8Gx6rSLrGNo
+jCeGWz3kpXnsS6KHfjnuKhirc3N1MFvvfSiADFZuCfPtHE6ZPge2QQXpetE8K51guetYJYd63IE
BtIbSJqsVJxDGdedfwkCgAHgZ4rUqJrm2uoGJfIoi1mYJGX5B9KXi4Zud+8qMbWLy9QYfEzYpfCd
YGrTopBDr914+1clyD/fn7mdiAqEi2OGxYpJeNcl6NfwfLYhZZTUoV+blNxU2aP9J0Ar73hHiUHN
RllOGFpkapq0HBS/S1gW3akES4ORiDrKOesxMicjPBPrTRK1UpGd61TRW0LBsR5mdVfnUgAJscki
maa7o5gf2XBfwJJBmchN2Fafd6Z7ZH2BJwSo29juULUTLugkL0yCvFWWM68egrh4uTOsw1ndVvFz
A2bpZon3Sy2totGe8Axn40KjVVO6+JDWqz7QBEWHGAdJMvbjYpS2gBBWgJMxwsak84i1OG3Vppom
HSwcaHKMfKsybcGjtIw83FJPICF/Wy2pS7SQthAA923qi4/rx/XElm0BlTDaPr1rG5q2FNs+e2Uu
QtmrQoCVgZGTw5Nw1hL43ZlIt1k3gk1qkJ/SJOGzSx3kZ9VRH02P0TPRdT86bDsaBSEk6EvFeMgx
HZvVilxUt10zYQ3k+uQciyi0kH/Rnd1ZlENETqL3dHY+eERJXXQ/yM7ofpJiUhN8CkNEiHKR1HCm
DUGDkXXZHf7Tj7FskE/8Ao96VG/e4v/HIiJskCHWqbSAYIp7ahCWeoAtfygCP2Y6zo6f/L003AyQ
+B/id2c+HOE7hZd5faxSBhm6Zl1w4ST+TsRjGv+WejG63I7KT869ZIZKzjm+Bawa1sbN729zSLAy
INEF+MiO0XAwQZT2UdQgmMsfMCFVUQD4sPGad8/dMdNYBeaqTDEK0rShvF+4xOnnKJrJfYXzp6p9
qRrwIH0aU7aSH7y4V9BTVHj2SZIMEOBUgMu73n/eS0CtAkvmwOEeNAjIo0r73p2AXEDV22xnd6sh
7gk2zhVV8neSi3fV5/+Rtoo0JXO8WlPAdRhwHQ4Tiv6fjMA3K4iuEIggFqpsMu8mTfnMRaN842wE
+/5nn4AJ+9TMg+hb1mx3ha+Qt5wFoFjJvRCLLTQgMrgxgPZsZUgH+2w5Lq2kLUqpHREgpyRLTnQP
msVBnBN96FcSIdnEA9w0nEk8E5yq3zIh2Ma6KPJNO01/t2FsSMra5T/CsHGdeXAdPyK3cR35pxAy
Km9vM/tT7apoSswe3PW4zDLrnRhHSIvT4qPakuXL4cgUcggYVK7gP3TRzejK9qDbo90t74OnWhDC
/tSI1njGTXO1ICeq66P1aWCsNzlu01WR7NhwzTj9xtp9+X0dzfvJllzJMZEttn4RxyqyrNtkY7ak
Q5pvqpLFnaWNFb8O8sfGA0ASgPp9sPbkpQqG5W/NPAUAviNVacbfo43CdJmaMmZgsGgdHn3AaQrz
M3XC1xWZ3a5xtq1/eOnBy/DkM+66XjRM04Y0kcc36R6sSQueZZ5Bh8j/EJFLdvNQcv10HAoZvboz
+Q3Js1/uEFcRJajwtIq5f9R4+mY5MXg99JzrUBMJdQrSk5odqRjVGnzJe37UDaZS9jf8a7aHsjEI
TQh4OyxQZXVV/wNvdsaeHVB186FvioPBTc5IGWHCAaWHKzal6Mgaot2GBgOY+fZoaMKcm7l5ywUi
/9SaudUbjL4f/Ax3JTwEckddmX5lNRx27bjp33vQY+WCz+6MYuLDPrWUS57bagwEsCT8nkUduwIE
VsVirOQKQv8Drs4rnASH1V+zWhrSRBGbdjqSuon36cVHGeyFl/IcsBl2SyT4bhIgfnWQt2G4VKGS
Fxed5ObtsiJ1rx+WWma/hlzSw+3inBzaefYgR2V+DVt0ccpvvD4Jd1BBGni/iF7Gl7Nq9nhWLFOX
vw1F2SDWkIWp6VqT3fAQh2iRTSeKMAoMxhnOXD6JE88C7gH3jAWmfuToqgjom2atVgSrx88LeFIc
jc+AIT8ymDDZjyRnJvURodpIVp2dvwjv5gUZotpy2oKnPsOXMCbwXcg0yLC8lPlvzbvAOwYTqypm
0cbm8cY4ChH7amG5I9OKrWaGbm3MF5D3kq+qftbq1LkiPXak1JxuwGgJEPXeosESZ8S7epbgpb3B
Xa4KEQ5vWGeOuvXerDvcDcNl6NKVok5qxSXL2u3wvF4lJPS8FSYCi9Nor/qRjSUh8fAeZKCvcA5B
V3dm+DLL2jze6BvhEDWTaKPY798a8UbkYVew3ifNUsoaWj4PR+g9Jlcye9kJoNumDUlsy3db5dFN
WA3zBQ3G1Jqr7X06hbQDQlivAsxOJWMX7bEdaKNEhSJEQMDiOWW5rZJnwazQ19rBHKa+la2QU+od
0Q83X5Z3vrppFvEgJcwF4RM6ppbtm8xwd6bYjQ6eHD/H5aWCfPhq2akvLwMYnR6o7qVpniCq5m7H
TJGRln+xkh+3cEDbIOjoHb3Cf+MWgCt/vIUCQZyywkUmu1eq1OIFSjCffKy6M9KeceXma7tUcaIv
L3SxNkHALppagFooERpX5v9zJjH1CN4FL+/l5w75Z9+RuWXbyXz5TtQKHL0Uwmq+URq1mp+KOw3W
q2lLj1YA/4FSZxPLuMast7fI+o6aXaaVi9MwnZEse5BC+6aXh2+IS/z+hQV5zKLqYp6s5R7tr7Al
G0IMGWI3JQoGd9b8N1ME+H6REvHAMVX1evEKT62dzs+J6VcWFow1HucMOB7vD2Wix9GDdcESqPEH
88OzwQowvHXf2/lirt/H4eOYxWJHYBL5VF+gMvh6UkNkBgKVyn4IJj1wJFc+OkX2KZCxTGbteTU/
KuJZhs8QgAdw0Lw3vZ0eh2Dr4x/2tkzqnsBIiwFrB1kcbFVxWFYnG131n0LzJjiuJzhod3tN6f0T
Tyj9nreq4hCSonHgKKZq5FBekUISZq0ymgwiWTDB+kdDpozi8vfCA4+vk4DnYvXhCVDB09ATVugd
VCXBJiYazBz4XATQUoZZy8HaSGhWUtezhb9IuVNtoPRwN3UQB/k/82U4F8D5L50Qh4/SyIAC2mfZ
S+IuHdKYFZ9uzol87O8WUF4iPiKYdki+g1g/0lRpQYf1hoq1mCfNleIPCb/LncskU7CfyWNORJuP
jcV0NrOP18WZyOIa/ObEsSykgQ0KG82FEhrvH8hL8opVhR+PB1Wo4we1NbwlZNxHXdDzoe3WPNYe
PaD08Z5hCyCfJ+t6iSSF4HA1BHIy89olJQuzaNsVXRm5KO6NOEyVcknmRlZo7N3Z17VRnSfAY9dF
olC5rUR7diXOqw+K6BYmWYT8xeevzhJyG9QMTRK7SzIGbp5VM6NGuXBgxTxuwiuKnX3oeg7TDT4O
WNBFUXNYSciHm7QwUzK2pcyEbzw5tWrHb06ugn68WXXzYCRVQ6VGVF7Ovy84mQc1FaWZu1GVEod1
RHjFsbD+R++yMhf9mxEliFerLivaSNNPcGKPVsmopAD8pchpVQToDNRXhzhAmb8N4/d3Jv0w2mP8
QyJO2wa+mfv6t2cnNwc8fwTWMvnHx5baLLVpgcjIs0YEEnexJ9xOt1EUstaaQ0rll5rq9aKGGQUX
DamzfuuGkG7Z9Wvfe9OXS6by3S8tH1RYHTAKKHQEt56USqXutMiTx5H4z6m04pNSw8XhO4ixV7jM
EEnLl0RRuIU/Z6hG47HwAN7dHfrZ/dpd92btqDnU8wl5+6XRh/A2DxJiN10RD+ybGu35HslvZiwx
vWeSJ2HJKi7txyCDlNqKJ2CCGA+fJaQmNKyf+hbAoCZcqiHNwS5tc80TREnKKE/QrxIcq728OUkX
qcGA4CPfTFNQyK808yhF+2D0IAAFbAAwXx0+0vdVWIdHdsrwKSoE6tNmNDSTb4wbrMJD+5tvallc
QVTlVTGhz8gMNTUs08NAtIMXnJ0Cxpjtk7+O/oTwQXkXPrcAGsbtffCEZkh4WZZvvphFBycE1q7k
lv/apBvPBksx1AGbni/Bs27QAxUYfUHDhxEk86Nqq1BUVe1Vvdutvc7yqYdCy+XjKF9LLCEpAkiE
kz8pNFwKTEA1G1KaQYHSBi6IrczbZMWtzFFebnZq77qE51f4LERTwcn+uHiAG5AS7LIDsEn/eEmt
B9bCwzZvLM+xfEhMSkulKFRRo1k2QsUFm+YBxaOKmRMgq9HDoh6Qh6rZ8C5Vcs7n0Baq0nsaIY1M
68dm/e3rWidpPgEaMURCmWqKwEzMB4Lma5cBfvaLKUzubYkAG2VkRiAXBiugSQxYsWJGb8pkl80j
2CPpy2heClT9NkylAzVDJsnFIuT5BEjP+NeIb8caYXO//B98mFSjfd8dWEztGEwsJ4tNkCiunfi8
mtjzb/f/reFDzxyAUZ0xduiRlVUVM6oi3To2BY6PCVw8zYSMmUNURCoEbYXie5gFY9W+At5+Saek
JJXYijS3Kh1U/ThiF7BdyEQJhy7tJlNrMrOBotNzyAEqZPRyHaCDUFrzZNsdJSUClo26pwYrg59H
Inp+TShZR8ZApc2OLCMLSelWR3IvG6Jv6j+sPuydwENR1t2qeIS51R/ezkZ5+ML5WkRMuIs6li5h
yB/wNVNSrFpSFQu+fy8REDGBrSRXdR91vENbOT/bJOTWkDQl7Nq0OqPbdK0kIcNuJviGio2PHDA1
ehYUz8oY6Y/1mKhcOSUQEtzqV3moGxTrl1qzMKCYsXfhozJq0WLQayc8noYEvdrIHsipGgh8bonH
8Wvwb9S+gdsU2z6jCA9EdiotNBFqwEfdTDu9nfQQxq6XJm6FKHU2/bB+2TpH38TXmlUM8AzRxjxC
aYYrs2JOyqWZSeOqikJqhdx+M3E24h1+K6Yjlh2JvtsG6NWGkP/+8pISJgMQFhoktB9lbW4ZPE51
cMwv58n3GlKCYb+QI8mC+2q62soQVg+T5gUCF517/IvP4r5Nb6Px1IQ0gHUaCCrIR/5ggkcHHrje
0bGDMgtdFUjWkmmzzT2fv7QCjdVRMtKuSP2VxZelTljRTtAjnYO7bLYNk7Mh7F8Fsqkcv6FFGCDr
H+aQEZ3ljDHAPRme6jIQIqrPR+boQlD4/anwuyikIQHLkqtTIoWmUMXcAhn3NyAsD/itJhA/7avV
uJSpvXTikWIC7sNHc4C5YbjYkiSQ9joxqmD40KLK/wWQRdKNcOHGbDPG2Ea01+Ioe1Tk4mqaqj7K
HXcgOvVimfB4lLjRTFM7NasesTZUBPdjcff4+WAdbyvBSrUzGZM9+AK3ltpwtFlayNAL9cA9c9YF
grt9HvZXcxbvbg4kaHIkhjHSSHr8Ih2i1Ns4oaoV5VE4jIP/nd/1YFAGwGuNtGyTl3cQoz2IHpz6
u6VSCF1CouaB8Mg077UwFQoHao+FK7yZEOdmH0x2p2ZA1T9ULvrtrwiGOfwP7zyleBOsds+hs3m6
WsNL1yqdpnHeqyLtTa4vtshjc13bR5mJ+ce7yrwAiOzCoFmHVpXpxBWIergomgUKK51maAZ8bUTY
cU/EF2Mfn9UgUQA6lwycKA9VEEsAI255rfs3FXeR1AvFuKHQaVwtDMYa8GTMVWYSRLnZpthteLIr
jsPq0YzA2+aOedZqe95Ha7rNvnm5Pxt8Eo3//eVuVm5HmGv8WMGL7kTJU0mL41kFP83ANVVNTr79
XDJcwsoBZ2ft7OJAZfxfdDDBK9jcHSLieV5jZBMt0sFPQoK9pa8HKSkQSthTJ9HJbDhL21KHqNah
XMBeqtZWy7BN6ypcaAfZR3MQGEXR1KZCXFD/xpoRkP0mfuvVBvoXlhK+gv4Mt9BH+KioO7+V6YKi
dE/5o0Q0pTkDnC1NTcmsOkj+D2+fgD0tMUvhdRbJ8oYMGWurAOocwbfPWTIv1ibQITp3CERyjrkx
LZ10hsf3H+jQh9ZVqQqZ25BIuYGxXd20uaNey3NBi4QBSHCnnYXChEKzMb3Xi7bXN++MujT4/bXZ
TBy07H3P8qoeiid8WFLGg07KTQSiK0QH+XYgTn1PwpfQSRtm6Z48dvJwKECOetKBW6O8TxJm+0L6
UiazKkFappXpZTSTCZp+vfepSD+NOjLoLv5wb74UI1pEvmyuiORk7Jm6QfX2QkPGhUiXAxobK+ha
e7Gk0ZIyQfiKFG/Lwq6QAUs68V9EEINw9MeLarDCOXZsgIoNKe+cI34oiU5FkzKELhDEYHgAmXXW
YrpvGh+4Urzjw3imUDzykUz+G0FNPBhTOUwuTvOh3hDquQaHcHzMqHTfopAx5q6aF7C054iYae4D
NFRM6i1Udf9Orqhmu/JQS8b20nKeRFkN2EA4hUX52dT5LURXRfo9nD5jpXVyoRGJLar4J35wC0HX
B6y7ZRKniZwAI3eO5Z+GNwIQbTW6c/7oESFkySMxl79qh1Uyv0FKjuN9JZd1kW2GeAk3jeK72Fgq
UMnhTrOJMJhI1oMyC5Cjvla2pZfOk7e7KCTvPz1TvuNtYdMTfXmEUDyGPkNhVwqXUJwUuzpDGm/r
A2AyqhIOAIcgOC9I8m7vR2zsFxZwJMRk+OuU1+K/41Cl8HHfOkysNS9WlyRRxRNIOZcmZOHCchl0
pBbdM2jY6GyXgPJoELrgzLZlMapztV6fDi7gcHU5ksp+rcZcmlazGBd/CgKCvveSJE0vrH2sdOj2
56TzlCQi0twTg37XS0qWG0VcpqI2R51sDvBcftRxdnY5DEb1IVwwLeioXeZdd3v5b6WBBCgWyUVP
iOt7KhsKCXHdIZr3MFna2u1pid4knCig1uxir6lPXgMGqho4ZA2UBPCWtKYiCGxMWy9+FTuQQrWn
7lDEcB+g+UatmoVlQGyRLsw4VqTrxmymtAFd0PCWPAqs6m4y8dPIDwig9p9irkYfijkN9nGrZxD6
n78OMEFfsleRaz1Al+UvJv89SgvwHVp6qhu114Sw0Ckjl2rku73nBAvjdaJy05lfiMOkpI4y67JV
aJ+BymM4TAwJwZs3exSsksO480dTdGGkoyNLtEAw+HWA0Brs31d6zm7dMtXl2wMhbL/NXjVqD8x/
rJ7M5URrfymZmcAEswCO3kcy2JF9BgQTlqIxtJssT6aY984jKqIg/kdleY/9jZea7N1y9o3ZiRNj
eC1PMtMrUw85ue5pldvfQf73jIZXiPSW1zXJrO7e2H0PBbEtJvH4PWXq+rwOI8e3F6fD3TLiwsUE
cAMLdJvFu9CSrtEpoh+GMzIPwUo/S9zYEAmFNKrnO0MnRsdUVri1kvBIOTI+HHE2VnwSjmdOCYqM
CKfnVfapx3Aq3dYtrri306LtlQ1cNydEYb3e6BKwTj74OwbP1+sAkImIU3H0jxN8VcbfIV8y1MCe
Puq6CLkxvDxOvw/zqQdPnqHT806Y1XGcXkD0FHDc1WK5dtdpN9xG/NatOpSf3nLaTQUERNWkPLT4
mCHbeRtmlKfnM+YV2s7d4cuAqnzKBHriSKJH/Sy8nzeEMzkwFKtIUrCTqYz+nbkS2nf2lW7rNRs1
9CjoXCJSrdImJfXQoF05VuL9ovFz7JPvINXc/CSDzcZ1br7P2TFp3AllXt/TJLbqqW545kcpSTE2
rbsHdISKclF8PejXsxRwpoPtZHEGcDhkkGXuCtPpygosWkLAgCTGUu57x1ZbYS1MzVZjKRO/1vZ+
Ixljtw8HJ6U4W4yCneIezwj4MqNWEvzcAyPXCrYmt7KavWk+IHsoII/d6EERHs8Vyn8+rNxi4gxq
fdc7nz3Sz12hU8rkdrouAvIgFuw6duLEpnWkgzvLcQ6IYMCqXufaOFkB2+XOzM6oBqf7Ose4tzXC
SQ8WxGdUY/4Aomi5hp427fbCAvjL+ME0G8I8JU1UVEu2CcXpgKHCBV3bXGwHC0ArvW4Jc1cmSRXv
laXhJOBVRIE4bxKnSKmyTbOU7KWX5X3JCSK47W23Ju82fgHC/Uo1acwCBvdrVb28xpc7bNphD+uW
Q0Fr3fNCq7I8SJeXfXBg2G9BAdW97RY/eF0QKr8rBQSRlUFiZlDACTVI4LDMNVgdygqpNS8LFBej
ojosj1bCbf4C671EVWboGOMnniLPa2b0H5cxZ98Qez66eloRR+VVIRG4eHgwZkfWt0bC+UIjd3Ij
Ao8MMa/l7ZgrKhO6coWbxb6aGhqQFY0QBuDpb6I49TVeji+wdgNVhs6IbCZ57CIz0OstGmsxZMDL
PE6FOJzy0t28yyG2GARhguSoWr1h7XcnhorYBS0m+mp4APi/fo5VoW5m/hULWFurfM9Suzzx89FV
RC0R7fYq47JOBhkt9erqjNbmcEr0/uJdjDsU6BEmrCYoqJ8wACp/yUiE+5m5g1Y+dDNsr4vQf4ua
49et3jcKiZSrkF2a/rF10DL71WG887Q5X3LJ+3l32rqdyi7suS50sO8vI6lmdOfktVY5/eu6ZJWw
xQkN0IQf6/SAMWeSTI8C7WsQ2UsAd8n/bITfx9yuAnn9mzrgHwGRde/plDmqG0JqGre9K6uOcOhG
Wzd48h9Yx8DIesFDmcIqJFBJVL+dO6FO/8wAwY1kHicbJobqlSHOgEX4Y6sRfX4Sxpt1uylsp0fr
SNrTfSZ3tPZJSnAasX2BYeYoJcfaoDA92kUTjBCCXeH8sIa3B7xNjIGZ4DFX0xClmFEYldBzVIem
xPkVpPr7OXDNDrb+V6aGJEiwx96C10kRT3dk6KBVD59wVMNPq58p4U0PN1U0kP2NVTfZN5MPl+Gk
JxGjVcmRwyvcJeJ+mcHKQFjTbhxroCQdvRWpVGWxWjWUm35zUdS8mrcOWRtu+uAuWOW3Rb5A0baj
bMdOvowCaicsgrls+n0+jOwOgpLFnlmSGO7V7u29gnEAu50g7q2LAW+S4XB9XQgfWHWL8mDaNpl1
oLlYK5pqAblTJTMzwS/qDarto5zmxRn4ZrJXouga8BDMSqAmqTy6MFmO7x2YMYdHFD5OPBf/klSt
pWs5bq0hLHW0ay31ah0RhBiNy4RJeWwJfdSNKYg4fauZ7OkbSda7exAnIyWiLXqF3uwFO+mgeejW
XBssFnoNUfrhk6O0O6RYMH+kE3liv+WVRyx5AcLYSWPKtPKuu2Euc35/hqAgc2HZd4mT1oD0J0pW
Gx0CZK1MRn/NoVAUL2VaTbAy50bB7yn0gPQ2zppHCPIhZccIRfKHi2TQTKDk/yhrROjscGT6uW0x
7k5kHPmvCdP1GKVVuk/QZlqJGbHPSBCOmpEpybmiYLUbFaJhx87Lx5kaGtYcxjExjUKJM+LQQT50
DuZ6W3sWWThXyF2itVwFyoyJ3kzofuBq6UWZCeOdWvDm4P3Vb0wg4rbe+QeA0d048sBKa0eTYgjt
tM4jWy0+N6sL02I2pJf1fbTXGSZZSEegHQ3ROu7AuHqsHH4EaQAg+gtsniNJczvoO5or4G1E+d8q
ZTvpCGLkW5x4aLiwfLEvLRSXc7hrucoCzVOtZkQfCNEY2QEmC2Z4qLHM4wS3/1HkWjjrzomOrtTk
pzdLqhqyxBtjQMGyJ1IxZ/Esok+ftegc0akFMgXFT4iyTtuVNkSVAhGQNNaOxjZWLio8GK3rl/pH
/OzYi5HXeE77VFKP4Jv/Rd8+CxCTdZaX0YOYUfRO9n2FC1ChtdPcHCEuDIk6acwdg0YlE0D4U1L7
9MLpYIJSESRWtHobkC0fVkDJ6riluT7iqnX4Y/w9TYpZA/9RqrTwuTWDxCZt//lXpaMdrdipdU0j
vrsbkz0kF9lyMTtTRGj/gES7hWEeO+DB/miWzKz7UiHzAwGJpd9XjeCX3VBCd3FzJ/2bPmAZ8qWB
cLNMPR80z2oHvnAqTVvMlnvPK/c0AydHECRwbILBwzm1gU0ZLbdcY5Ar6VAoWJkjrUUQlQMWcpDi
1MHKUW0WKlmWk/H4p1/0uf15qbT7B92KjqUASe96q+tUR49bmrgb+f31GNZgqHK1vlOuMhwSqhzA
GYqWZmT/MKFiJdvJ+NCX8cb2383OBXFx39ngczRZ46DDhjKZusdhRUZuk6OakrnlkSN87r6u4XBK
up6HlvWdBP5v9yTrYkjXHkV7VPB3Lmr1nniryB4FWORjvk7pcL7x+Id4N133o2JoCV6IYNZ73r6x
ZU6lK4O8SmbCyUnizU+PPPy8By+W3nRHcsX0wfKsSzhya8K55XML9w41cgQ63qJDgyeaU51B2Pbr
Q3PsKe95TaIrEZMum+C+3BIH9mEZ6rdLVOsY+WTKDaLHZl36DM2ncv0BEkAzmKpndkeZEjK1tnLJ
AFmPzEwvpWkiH/DUGMphlH0DW1LB1dYn6JJe4TfWpiXMTVxCLH7ov7IkImiK6ZurOGqF5z0qQrY/
/Y7JT3D6RU5hDD9KzUJW5Zi206mYHTthX0hBl0i9fm2+kv9uywTR6A61IYJJmQSVMtVX4p1iYhC+
RrrXNHohi/6h5OkJ4OzXkrQLpdS1a9W4HUYj1rC/KBuoVHfyeqJfGCE3ZFCkB1PXjaYmpaKhhdnK
emzGAmf5ZYwlpA3MRqAGyTA4FyaHOa9hS1+jdURWzm/7r3O01yahxQPbXJKkbcxDLBc8fEAPnnb1
5CU1gRJu159IwWj0o+/2H0M/CSEfLiNIk66UQiITmbbiIVPQj59bM3VxpRPgsIr+UimQS0ROvbhZ
fGqKEctAgDM7yC8WxneRt3wuMLmk+XJzA7o13pti0078lAOwu7FZBIbl7GMz3/dIO4QATS1KIqGa
Kdz4EBzgaF4dQpdAZtptreZG0g/VfWiYs7z4bi0SC89C1gOD0ok3ht0LfkgK13KOf8ZK2ob/9tcF
/OFamw3PJBLzyNZOx2SncrifmktUX+8JVnf83hSms+cj/nt5Ka0wYtlFUwd0ru1AW+dc+SQ7tEl6
LfRLZPUmoSmqLOYp3YDHs36yQLtZvDO+24Hnn+Ga1X76h8elRRNrzrBPRPNUlyr7XcMK6gPNaTgD
1zJb1KBsT9GTMsTna09oxx26PgWsd+lZSiPJly+aLvK8OLMqHwWkWpV9czPW1petOwozZ/eYXyML
+ubOlAeRCkYxmCQ9rL3pENnCAfXCLNcrbYIzEsj3FMumPxtGltYgQzK3JpEdjpOh4QzcYGyparA3
dWZtSPwZCxS4WkcB2S6UWO8MrCpVdLyHkQxicf+flxWf40DwHPCGEtCM3bwzyCwFfevheC5ZPZhW
QC5cN55l5A09H0FVocDHCpjczPF9t4zXNou+6l1DKn7sNuY9oG6vo62CgN2bVyrCsKqN4nPw0Uew
mLF65tLGtvIksus9iVkxuK7T8TyEsPcX1DEUTgNj0vUTz1KTL7xRNgS1g3Ug4r3jxqQn/ENjyCx1
+H7yfwArTeQTH3ciZNNgdn9mWeTycEUUcWD0uCWxHJRAsyr2ZLZfxICukFVJcRqIp7xwYwo3chZA
7kyLRPUp9dHx+0S5DV7Pecmm6pNUlhw0uyLPl35J0WAMq5MTNM/XCnAaitd0dXIBPuZT3rxr3SQy
TrbXE5x9DN0c/tS7ZCkFmDM3si6lNcPEpagNKVSctSx6vnwoQBVoCDyAQi74AmXtJZDfnP5Xqk54
o1qWS8esOpiP0AuygQ2fTb4cf0VsffqVv53vjWqEnyb0iDgKExc/JXSWcFtznQVTCYatANrwrdMM
wvHHtDVWGioQ/ar9tJvEo/UE9VLeW5b4kNTW3tBzNZ2tJGRlmoxdA4KubqBV/LyJtyT9kSfzla08
0LBw6MSyrUSEWEdBxggCGBdRq8pgiZUPUIeRHsBBitROMQMwv1ME9m+JgV/UUyImdcfWzp4fLq4E
douzJU60e1q2/r/Fs0VUmSuolr2EtYDRrFzAfuhcRAskUHVhQJww6fewORuwBYTGEhO54fdkPIVG
6deRZd8mSVYxsLhAbrukmfyPidQiJ4OIuKbDst+WrAL7wvaDQnO1WXXVA0T42IOMVAc6ktOqY6xX
kVWD2zHY8+pcZheBoEEMgMbb4nORZOdx52CC3t+kc6UkVB2pzR9uae661k5uWDP6g58itBg6djtK
PhFzHsaxgMgANfcFbg6Ri4s4KwXC3+mB1S3HT8fJTd2MSaA197fzdopCI3IAxb2HfEReBgherF8q
hOqb6o3P93o8sUnVVrz9jxh+JrfGiqB1kVwE1M0JwFDNTfkHsafcB9o6gh+skjo/0NZKGqt7eVgi
vx0etKmBj0xqI0h37J9LWww84c79XN3xEv6HHTvS07EG/a2Y4EqWm5OAfGZDn0WDSCW+nmGH6y6p
3NTyYCITOXj0hNEXSTrtF8ddEI7J0PwXb89WYNQpnMrtKtK5LU1LYBUSFo/op9Yh76SwVkdv4Km/
pI4M+5l5qacz9artw8oHFiWvWsrW7cJTzeHuzsarbF+twOkIF58piRrBunF8SqQtpzDEUGpVS24b
d/MY5iUYxYyNqISTy0ajvf6FLmN6x3m8x7+BycxTk2piK5orhSXOiNz8K0y8WNXFwBKrRIu0iJv7
BAeOyYt/JVqylY2G2Qr/p+9OdooxgWnHISphqTG0NQ9LpxdGUqwZ9/9RqzOsTksNyWTlqiJMT4M5
fNY4j18hWfBhaYLwEwGs65X1EsMfVBXM2pYlef0UDyem7zB80XFlAndAIMiu8YSRaqCNk15tLaKh
8StuVPpXeqFgbVNHt0AC1gqEOUya1ndeOrI1Jrqhp3J/ENEq4hrulpn2KEx3oW+4lK4qPX1xDkYJ
xDHK38/lXcOr3XiJLpXSQbxymirphCYgFtsP9l7rxYz9ZR3PVjt+e2G5XeCrwcAGcrOF/NeXsiu0
ghQeMwQcZL12iNQPMgflztlif9wAk4BFTgyUyyuaVbOO2fCtCAFZ2BV9GPgDK5bbqr8c9jQAMOzP
bGJlsY7gqrzf35i8BxYlV8izcJSqneKrEBr4dRfv31i/S8gYTFz3p+lcdcxjnHLRPRUfRs7lKvJy
K2m+63G2HVHudFmecWmZH4fhLyqZPLlUsrPuxv1u83hLnD+seAWCnjrnvbqPVUghFJ0JEE6euemT
+8boo6Muz2AnV9yiPHER1vjoOuHoZYmfIgvljXAAfypMcwoy7LOnDsp3iSM+uIezgzer/7gMF6ex
zJNjCHKRSxv7icy7yIDsMSYzDXrfptSgjgnOn4KmOk9i1qNfiEP0AM6+RiRvlY8wObfTW0j+LfC9
/N1N6fJOby3sqnFTJ9kxuvu0l07Wg4uVYjMhT8EIhQZNh6et7deaj7O+h/BEpDU9CbfVZKx4b5h2
PL6zFFZnzdteEsKJ8b2OFUK96O0rtboSGfp9ys/IBTBKNPOsUjQMKOTF8NYjyg0rbO6zkAzxvuTe
90g7v5mBF8Q1iUJZl30PCJny4PDqcXK86R1HXPetw/oyurlodusG7lmF3Bq0i2yahpwrNGn0HQEf
A3br1XUrTT6ChH24TTkT/JPdO8FtF2ljKivAXL3Pyk077wrmwcVhgOGlbOdPQqIISQUdkurePurS
NISkDl8amhu2CmV3KP2scs4Au1SuiBuKrbDFu2g6ks1UeM4tpLGRJWSQ+a1ncq/TPtsiVkbT031/
+ex7Tj+ZSB2mzfFx9E7Ne64ldF6p2c18wU/IeADAw6/4M3mnMQLFO9Q33wCM8BK/6dI8oLHPw9tI
fAevjDyPznHBDLlYVOGb3Pb80JklTNt1/la98j+rjeiMDk4AbSJ46PVgFCQrvj9Ny8+N/nG8MupN
l0f77Njgj3awai5Q8jiqqzKbCXh8+sQGZTqsK/pot9AIV6JOOq3ylHW9WpDDs+L2GfFkbPOTo8j0
0RYeMA+jsijShsoRwwQEd3JRIAV5pwOYgNGqMv9TxFajW9Xu0OJ6qbsUM4x1MNNd27bzPOFwWAoh
27i3jt4ZDcVdbrPNR++6rU39LiEfymU21NMEahyC+SsJZj0SBxdhzfGZ/1ZYhun3v+4YBBHTlkgP
wF/Sj2ZPurBWaODh1or0H2wXJlkwzRQsnumVe2qhfkVqLK2Ktx1VVHhkojvqoMGe25VVzyA4sjpi
Y+rMfapRQTsfSGK6W57lHoconUCLlXh5gAeZekNFhxj8QpT7HA/hLyhivDvh656+VVE50pspdb7v
jziTCJ8eWJugoKM9qPyy+N7xmO8t1iOWe8YhzRSGPg4pJ5/HM9Sv9y6GH917nPwiZkIiyq/mkhnO
i7cjG2BsKjHlHjFjJwGcWu/Ls6PMSJ+Tiiaut6ZBwchIHFvGNVXhlQuUgXevf3nhSMJVSh8Bv0Gu
gTwqfiCbhXcySpF3AqFi5tAQjgyNT1lD7vF8FPGbf9LtZN7I6EAroxvwlPPe248kLF81djU4Yy3q
9oVvmhyeGE9k2iEn1awvKMPzF6Lk0L2spk0CJ1QXmnN1j9WprXTyXo62yrJpWeKSSEYW9dpKFqOC
7MEosPsL2o6xDvQ9gqVPkc9aWTECAb9NxUB1YOL3V+mekHLROYBo5ob0cgNpS1TdfyPCY8f0P27d
Xr4EL1H0CaqJn3b6Fplb7Z/CD9C6U4s6sNzCxaaOYRZqXkw+ct11kF1I5+FrxI6+N2DFONR87JmU
eVdFf5c2lA3Lm+vBcKuP53l4eGrbACx2hOHS0psX6HJEMSC51iMFEh4UrYtV+vV3GjIFupJutheL
MBKmg10GSHiNV7NldzWym4L/oDPVIgdmwtPBhAh6EWCK3hpJ56XghBU1bJZQDcvSx/9/SffVi+xM
YWYqPh1n4phVzaAlmdwQghWtxHT978DtIGwq6Qg56hdp+K8ZZJzGMxBfstrDysPrtVuOAf9nP2m5
ailUrvcnK75mwo5OvDugRCq5KYFys7xVESjSwFLhsUcnhJHzUp4YgWr8yTwCOQvuQyvpnKT9X7IK
Zf5JSu2m64Q5hiqVGm+vIDZbggeI6XtddCsrUTENHod/vmF6WiUCsANpeFh7ILJKEliYklZ7e7mB
jRfMQOVGWMZhiryegf5gUrsVLaZV8DIiI5WTkUrqm2GZyyQdR/WBCycqNvEGLJtFyv/YST5T5Yxu
yY673FzipIXBFgOTRIM3xlVqaBHD0cw0SDrRms9l+x89L3PRpQgk/HzzdFIdQxI+RJT8pttJYT4q
vHoQPiuLOLa87vTycjXT1sYjpgHWjgs84U4LnqjUq6oFvC987iVBEYQ8Ow2FwvxtM7H4ylyu66St
L09ODsOu16EBOaYa6MUtE364C7dCX0UehZa5aefjvRgKK+HrnEayT6UPnn2sHb4xTA8nA+zb4aKX
HQDVHOaUORIrJvO41qIl6AsDewVLvb5/ZTmK5rJgMn++yDopDRu27YzBJ0PTcwrGbsMpDBAFkBgI
PqBHMkpqJ8s3jg9cpLMLZcv+ikILOCfwX3MVwadlSLaJcRf+Z3d6FmEcByIYLvlmbIwu23BytOpU
aJ3+zytiOhp81cEi/COn1E8Fs6bllWmp8XBhXosgn0l/Jqfc63lYK5lcCUmFq8pPVFqvfbCTAQN8
aSyr9lYZcZCa2XnlQBVauZqlKI9onxEMF8Ydf/eV/aOc+Zxk+toiKb7LZmSg7LaAz8AW1qk5JQMa
cAuTqio3pWKxyyuFR7ecLTf2szto38bWI4ewHwInKZTFhg9k+VsfBp0uDJGoDdvYcTBgFROs1aex
eN+42lBDZ+GuzvE7szundQexy9x5X5PuzjgCZ02OSHc5tbOWgWk5fnaRoVgSe/zzolh8ZU5BAgK8
sRdtSFoPxPMHii5H/7dVdq8tZUhcrLaldPmoRN5jYMXu6ELCt91jXD6KaElEgXIzKs4Vle2wpBjg
vQDktihuW8aj+h0tNOxhU4jtqElvNSqFq+aaUIVMzevr/Ob6DCn3eSYB+1zf7Inv1W9MDq/RElhT
sXbtvaqILBgrbsWQg2uJMJ5eY4yavecYrFokjo8uF1KYP9CgGeeq2IL8Xa+6D7hwIs1pQrIeN7SZ
UQI5v8DiXhaE2FIytGHKASCU0TvleoajK8ZEAPZzaN8xgM49LqB9XIey1btwZ5YAvnUuNuufgo06
yJRwEossJNE03Q1bC/gcq0MsnMRBsTxBXzSPcoiMmKuhJR1MZQd7tqGyAHjZbyxu2oXe4F25S6I3
keC7DLoFnnUsgYCjWe6pNDnlTIteWKeoPvcA2dZ/lJfGAP1ZlB8b3LfvE/S4UyX0OJzVQccWcH/w
VzMBcfpD7ST/IRM/DuM2WmHAuCyWO/S8WQIVG1MYNoXi6WgI/goWApdGrWHr5eCF51hh6FTc11oJ
i+3slpKgpvZGerfNzP5j7uA+Q9pn7XT5+u8oFsFEHO5faWzvMXA5BtJzpF37PNjAdrd3/fCSANE9
F7+H4k7jSzesZMcftYmx3Qd4fYjHiDdFRiCVXIrrPzXApbOgZI5PmHSId6K1Uzn9Gb7TlIdjCSRt
9vEb8/mhOsde/FC3TZYMIJQp5Q325VTBXz+wBoVX+xMDAAAPNN2syCceglfUH62rQqLka4AAtgAO
6HdXA0+3rkj8sGfHk9GZO2Mf31k1tQBiAS6o4faKA5UYXKBBbD1Vrl6z/em7/SPF85DPgnF+dxtd
SPbtd6+N6LqGaWjZz0RXUphHvl/6qvwwBT6u/QBJmMZlDB49ikdJ4c56gd8UBACDs1MGkO6VYhbR
hOb4eN40J2lIAz2fJmumdTyUmrr0MQj3QhoByOorHWNApi5Xzkx8DozKjexB0EFnt7CtNvtiOByQ
XIGuUTZOwkET4k9wYNms+MRR6einWpBhdu+4HlqfV6ZrKLMgLiAe4aKbcru8SplW5rgkkqaayHKz
h8jgMq+IZuClBkOinJIUtCSRlDLZK8WctTooGN8A6k+JnJ12vkH1a587r6XqeeMzWHCLtLn/0HoT
feRS4m/qJ9AUM0s07y9tNE4ljirqbfyhe3umPa9hWAPxC+u3NB/jDEhXzxI2xpSmuakZxS7ZP79S
NCQ7xX4jpExeo4LyYH2XV9rAJBUdPDXPGjCElA2wIjdwnxS8Dg9ycDDG8Hnm8jOXOr+5Cn4cCcR9
QXIHStvxGU6WZocryRF4pCbdsp48RieL1za2tXDcUXNhr6SkgBGLS0MZl77TS+M5eL3/7Aaljnks
I0i8Qh9yG08WwhIL7qLry1sjMYOyL4nwUyk01o/s4sAcZZIr4w4shVIGXPhABXFgUZBsY3EeH1eP
fQUfSEhhPaqI3svABmVUe9y5jbaRLs+5y4slbwuP4Lyjuuh0nYKl6zhTsv5LYPimZmyg3VaUyEFc
vzr1gOCAxN42qKSrt+js21xZO2F1jC0L2wgtfRD8sd+JVrAYwaBoiCE6//N2ojUZ+TRCPno+n9al
12K8ohWDj27FP/wahWby+jCFCYyljbvPMaisNKX+VSiFZDMMDRqx3AtGcp0+jvtmQbdDnd9tEFyZ
gnHgXCplb92xx6bBganmrebAR3+OxLLyNiweTLdknCSqIta6hLYZd4qgdrdR26Qn+VmLML46XP4E
3rW/gkh93GDZg540K5FMXVh5dBARFGtXpCSyW7SGVKU/dDAQnkPCyzou4OfrUJHAY90yLsw9E2oa
x+cKQrlHDRV1YB8A0XOynee2e+MEuHdCmft49HVKTVxqnUrUmkWyp0ctS6N1NEqXJnG5RoGWY1yp
wbClxgmy05GHclb8OPFVVwH0eQqp4WARrCF2zxxPyoZz2eeZ/5BfXR6RkKqeHUqhsicVVYBKgbtv
f2Vbitsxi8mfsdkdfzfvGkbVvptx2CVrx2ycrrfTcWJbOZlGi0YPb51UkL0BprSIGtyZcOripBIr
vyAuIpAqtBBoCu9hqw2CfW6fQ5KdxulEYX0RbD5HC0nykiiSycPjXfxIYUATxR3pyfe4LBDER0n3
7V4UHuxKzgo8UYZnllEvb7VH2dHVo4a4MHfqt2PN5p7/3jU1e89EjDakN5HnO6bP0E4sIIzGFF1o
BOloG4EnooAHuhw+BJg9oYJoiUG9gTbyCqn2yJPBbr9NIzYkhDGPKyMoGktdTAQ9Y3eu95+p4hrf
Ng2nR7xSHoUlxE3edXdwISyA5o4yI8+98uwcKYkmiQumcaroIH0efVBOc2hTzSeHUQc8+jSNIOxp
1RDHZUCiTU5Rsv8TTJU96uagDo7gqsIKzThIZ6fW0j6kj3CXqpPTRsUV2O4k6MVxp0AhgF3vxWhj
VbnuHXwTnO4zkFuiEDvGGT3NBensVHLQ6/8eURKXffidxb0YswPGsAkvhEMk0FApkTNGmUK57ZHG
RmmvavryNK+p5j4hHB2fhmJXzFBmYZeoqrhH+2CHpomTEXgO1NgIbgqiHBlfVXT8d8UXykeXwI3m
ZCZcqhaQHklMNoBhoTjmrrZ9i2ZPvJOIE5KPyWMnc5Z/+eito3HoIXRR0h6YUg/vcKn2dSt3Wqsb
XPb3XpQIlNWrHkwlYqycBnfBJjW7zm0aui2Wk99xZ9z4kOdJ9r1Al69Krtv203kKfRER1FeS9uxb
QvThRIvvL+DDNkrWhyawuE4D85jPgyKGJs7aqGsZcLUeMW+6zmfbDBlnxKNfz0m0RgwG4HLOEBT9
dTwsTQGs/cNNlYcyJOBc9Fbmo+eIIOsv6A5/2rdRxUEM+ZxTywQTNkvE8V3vWA+uH0tTIo9uYE0k
j1/J0XcVOZ+ZT1bcg8nKE9Sxxl0kCMukIqKJ+X/SweLoPgUbhTQbV4MYSM8wGoxQaHNCifrLvylg
JD1fkSw+7ulkRjqyHvFWDVRrY0TG4kyCcw60wxJyDbrsHhkwpT5+QKqv5GGGcmv6IWMyhtWUizsP
lk3fO8HpKHkjLHkqsQd/hWds9YQEd5t06AQKHbR5ZkYqcloPzaz42UbQT4C+RW154OLdv8r7HBoS
6fMRiWauK/7SK5DgiDrKCcIfFNKxbojj0ceRIany2k1hd05sjzlLldcv0x7YvCXppBpMVSVpx++o
YktL0pQms0F9K/O86XuMWogL461WF3nVE4u+oYekT+bXqm4z4azZQAEE/GJhz+jkhfEX6U3VNBPy
ziVa1AXzymOLCqqD5l2BgI2E2wAdVKhr0uJPItG2D0CNJKy3FfVbl5lYl14tEEaEt7ZxdF9W2Zm1
RZ7NXbs8UTsag+ZwsHIHO6kzp7751fjTJWOWftY53rTEt83C5ZtnsOz34a8rZKJPUjI7SGcm2AhS
9hcBNFne9yYCM7YSgmRAI+lA4LoHE8COKot0H7TQvpibKnDTUZ7rJdZgyM8D7xwYZJqQf9KrcFoj
VwQJTTZ158vJ3yMyptEDwzH6WjRrOHjC0cU+HWMqqF3Xyx2RB1JxQhuPsn2ao80o3mJt0AJ/F6DJ
boDlh3tFLq3K/zkMinjldUPU2v+bpZk/XcGz+tdQn1sbyuPhP30bVEte4OLV4s9J68y6m6aonp1+
/iMFXsxhOBE/hal6MUdd+LssJDF+XmgmlJ9dIySNjlb3jg8ZlkYXsyG2f01+zSuiYZoKCubZahBW
UP0ADT7tKzP+XuzvfoWPfN5X0Gg+EbJZmQbp8vJMy7VkhFZIjoRUMGf/Jf5r4nsSWLxi8gnC5KmH
U2OfT9ylqD4cO9XXkRTxFpqvEHv4Bleu6Vy1MqjghgJaQshsz05ouYHOTiKVhE7+WPzM4dpS1Fdx
SaPBBqzASawAGYg4XG6QjUEROjlHO7pLeXiwe/xJsSrOKYjPYUY73xHQbR3WjWikAo+Gl6pOtmhg
nmCWRLDpPaJieeXBL+kTUHLPNjB4reXpNAixP56GrPsojTkIshHMTeHakR/Q09Vq0J5/xtOgV2Sx
DXtLGyPq6w7kDTKQBgTm6gI+fgoqTBInWCO3sZ916BAyW8mPpGjNwGnh4xNdblZ3HsXTQWXoBNyi
Y87LPbPN8GNa2ux8r6e1dfaphAEe21m6mebqR7ytxLbyb/cTnWEofpcZDzXfxx0R11NISysO3uVm
g5WB3E71+1jBBZREErwL3eqLYGX3gItXShj/AZSl/ozdxUQ5ccELrabbsiQ/L5u1gsjvqHF92Uia
48rL3E2253CxY6ckvbDSl8jzli5rBp6A88vdkJvGgfKrBMbuHLtfeMGEFAIMojLn0hfy2ffi6/3N
h4qqDl70H5v2B/l8cEIKZYzomEIsRriCu1ik46jW8Id+jGd00kLJM3fSpbjU5uXOWrD9ZvlO6D5h
pU3IoR242sqUDqsUKD03GDiKfFqZbSGfxB/k5UupnAF04jgzp7SpNX3VPMqKg8oRMNeJvnN4XMNS
sZcL7aRgoJVkjGd5VTxl+JpxwCjnBogjD+ms1M8thMIFWBDOtdXOdAGNH2bHsalxuJLysYmwiFOY
AItp6Z2yyL97n3k72lpTJPULHTPxKlf4O2INCDWLrkZIhL+2g8iRl0i0TXvBGWypbrVc/3yfl6A7
NKTM2fdrNhDilfMb28sQoNIkB4UTvmor4+/pBSc1YUOMMiwQUqNWGIFTx1eJF70baxTBBcCiwS/j
yL5Deor/DyCI0hWY5jPSYKH6IlQG1Wo4lzJm6PoksCtbgv37au815nC4ybf0TcOu1DQwHApEEzsp
hKWB00yhN4bNA29XYFIg42vZQE/IFuTr/9nb1Tl2k9N7wApO9EKZUSIKLG4kZRTCKBlr/ReCKvhz
Tf0JpaAN43MAAYqfhXvcDqyM2ZHIUz0mouojmEwt24OEVJYDTusF9YRbQqyUx+NtiI/lnzkJZvQS
W6kgBg+WK/8VLBdYJD9ufW5/5mhSqe4U9TgKw88qICX4q7/Ic0kOHg4aalPzccHTdIUlx2NZYuaB
f5vzUjsnNeGoQi3SuGJOXJ7ztjbwIv6qfnlgnWNKM6VNxVGDlNfjWz5AughcEUhFkTh/N5GuFWgQ
VWqSvd4RMP6B4KHFLHY2sKm7BYmWDmStrA5jU+pyBtzUS/NITwUBCkw4iEYgWDTZyh1sk0pFap3/
hIVsO0+Jy5CwZOt2j5z9w6MOYNQlyFFlatjSssxaz5YVUEzOWvjcCWxx248Req/M2IWT47mx6bBw
SM+Z+E0KILjQRn7Rx30NWicD9hu5gLkphK0WEysQLUu2xSohyB/G4V9/T3Aze1IE6wap8De499LC
k4bD8dtC/nElAaDYYZc0C3TInygCQWTne9nGSL2k4DBbqYzWPKBGg95xXdB9aPTbSYX7qyGCiYHV
GaG17GNKKJhD8NLLMTsxkSLvCCo1FMixq1Qyyap38mucrVf03QGou4B8WIL7SdE+P5mMSpxwTvKt
4xyWhkiLtQePQ6GpMLeLXxZM+mlH+j/B+8PPc9Be9Dx+jaGdx1KcwAbD4Bzx61H/EhpbXePdSS6F
xyx3EhVxmDvKz6boVWm4liLybC1UyJ8uz9F4euewI9glAXNOxl5etend7EOsC+DPgGhTTXB9n1C5
k8YMxTtrDtj9knOIfYnFNuysbMR4WUrzuHSbQz4Ezva73piWXXmfqrZqsD+93ZdpTK2aBYaPaiFx
ivt+ldSnz5JthCmpIPhWjT9Sbc+A/5GWMuBuDmyxumiUGaMbhpgVQn1P4UOyDnkcShZHfjWixbQX
EVY0/bCHrDPfjrhU2kgpjQxMW+cQLDDoYyU7NogU73bgwVtQkVXzq7m4nstTu0wW1v05OZihaQL8
rSPXjddOfQIS3QtNblJgsmUFpwPgh/B8A6w9GPjg31oPJJ/JWOBU8c0qNEJa0yrEJ1QtXDQk6dUx
8nM+ozyKbWLWxoFNDDSi7eBa+uFWbYn8ixEt0UlU37Nu+jCPeqBCpYGmfak/9i0dkyrdNXP7lAmz
LIguRNtIa4qX+9fehY9Yii4SH9fHd0jgSoMYdo3lHEeXFr5zHzDX9UPkWBbossjmnPI11CMqcSh6
oem0RR3lWlm9SvUsuyDynCFRULIsDQNMKC8K9oVcmMGcdZOUaYdczazioZ9nRg11BS2OeVPt01ZX
75egebvxLQk3YeG98iDF89yKOkOzNgCpMLg64feeMFdgO+WdG7fkMv76ARgSTtOcL4maGMcuRnvf
ajO1SGpB6bCcB85V4G0mUrHYX29Y4t/gqlWUlcU8a4epUo023arVLrTatRny995Rb2aW2OrBKPbM
eaps/Wf9zYsCBdL0812usQy5Apx6CikyqD0ZgckLTRsQC/f0eEhXBg4T41+yHBm3A6yTlh0da8CF
xJ09nWwF7j8JbWDlv72EfFdhdbXyrTY0te6l5c6kcnAoM45qpl3Ds3ZysgOy7tZhaKJ+FVYNhjDR
hjR537KhIzf/1hIt0Q+xVqe3JQyhdOA81KNsSr9dKMsay6S9kANB+rF7Rn6k+LujF+4e6pPwfkMV
eBCgm7xCeZLv3YLhKFP1nc2t4gvp4pFB/7ZRlleyK4Jg41oAwvHmmH973RX9XVoSaat3bUb6Drn9
tAvYd3GUOhLu6GLIETy7ZL4wieNPvDiLfWQucefLnMyjVK7F7AVD5xXAfVZJFS5N0rMnyU9qCHRN
Qf0V4l+PFk9XdgTabSt+l7lCzdZ7d794mBjY63kuyzlR/24ICannYu0ymJjWROtAh7R3BQtE1EBo
0Flfmg5qV1n8SjBCYY8GQ1a6madpfa6tSOLNh36es6t3XuXVB4++lexNlgt5mVASADHjlDtclG2b
E2Iawbuq6ludcRDCo27a85MPUCU9MNaGneVZz6/jx+TNF5v7zlNtUvm/H1qSbJx+hV7JpKibaQ+i
1uNUVAoVO4oab8FZq5hsib1dpLPzUn7Z660X4DKiVokzLw6xAGhw9ILH6gRZHEmSYXFcZjrYEDoj
PCarVNVWhVa438tC7S82+Eb0a6oi6w1zLguyFkhVTy/QayAc6j0jEMPSeGFJ71cKcoVKnpyqhCbD
KrTnNRHV2wffceE03aA/FkGRC99BdMjLZ8Wnru9lcnG+XubbdcWbkytOHModazlKmm9+aT8gxaIi
R8NUENoVvWZJvFesKY8DeTld/ayszvaSqiWTztzmqZ9/VEhbdsCF2uXA0tWyOclTLpAjluIR9azL
tVLEo6JEd29fXfDMAmSE6gYvFK9r2QEWI5MozK6OTWiVOFYSWhBxDDUMi5N/DD97TQwKNQDCsBRB
RnuXtLby0NbSQct7csbQgytmtzg0Bpm/f3ZO9jRp3K+isoM5OlNJz6E0bC4ULQqhOX5B+cpqRrIr
wN52432EE2xgF0n2RflY/22kC6DhAtrpG2zLXhf4xx5UhWyYyHeXkRloxhtiQP/Hl5JjouLkKj0s
8wU5koVoQDinilWQESm32ctTR0tZCLMIu1XKAtInuLyWyve3oVPieEdg4gS8PHz17+C4TxmsA0WE
hctNmIkDcT4Fe6yU6eeHLPYTTTnzfl+RvtzOxWIYqYOsP3biWXFfInm6We8DIRI2fz7T9jQV+9zU
gulpJtx0hsz4qw85NJRV03vRTaFhXFtQOSJM7TSBOiI7K+0pLK8xBufqCp9iUt3H1QD1lxjon7OS
SKTh0KfUqui5R0eroRX7Hbz1Tq9OCBfGrhDHJTZ1Z5eydS5f4KtZ4E9kLKt5LkigKp4HgyWrPjvD
ORXJu7jwFU8vKTmHDQtcGDTsEwLhAZV/qdZUtOqtxXW7ppkTxnH38h9FlPUMIFQ83PEFjN5rEA99
4KJyjkDyBaKYtBdrWpwD/+T6Jvs0yPqrkAo49BF5w8nzkLUN5Vj4VJ67W/nmir5ZPGLKFGj/mhNx
IN5VZ8CizI3g/U8qTe8+qy6vt1g3+IcpgvHGh+OkYfMS3KsM8U4ZqAb0PKrtFU0k/rBelUYGOXwZ
eBtCYo5Wvxr5vgji3wCUxfcpQsKB7Cgm2pn/Q9SyoJ35Ee0g845l0nMHB5T8wclC1WNOh5eQdcwt
5mji2MF2xzVg5ISOYH/fJt+EvlR7vL+rBtG8KphNJkal/Kuy3g8wa7cwSYSE9a+aCmXuO7YQUjWw
QYc4VcXJOrNIiv1KLZ1u7LYD0/P406x5PSircW5cPGL9vR4agVxwsKgxzD3hbqMyMvt/aWAEsVM2
YaDgEoqpw3dvhcuoL72fSIo8YPpcg9SFNlH8beKhpFDbcSLcGqAn2ILmg3ZoMehSxgo8do1FiZ4y
cFIDV044N1ZXDlHJ7Y8/9DjHBQ+Q61CEChPpFjgZE5sSZByNGU8SRcR9l31QpEfi6ZFZvqhn99Pl
xNkJJSdaIdxB/Ih9/zI3nE0ldhWxaYoqtrLjaoCP7CavXn5JmbW4umZ3ZIjKhxT6QccPac93Ubl9
K658G4EwxwLv+PQcl95gRExzWBGSRyVGfUjVp87OvmREQpAI7ascf6g66UeBpZhDOBCUKWqGDKmb
U/ZKEapMHPq8IbNyMuVIl5FCiIum48dgVxIzXWNz85FdgZ93x1WVl0Gz6iqoKi2dvglcrJDDBWj5
JgKdsYa4jWyNs0zWHeOOxEB9EGBliukcIyW4RqeaKBW9LnPT/0UuG2wYiunEfWvW0fBZtGwll0pw
v7NN2WqqrnF4a0Ma76ifvN5EP4VVyqIvCDckGMsH8IpPfYBb3V9ts8Fanc8YcoW4hDSOiI27A5l6
CyWAMyqsVpODPnaFqeb4XAS9WBq6XBCnmAbX59OwPAJESFRwKpyLBC6mmyFAyXNXgTmQ52H1qw5n
rED/bLrXTcYl89rfY2YWtO4+YJmpM1xEK7/aiqBO2yJH4WArIcxZqOhBlVS/0ikBj+g9b8x//xBI
/ZaC2EIAH/n4na31ULQ+9a9bywYbNbzYGAv3VEt5Zc1suScUMWkPcoEV452NPzZdGXQBzCokcA5c
XP3L0/2tHNED2vFBErL7iz6XlVWrbB4E/Dujbx9HAamXX7A7owIgRnM1P5zB5eUl7W7oBnAN7t7G
Y8gF6ae5q5aHi7A0jHIun+JLXufmrHo9uOK4I2CDcb6oMYYeYd/RWA1C3qdXNd9M0q+DZpotiFeq
UjY+7MIUqwd6t0b/bPd+GzWSvxLuyG+KPHZYG8SxGVq37w9Ap1lyXgW27X0VFbN4eT2F9izDLi2W
p0g43KYd61TfOVUq1eMf904X7Mep5kW2N+n28htXxiXFuhE4d3Y6NUmNVCfxATUEyhV8YFrx7UGa
uFLjbkQtCdS4Ib1fOgrrJbpoWqpUp+GmC++/+XpaG1XUhpqZw2iY7NtiruvjtnLtkqsdBQYwaeVh
oCJ9GBBBOQ3lhSjPCZGtyd6BSTxRpmCapkRyvs4AwRD0rLe8vMJ7OfFypKrAPFJOtXMrHi9nbfZ6
uxzKaGTPJ+s9lTL5W7gIeALAmP/7BRQ+R3K13j5EOsU5/a3ECaZJo3663Fnx8VgqwYkA+96RCv48
bbH6UU2SxYrzpoKrciHaNU2A6xIuifsWm2YAu8hAdPmEiRe8syaFyd1qr5wRsh59G/rmBvYvTTUu
0FX46L3uxaxp3abHN+rX6BVSJ8u5ShUVz77l0nXIpflerBLcxBV5/VP0hIAdZzHizq72bPqfz0wN
D9nas+sN9V7mcIProd9nsvm3BZ7WPMjOhzMlReEeYBE/T3Gr2wdb1w8Dqm3dVeMccEsOx0fWxxP+
NV8be9eQ+KbfL1A4BTvVjC3E0o35WADY6Ryhc/NarkHdSNLco4NZWJQnqk/ndv9ZyOKedjzZSFq/
Tf1KUOg9ossQb4q2uqETwiXUemF+FKHR/1hqMhJSk8G6r7FCcW4IkaR+qHLqXfCB2X2oP8Q3S/bR
56beTh3TnmHnJh4VZxVEG5CaWTC+oBg3llCEkLNaka/yCzDKXqQ0QZ8z9I+LxNxwTCTj35cvweRZ
ZSLnYT7zzlh3KEQ4SHblr3mpeXumsbFQXvYnoDSLdFIZo9kypFkNOY99+SoepcES4hj/2bFlqB5s
M36lbMD5aJnEam67lXSfaAOnqJQaWH257jnBY8u+4/O/CWraOsfWRkzwFy+bGSc9Nb7ZW0Kqbfw2
UXCFiofCaZ6ZJ80sNnX0zEg1pa7+N09eIKU6XGsiQvtnoKYvAXnDHo7//BZWN574WCHWyA1+5qY1
5NDhK4KDct5b4TAZZJbw5HaBKR70al+i6HtqHspDfFn3hw8jHptpvB3uYgwfiaS+yordWtBbe7vl
p6smZVpZXN253z0KatKjhkFK3gUOyD3l5vmqWCtlbB23VkttWmWT0mDaQOQd0KvmAhp2oSMcEAC2
XzSpX0ERAFI3aN6dVae9tlps0TC2npfPax+GM3qHOe/9DW2d9YSc94XMseWp7xznLdyK1JMKy8yC
kGD08FXCCHXTsDN6lxPqX3jwQ3C7LjWvzRRODM1RBLxYR70sZLprw263nW1TN8jnbFy2DRmSmkTy
lk64pGSRcZHTTZgQF4xh5J6GDb9WBzyukqgliHZZWTZbKQYgw7aTm7SqnrJQCuL7u/8h98VtPScG
sMRBRB8+wRKkHMuGfO79zOEq5A9rAhszycMT0x2coWft60EeszN2v3+mAV4T8riUUnEfOIgLB/dm
AYAIfdlXkKTr7aHci6RJ1EhFwraDoxNnEuOxPYggg8keLzQsg758j3xCGHpWiQG1haduGhspdfs6
0PnFEIlawBP5BQSCmnbmR8H8Vv/3WaixJfUDI6Y7SIn2CfFV8ris+l7M24HCINo1IkNZ8x6h1hu+
XYDTIpqxpct0BXqqDfl006KSX4kRHkt+agjT5ehneuVoUPSotlOQfJ7gzXVNZsGk+X0t4cUtzPcc
l5mFl/qWQMryyTUqp07ltzlO8E8nAAxHZbrIPvzlIJup3mHjQVc1MP+VOQFtZjf9kchXI5fKtT6D
cBwdSoSX4GqrMlPmCFSdb+DNOAoYKIm5c+Ur5h6pXsuCISx8pgIOu6P60zBsTY8izKGPwJc28T6n
EeTIntCCfPzPm3haF2/gv8t8SJWTSoPnMGifWtqZWURUNupo1Z1M14Wd9pbOrgvjuYUOs75GY4kT
vO7x9Z4aao1RDSmIzEgNny7rVe6bS5pQcPxI6SC97WndggunuZzqGEMTbLrVPeKSJoDpNvotu37n
rtYbzApctoIgd4liaOBVlAgsfH6E007AxBaq0kIS3JII9Cr+K9PnxBm7ASRSYZmfSFwW1INQbkCj
8ke1M8diO16v2LO5rjj0Nq8wvoAwg6b/VIxiNTfu9PqnVAPtfdtjQyWHbct7Mp6LyBT6uor28oCw
3PMudMIaPo31cGoPjmLJzZUeBxMVklq7PDPQVrv+chYmXvRU7+AMRJYuLhHwesMfxDfAJkT0Dj6e
AiNuE6laXR9h0wIaWbJvJrrf+4TwPhqyD3gUGYCwyNAdkWMpfx7WLTLsjYqaWXMlkXSii4s0EqMK
iGZMC0oOaea10EHe4QsxmKA8m2KDpJCATuypufrlY2r7zGtMKur413xr1ey8RBbtzcWxcmOVddyV
mTEXM32tF2vTjeqy+9rtngbuzPipHOQXVUH8mw19XF22aY1Hs1khF1rWCRcp3gjOsvxMfM+K5C5M
zlRXC1VmM5+B2R2TvgrJUmL1PFUWknI6JDGnDn+e6ww9AyBBHA9uSBfAigEDilJXcW1bXQHbbECz
/wUDlMqWXn/YqLp68u2UkmFq2AFt0GWXEGiWkjKSmDYvSpw3qnBbPlW/v4ZxmlzoRHqUWFXmFy4E
GgWQ0EuHjaBF19joU6NXx72goGRTTbzt+foqlP6LTyR/twqOcJU5U4Fd+oZpc9ae7UxOqIFpz8uj
Fmn5/ats1lKEgCL+UqXW8KRJAZOQ0e0Ztmo7u/hEuq4yVWUalfLRf6PAxeF15HuT7jaQ8i6ySvYV
Zv1SslajGaObnwMpzJ3FAu7FqHOwe9Q+O8ocUxCjIb5YvUxi7hFFoefumyrtrpuYBjLqBItQ8w8l
oXyIk0hl0nsWDKYZ4vz/iCaomfyy8mGxo+eUCuEJOE0s2PTXh1KZK3Xs+LGFbrHQqNQS/N6hQ+8l
uDlugYshRKQJnKfN44uMsLRZ0WhprklTzqfRxR8OYcxra3CV1rko5tW+MOF+jNVQuJGZuXGr3fG9
V0fIbdQXNUSMEuOGIoBS3Gh2TmvMs/XGWuBEglKnxjeRXMx5MdD5ofgfcVTKl0VwfFGcpvkZGous
YfpSfYZ/FVgk31gv42oY9dGfMc6xvwsDY95Mrdhu/AU8cx4gCkJXdIfD7g57X/hA9mhKus8IVnRi
ixls5AxNnbd+VpNJiXRPL9EDqKZNUXHBGBQXhkfd8Y6hXaUdseikUYLNHSoLJKxRAjSWBu0ZV/IV
kIshtXMdHGUwtbyhkeSmBbFQKJeB5rpCQ14xNLWsN9Sk0BV8YM76v+bME2koBxEZIXjhH8RVbgDZ
k5serRVXqaeta3qKMABcYLk6ZKGFMc6xl3rf/ne1wy4FdfKJqwibfLHx4pRwtVzVRBLnHVFCHLel
e+j9Ss0whUdirMj3IpLgJHpGDBQ9l/57BKWR1mIIZQaLiV7WmByaFpBntFrDM7PgxHXqz8ylEiV9
SWnOfTmI+QrJb+xke8bTDwpxVgvWCBMx5F4JgMAU19AqgwRsuya44hm835gnzF/qutRNH9qPq6gO
wwOZP2RKzXnsACagjgyHWuLJ9Crcz38dFgwyye/eYoTAkRl6UwEVBcgI6Jk/rR2q4g9EJtmtsJyX
h+VixDNp0A3Bf0mKNoWX4MnyPw4dVBpUXEEB16lWdD01nxHg5sqvEx8jgSs24Z+FSG0gwnFT/qax
xYYFPowUyy7D6RDHucXSdDDsytCdqQoIPQnSIg7IsjcGSR+Vm0abCgz2F18HykCLhriyzPtogYLU
R5a81fSWDf+E3/cv/oObMNrginSy/rzkNtnVMwg+dC498OFQ5WIV5sFmyJb6B69xLs986Z3lvi4j
mIAI4ZbFt9ZM3lCuLludOx8LaZLkqKcVHPRat5AdM4AmGrx/Z3L3Snu26QNnkDgyRLwnYYz+YseB
rVugBE+rmILI07eckG+lj0cl1IjLKe9C6FBYffFXO54I3j/W9xjtpqdRfDDWeabn6sPAmlouE7nk
HfuU6XMWDyE+FNtpdhEL7EEgioWvSa7/NfYjN+2wqcsf+xyq3RHXKpP0joRd0wi4V8L2txfA5yAD
pS7lmeRQXwHt6oy6UMm4ixm60Y2h4pl7K9MXFmaHtktDGt+M3hxcjh4PciLVUWMgSG0tr8CHrZPa
Hwm0ATxfg6y4cPeht+Bd8pMQFzHnC2nNg7LSEw4bBfYx3P7CRf0x1GjCZadjuRlKDZ+T/DSFEM3H
SlFHcxitsV8BmMyhNfFiIkkraTprTErbEr/FVszFx1K4xZoxIFy8ROKg1J16uLT75YpvxvTD8Y19
fIXdnvNgGZi/LqPh4Yk/TuW1XJbScAAY2NCDH3tfAgz21/S7Ke0RITbLiS2NreSwRVKUxZMfM5W5
v53VA8KEfvUu9czZ0WoeczW8QyMFtI7x0vQSZJJaQU9QNKeaXX4RjvbVNXjWePJZJ16HoRT8SaCv
1vLnEJw2EWeLgWgvFNc4zTfBT8kfXc8YftP8ErBBYZ9ig8cGf+xn0RBMlwWJZib+3aRiYfU0wh9l
ysYMGqJKW8E6/0W49zgrZzlvJSXy8BRX0VpVTtaJrPhjls6KxOZ/2fKRz24RYHkFzI8a26b6ar/5
0LX1W0e4WJZL9Sy91IsEVNkcLU5L3a1SYIeyJdD4jJdp0b4uvo7rbORRggW7djyKHR+9RIue6jzV
8d1kpjAxWEFAO8O/wDclgOJU4KxZehwz48PQGWa+yFi+m2ydUivR6gxIDAVlzFUE1ISDYsUsAsjh
7LDjAZ+bSUdFwKaoAHdYWz9fPzy6a/5XxopN1t57EjY1t6mttB+3oKSosXNOfrHGVc8CHMaxmQyL
xQKy5Toxc1mBzD0kNqGf8vWGIx6HXQxvS+QA0HmXNzT9RrXO+JCYltU+VBMjnnC1oEtJDuS+VtGe
j3gJOsqEMJSeCulD6bvpYcOORXpCmEtTLZ88/kOBJUXc7xbONuV+TAOhI/hOsiBix4cys8fSOlVI
d1y25555Ow9HGv4/QdIIBpxr/9vkxEsdZxBpq6l+WwlIVLpB4BrbJHroSeRsjGeto1x+dh4lc9fH
pAPcodftNGWbPW2WnSrP0oWDkiRGliPM8MmOuZ/v9O5zSpsw3fxjIlS/8t6PbkNk15tblhaJM892
W3cvXRY6nVHNnor4PWcRSXw2qfXbm0sWzsCggB+0evc35CSdoyMEXqw6sC5MFodWXUXGAXTX7f4r
Z607JTxDgoOZbj/AC0tCFlopMuzuJE5pb+pY44fIzBVm/RzyVA7b5FAV1X0nnHUkcj/7vExMrNmh
49wLF6E32JTunH1cXFnx9EE8n0f9VNqGTkaE7MdF4Gk/bnKOynVLDhmyfrafAr6JTNwRFhoYJghO
ehol4VKu535hK+tcSIQXRFBQS8Qg4srll50GsxthHoqEBbQ3Udc1k6ewsIQflY8cjgfD6+6MARHV
LaXcKk/WYg+rFwSp0u0WKwc04HbtEM71Eqb3zoGPd5u2yhsKfIQgxKxy1/xx7n8uVTlHicyhRJFX
mTX3azar8EHAoknLC2FTiNEvmfUp7K5qtNbTXBYB0mQAocYr9aZXbvPIgmjQDUEIYR+BQpVeMhZW
BW/sMc5ywfQhncU3NgOsEY0goZiRttddpNxzOANaaBEhesy6a6GzCDbRWODNjYvXXXDkyAde0vKF
1ipVoZzgjSQgCKo26hnq3euYEkrfKXIKeLk0UN1eCN1tKx9BRTRMtEUkZFoDcm9h0fopRduisypV
ibI3torKrba94gBJB84j4fCjd4R1OmRjehzBtfASq2G/jmB/7mTiA/0O5PIvQxcJqbD+4ccNEcTF
AB82V7r1EGUcgSW26GggrVlvXnlQTurmpsJbWcfROkejXmZ7hI4MGHtLlPCudqzRIKLRQ+btrVfY
1XfcL/sXijQdAzTwP/gKK1FoCPXZaCVFREHKZ0Uaip+bTF3Ww7q/NXcRNUO235mSKcHwzRHvPnH4
yHn7hWxbsQvuOK7eU9OPWbRFEs1i/bYtHQpbaThp86u6TVDvMRZdW3p6zXcZfPZEqZcxqbBfwlbE
pvG7RKdHp/GIm7Iic7ve+F8+q3zYU4bs3S5/xmFOidDjrNVEizY+UMhjRvyfygtL0opLWCMem+Ny
ydrQLJ7dBQu8jqrWB+FoXC+6UjCjtdJARaV3oKe7Uq8q/H9KZmAh9lE2yThqcdOmBBxLeZqlfo5P
XsXEBnkuUk57WeOaathNKAcr7ST1XQ6v2whkVR76c4sqYKUhX6gkWC7HvU2KCJ3JrvI/b/57SNUf
flwRKfA3mU88zit+ZYIxmyQ/9292AGfsmy0KRu3xXOu8/wB195M3XmaG+ZcC7GBu+aPC6EsJR5Iz
eNGCbXSucO1dF38+FIMn1aQaJpMyoKhLY6MR7quWxLo8q3EhbK9Ppmh1ef5+u2WehTBtHgrKYA2h
rJne9RriPhVlpzqMAecGhKhdsE5Yd25YS4KJIK4Q/JhYNSOcQUP9ZivNh85lmMBKEZ/pM00q4mKd
3YUrwlLgQQ2JabQbFkl0zUHGAEYEyAnyola4+wzW2614/Gw6Rf7cYuK27iMtlBxMi+700RvcWwL9
ZlQPoq0ToFOchvwzxQema9Gumg7aTN2kwsMWNIRxXV9n7UemwRhKLcY6X69EqApEZ+uSpcFXUEO1
b43lrx7aQP44ddOwgtvr5lzp2eXxxS40JqrrKeLF83TnDe2xKtdwWXlYCcNZ+XK9OhjGwTTthUbY
oT9er/NZbcafRwIlzKlvJfO4SuRhDoYvXRzWVhvimT5sgQXmq4TD+hDsz2aoZfYrcSOUytIags4G
RGTsyqiO+8M/h55k+8tZ13dzpBYSlGbRvrK1vcEnXMxy3Jq2xL9VtydM5ZHU5vT3VRY0mh1ql+q4
s9AbfL8oryCxoO0N9v8kHFIvQMGfJEvhC5WZzkVG9E6UMeAfcZGvKY5hlruGMgWljIDmDA3hSFnK
M9DDHzEdAVO0UAGRo6pXtCaXJ7Y9XKvjghMzbrZI99+3iqqNU+8BXglc1m+y2LC7VO1AT6kgajSh
ZG68UiU2TikmooRbinxyWS0E+9GQTxMeS2sEN+UCU1ahjIx1qEzSJhjgtXdeGxUMu3Q9OUtl3zXd
4Ro70Wy3vLecY80svTmBRZBUfUKxEUmce63C5BmtAwHCik3S3DA4YEt29tFqeShlBZL784ERAUie
qE/MJPNT7K5I7A9awUpriVCdh3Yt7HC2S5iVE+gLBK6oWp8qE/LtgWVeCsLARTMmq+qdKcCWLcMj
QuCCxqqIausJxj6Bb4fFeeHsj+tOJFhkqf/YfzgtFbgCD8Zn84znjW0Oz4NX5VT9Sxafvkayda7Y
P+Qqs1M9ehSjW0cIw10hJzMuTxS602J7jhwTrgNmKXnhoH7maXXtXcZvsHEO8luRId3Q59qbF6m/
kulhmt1uPxqBDw/ZDu1ZGT4vcykJEs43XkkfOnJLiHheKeq7NqK3abBtS9FiK3TdsSsGsP2IXV8Q
s6/5aWR0rwMVbggKDSkCxijJ6ost3XZJyLVA2N6gtknSAYi+3B5ZBpQ+riydrRYeKc/WxlERygWk
t5QD9Jxe5d6ueWqcOcjsqVpqkH2LfNqdZ2jijuWBP/Wh91f4mJgN1vh1zWW2WRpOKN1I0GJzo8R2
M+oXhS8L3JPgnuhpr3MmmNjupH9if+p3Zi7qx12q2VOQCQr8eTAA2W+kRi7JCkDXAL2CSNQfLnoH
oWpuooMeOq8L1EyfVF3Ndeilfj2IU1srRAfWfHpxj7Id5BR2vBxCnm3tPTF9s6fE0gA6+QMsxvj0
blIRq/OJMyDpHPA4/IpYcXnBIMB9JuiiMWC08CIBZY4mq0b6M2vNr3imVrE2+Qnpnu9x0vhNqvYl
4wD7owSVRUyt3TpM33VGrgff+8qNyXbqST1MOgrN+ZZ9w05/K3BZBdAWwu0fhvyxnQgal31R1pLb
yEgbM9oBVorHEoiOvuP9BYdo3+qKQ7zBp47Qwn0oma3mST6J6Ja3/7Eh82YKOPIBd0PdmM2I5aFM
SujGJAv0umqnYylF3W3q+3a8y0EHwOeLdrpLEdpTd1Q3BpwjqM5eb/JDldSbc4nin5fbH8WB/y9O
Q4ArKDz+xwGcBRuGNWUJW8zYAV4Iddqx6FZd+EZqnoBI/YESWyrbRg919f81UQkFf/iOTeI7hCfP
aPb2hAOOYEn1+jUZAZCh0CDzkmnlWBcp0fkXoHBfmk48By9Iqyzpm6z23OYGDW9M+S2FGEXU1dX3
DXIoXYOaDf+NZ4KmtKPOQoKUI7JRlkkXddWxXEyVQaes3E9fhJw3ylzzbqGcTxfVM4o4xhilmgY5
U1cB7buk/jn11Geqtu1XhPK60ghVGQD4wSA4ailwXD2QWFdNqAv0nVnb/gO11skciaA9TcPDwX4U
wiw31BBNuttAk1t+OxIAm1RvxnVlfGC++M6qZGx7WkRnlVf62BkDGiQ2JiXD60VujqhNAEae8kj2
Tr+hT0HQZkkvNMQVHU0tQ4jGZicSoPGm0fODTvzmn3XdCbFAnjkX+RJTX4L3uaHncnhNh06V7uMd
+GqmDq06SrZjZgwUudNpuVgGtqmXZ2NBEwpQ38TZMPLW9UF83vRfoS/UTQfzTKrTz6wzvBJlKN6q
TozH/r7sv6Cq0oYbdhVVWuUbzR5R5L/PUNT14uWzkrf/6ETFPFyehoklFTdl8qOetKMuAegJ9ufI
a4dNfsjwhshp6BPZ5upRID2WLl7BZLwFDl809CG1yp1q09CcQHxfzYI5KPIFztQ0xYTror5Amdb0
j/mhzmOvHsUbhqurSDsJs70zDWjLbDtc5LV4RoVryyezHmXWi6JL6mhqJMrywalKXDJgtBOLWzl9
z30rUJSrH2rUIq4aIuf+lhkZF9Z4j0vakJDOhsr5SQNiZhRJsMMrgDeH3yTcsQAVOMT3EShtNhFN
Lb5kxXaNl/8379sKyyxhCgB8flm1R/uqcP+8ke37GmWGDn55ux3LAvkLThOwlt6lu4O5SO4PxcUQ
hEQOQFNhF8DyoKUDRu372pAef1eTsltUyJAXKBPVFVqIE0ibzpI8cvNziTn/GEJxDiJMhK2qoHRb
WVCVQ3FexseLtm7u/kzNrAaeRi+HU4lrN2/b3DoLCV3FTHdGgWKBzxqT91+7+/epbL6o1Vv9Fc5W
0udA3EzuLLwqxwKlrxScONKdDjhP3wLvu/UI9sx0xKQ/sgbS7pUa4ds3WlR5BorKh0cqnl+5s6n/
+greI6DFY+L8BO38oevjqJgkBt/mxq0jBL/o8AB/HvfFpEc6dBbEZgZzmgKfv1soOUraXBjliM7v
rjPQatiYazBc4tynbjVlpHGl7Ip4xNkkBTjDWDuXnNdYyPWoa3XAhDEqUsc6c7lWSVfMsQ9ZUz5A
7KMikOURHg1GzyEEuRBHWI4dI0PwMuE1mKR81Qwriw5p/eHj6oOyJzs8nVR5mHZDiAe97+fB2UDW
aQJPQDvRbuMAAXgneOET0qXjK3kHY/QATpLJSA38COnbtUx7FEiowZ4hg5/H7BBMj4tfxJBjs3pG
cHt+MTENy21PctYohKKaokNf4hM0N4GcKI0h5bfUuUowNZ2dX7cHUij4fAOlb0QSn5iG4vmSIUlk
Ya6brDdsYhtC+txstUWS67Q4JVKepFlk7Sh6fF/lD3ukGWf0EgBXORhco6mGH8j7JH9mvJe+PEgM
oWYGkz5LZ1CZfi1vfpb/ddWhPuENx1mFAjqRiy39i7Njcz6ve8e2NpSwubQT0M8YojIXOwBUlKUw
2X3N8NSqrKaPx0WCFYtW1XiuY1SlZ4zaZDW+3x6H7D94ZMcY/K9QZyoD7OGRmz2BFKW44b5G3Wtp
cdtBbu/uHuGb0Zz5+bmG6i6nEv/B7XtyG3Y0aQqzCaG6ap1/fy81fbPglovv+W3tB5M4zMZzSK2w
6Z+LBIVd8FvbH7nr4dAs1N1UyF+y4if9irskEphgc278f6jQr/YrNNPUGvudQOU2i2wD1MqMsLbY
WlhycpjcZk+NQbnOakyUOwJPYIAB4ysEyqVglsPZCrK4maCnr6Rlv/tqSlv29ikJdeiNRiF4rhVb
ZQ0rqmDwKtP9ZKhywNHVegxaozEvsxe8lWUiyJXD02DwHxDXkTHhJOm2PJw2Qvm2LFDGeWbfG1P9
syk1leIo25ajH3B30T8p6v1bcXTlVVt20DZdbM7kv5mIh3ORUKPaqYSb5+v49BinTYfQarEuo0LI
z6E7mR7f6RIx+JYS5Mrwz+7ZfmE/FLmfATcF3Hy8HsZuIXKbIjO3O3AcEmkI/jCDoI7lfaG23yZT
61zobv2AfYBOiG7713dcKu+b6CxAluCBuLyQeyfWyOqRaea/l022cEvswP5RhncntwL1s+KruOr9
cLAiF2ulX3sXug7UchOtvNjJs4cMNaI7Tu6AveWNV3ao36wiiwMIdEjeJ+BuWswSHUGTmuBtzkvj
hOrYVxx7wcirkesDr0uOVY1zkYPwE1qhF0tF9Yz9xz8yjrecrjOTL1y1t286jw7XHbWkJ8146Dni
7e+D5wmXy9+j7T4JgBQTwiWp7y7v96iv2A9w04cVNjL4Glqxz7W7vIRO3nWgrxrOqwsvCCRSxqEP
HDruJDu9P81FFHVlE8PwRwoaocu0Qma7TiGuGC67q4BS/Hq52DngAgBaTFhIt3EipqX+HtsrS6+Z
5vMkZbQhYDYC+QXvVh2q+1YYLZKuUFlbc6bcDeMuOdz68d+6cf41KWZJpmDH/tmyJcn78Te1cxYn
bvgMbDgAIcO4Ni58DL/VnkH7gwY6Vp5sCeoCLnH3556B2/FkKc3mcELcPuwhPrf8kZ1GDkqnUxDG
ELMroKo/BZpsWkBUibP3XCH1fS8RFH97QbSHkXnDQkZRCL9JxKpUDVslENywmAqH5DtYNh7nhNOv
xlRao+e0z+9fq3F/w3cKXTTZTGbJuNYk27ng1hJhIwh6gAMcTElOcNpT4pv3yo7LPLwYvB/WpXTZ
lff00b+6o4pSd/hsdX4bQkeZCnuvJe6VQL7TsVejvfcN4BAmNktfteFBn6Gl8phvv4J9xhOHzZlZ
eTJr3u7M33yP3fEIdQLd0XAsuKI3Ija/VSgwUu3iVrgFxn8S4dZsfYgZSoMf9PhN3HJF4NIeqNwT
48GcKcLHvpiigXiKQsh5PQQZ/X538apHKHwK/snMQzbYMrCOTtUDMdhIAelyyaNN5VTUw1WWtfWy
Mt9qylk546oUGG8bZhrX5t4/s3N8vVBW1CgIMZxuHkp1BoaPyNtPcFtqW4b4v3iILHg9OWDi9bsU
SpRaApKyh9g2rLe6qCYPxiTThSxzGzp0OQz8PTp5RkYKjTGSArEb6CNwh5Hs7dPBmXZwqbW3l8g4
wtga2nVWA/I+NVHa9MBMN5SUp+ovhLvQMS4D4xcxmLxgQxL+3Qw01cPJ8cJ3ddOcmPPP3jWwll46
vov/7CP74C/0kN5hgqetsDp5BNPGDJqQs+G5opJ42c5E3Oe7RSGlBBvx3vUXpCv3RA3VRRAANsBy
yK1HkMwuLp8P1iEy0jMFqIO9fzRCTsBUDj797WmFVH6Q8l0UWe4AmlfagH8O8ETxdtflGzfPpJai
ZrlSDLIo2ayqeeGihtbIm+zFsBKG9gARswK5PeDHWfzVKkli2hpkish1Lx2BEo+RiIqB648B1whw
rJ0HcZTcfpWdKUAL0viYX/HK7k/KBI1vlyreCyLBWIX9k8g96IZhGuLf4vrxnjkR1iaJw4Hqy7kW
qut33Yq87BI6ZPBZbrHkkVYAL8Ce3U/dmBBTvImvBfBgI/YGvjmBVEj0r1I6wUofyoqGbuF1Foy5
laoblZqUnGjCKogBQeyYYYxGsc2YZg97FYhjz2qUw/cIdmmgd1in0xxHvsTZkyQMYZGGXI3bv7yD
zGE9qgHJAtw0OKdQ5vSVrdqzMFRd5BWCjWePBlIhKJlLwzGXbCLYXZk4bZNz5xlNlf2LeKtWfI4u
qr0v28h29XUoT3wdYEGxf4h3Rfs6oymt9pUk4DTozwUbpN/NT72FzcZKswiJGkvH50J6xxe8RNR+
3/KwdT3PRC3Oln5iTRr3WmkgKQc4e2p5QTbR+POg22zZS+vEZEBzfre26iFAfgps1ORi7xDEwxFI
sV2bceNa/XxR4NuaYlCwq/6EkSl8ftI/6dt2XmT+rYHB2/XE+O7Drb+UGsaSoq32t0xOfWrFgi+o
zklKb7wknqBgKa9UmDDA+kb9luNhLX1wGQjOik1xdMy6FP8sffdsgY5iNjJqQ93PHZWKIQO65s0C
O3Mkxs0Z74ZWKpN9YB2CkwDH2s9Ourw6vZW8oLoYkG/VZ2u6EYDnF+VILi6CfxiX6YESIrtwkQAx
OrcCxBlXZKxwQWcDJCPCKK529ufWOGo+YoHyd6y5QjsldxJ9Xr5d9lt3WgWBeHbMqietXs20CpDR
IOhQVQr1/UP83IQpWafWz0c1efdFQVbJj/vPnMXRKAcsCEk9/9z7udK5wg/DsxB2XjzvTpJUEvIP
0SakOqiAjoS1NTd2kLgPZsOZ6EUzReN/SGMza4CG4Q/4SqZ+GkEAWnSNvwe6OBOfuyOImSqwbqOT
vTN8mjqjngNS7M4twpBIUlaY5XzpTOL1p0loNlmBFMkBF4yYwMnt5gVVDhDE22bDekvav/Rm+d9+
cuiUTxGF9/i5MmJ6Kga8Au7BMnzYmMpoisnHVFWuCHi2pk/1qunF58OO9s6szrluLzMxX/OnnJrY
0EdFymcJrL1y5NzfOQddeDZIfi2J0LfRnS5erU4/I7d4iwVZYWjH/9Q8cBTZz4vJWRtVsyaYhA1k
uBBH1w/s4MhEsC5kTrvR/s5fQbRt1ZcTkrs3nZbYtWkcIGpSHxoSMJd7tNpVXhrU09qRanycwjYk
zplK6amsDRgosmhawo6nvQMzy2hObDQIXgmNga3IW2WeKR8N4pAuGbIopLhPuWWvgW4bIRWf5dfL
rCgS9pcUUmhz3oW3y6kjqllyYd/9V7ezXitq+KPvouWGbXo8n79b4CR3GAqm4PcKW1W4b/55Xs/8
cEJ8N7RUaF3bQiFStTiBTL1U0qE0WOyhI0mgcVSRy66TxxTTMqcfLJL+gN6tC8H9PkyZvG70Hnnr
b8YreyoJwxrv3qc9k8mydu7vfJ8kVlACXf9F9RURTl8lpLhwD5YcSEJRHYkcOdJPsvnrZgJa4GLL
TgRGcesZYRA2536ENA7y74O4X1mxxS7JmCqggrzWADq+HGW7vn/T0bl3gM51ZWUzHXQUafBmMZ+V
1wNx77Tg+3hCRA5f8VupxGC6aL/xI7F5g9c/cdxtXmXnTnv/X0sgWFlqO234KMRCzEMyYf9ktI58
RlvFK5h2Ah6r/52xThv1U7ZJt15ZvDdM0oNtBY65wljN9Y2uf4tKyYQLT6WTTYB5QwS0iqXYQcJi
yFmFeO+660Yvug1tjoQM1gRaszbv41t8xnAVuOJ7HSc2BK58pEzY7IaWBYl3iC+zsHHmLMOVWRcE
IEsIpF7geen91XulT9yBRhhkOMMoTMre749xbDlEcQMuG8kmN9NLN9S+73RbBBFwMxaVecUJbj1b
9NSchvAxnVW0fFG/JGuFWEVjz2b/agW4f0WnGEP789TZIUr3nQRirOBUdK5JNC6f0NVMD5m5fQpt
QW4ym5P3/Ecxf43QRTRVtYQvk4i5uNxSBHV4cta60Z219l6yh8YMh9BXtV5z8eIORYhud/eMLSF1
mi2+sOPn3GOVaOQw0lF+QKRF+6IFxJBMkFD8rmsqyPLODwbmLBgGDrQE2EXEWzwkiLJl56WFON57
Tmhv//VEgQQnaS79Qo6Nq0wT3nctEbkeXQGRj6bPD54Z207T4EShYnAi1g43rYFNywr4kCQdCvGl
XlN/cDxhVZVUgxUepwBox5h3EbUIyh0MWfF2kFf2hdhe/S2BYfYiPa8M5o18vyENNbeMf0N1r5Ur
g1WdQboipqRCMyGkwEeBJn1WXsNTWR4IeaIyH4Y1SfPx+uymv0H3VGSoQu0KS0sPFUisLjDvv9Zi
376Ql2dpi1RINKy+OxSKkcW9byu5bEHmBaiQL13roGl59S3gcLbnGMINsLjCR89Ii54BFguQ811k
0EPZg24cdJ1pe2Y45de5x4FwFSD8j1ile9OODipFuDRemY6cH9edVleR8S9bzDzE7jI/xwAoFN6A
HDRf4ACQiflgcxS0b1FE9/xm/TUtYp3ePcFFTUgn7EphQzLgLM+GC2Qel9p9Q3TXOb5Quvbqz82i
+FW8LvgM1r8kUbW8TmTiBZFh/RGCtN47sorPClndlzHIWdmjenMT8KvQ7WiooWcJEZCTuqYO+Jb9
jmlt9YHKRjTCFnR00MZmaysgWMaxi0Xpd1tn//besAu6b824suFx7x7o9SlydEGG0A26Nr3lgB/I
t68t2d/1BSrwGkzYbzH29lMhNT8x0gDb8ocLRMYeyhWw0LBwF16un9TKNYtJM+SGDCEXmlOIbpQX
zSX7NQHXdaeBWJNJZ1KWK8W62WEQtALxXeYYObTKU5IT1XabbJwqHX/Lufax7S/N/xVPib8qDDgV
eoMjlLTrUTTB8zv9YV0EH/v5z04vhRaLBczPu6P9TiqB1+pRKqaDVj5qqV8FljSIEu29fGxTOzp+
Obpeo3kH8OSsxw1wewGCk/yA30n9UyWzv8qouffe+2C1wXYt8dIaEidvFnJCVph3+43HKSPDBvkP
77vXrprsUwzMk4BhoKCcl3OTXcxl1PJsLSLP1Vs0Z7VZF6HgmdxsfWFMQkLZVW7tc97zs/TUnKWM
JnaKBl5R3HB/D5CX2Y2hneg1KadPZ/dHut6YTN5J4kjhpa1bbf5IQDGuraF+na/2OfMQQruB0Q3C
nw47RfUkir/9rnhwp+pcVel5SkrufoCW1Wf9ezqTjCmzeFVpjNjHhklkJ4JVUUqmmSA2shNQJv7F
kXQzC7db6nkymuDWNn3u0qal3zU+KYIwSEChYbKPfSp8mvnYXJoVIAIY1DvOsMU1pOeaqzOpUCEO
bh3Zce3Y7Mro2iYJEDg/AcLfFG1E85zWtFWbtUOiyX5DbhoCBRh1P2PQd0xmRNDOcTR2bY6gGMWK
+vXqIwfqED8524V/AmExGiEjP5jtnJ1McWZpdI/EcsQNusUg9GNZfL4U7vpRigvbneBAn+h293ZJ
atnxuHfPxuT70Dm+wlGk/G1C5vhasDFNl5huhg8vhswljp/rdR9Q23ky3xNnyvwv0TSEiAC+CSU8
YAc2RZLlKieETGjlfkbNv2fI8m9BqMjvtxFqsHZaBlBkG3RXi+29X+NxGkdciqXVJ34g3W1n0l5F
m7PdCYhkf6VDI8FDp39vRL3iHesdgDl/ufEKul/Z0HOZllnlrCAseBihyOTTM+SAlvOdUsNeZl+B
Vc3OV7xqrcHP9ap586fQNetSULrxEightSWXiU7Qlt0IdF6QCtM5fDGcrF1e1wfUR/zHCKwbijFG
rig4EzbP0GtMta3+Pi6bAyxbhHgFbCnmOxM2otLyEAERtyPZFSgkSZeXfCyZWVYV0ZZ5RNRc2CEd
QLQnlbjCqzgxtt1dH025yY2eiQshZqc9rwwazgzjAY5lPm+SzFQ0+dj02IHi7nV6YiZGaQW6LHqL
QcUPhTOoTGhKvJL9vzJpdu/9/ZwdTOd/yELlGvcoBLRdeWf/7S8uMOUsZVRguC32tpNQk9reGbP1
qPpw/00JXzNuyoLl3ktoeQh5lFZI9tEfIYLB7fiAS1KE8L9nFi30XR4RrKzVy/lZX/2Sp3JQA/Tk
b7ugigE14qKgp7pPJsOmtwlA/W0tm1iCMfXLPcZ1YXbw64MBl5OdcnSUuPYmReRgrmrqQ0qsqhSn
gveXEKIuTwPW6p6Sq8CrlZDjdkeCMDvIXStPexxNLKS/LOIiTg04UgAAzEbhIG+jlRdoPE4gdqgj
uz0oWAa2qFbZeWmzRaQhSQgTnjSA5iaa9yxGqmnLodiust99Wb+yz0VoG8Gu+jMx9o/dsUFwh+fF
yXwN9LmI4tRpAVLRCARq+RECjikSti4JFIYybvscOtgYsgt1RO3E9EJeKuVCzksHzbcW7WQ64Z42
Gv6gqTzg2TrIdTBtEOzO6Uv7nGyo8FD7goryyLannJpnFu39N4oDHnOAKZdvArfq0oP7NEWt3qNP
qG4Z44LuzCSa1Y6XHwAC031f3NBUZLF6m8xGjpzBRLoPLPsONvki++TA5gy3XcGiGnv4wui6zcaM
UqswpvpHZbHZss9A4AeQlaurc/qtIAw7MiDmcDVKxVXKHWnbncB5ozJNdYZ0bZRaRE7yCFoZ5khu
Wd6mZe8kyj8fHD4wM4ZSPnkogLVMr85Pqqaw8w1y9wd55YYpsl0diRH7+OwdlV74QX9kVdEikqjZ
S1Zd6QYh4JREZQmX8p0r+HX4I96g5BGV+MzjG/+vWE4ncfMet7OhAcWQTxStPBP73Bpi+AezscuN
ekunP3RK0yK2IYkO7okJCA72bF5/ooezF/LaDGE66HYnG7agzEl9kYhKmeRqEFoNUif8GG1P7SJt
atn7b9DKcLneUwpIs6xs7MmhVitWOsGqEu4rO1jblam1bHc0DSYAFwSjYwOJ8o6S/F84ZnNewPr7
WdY51MlWZ5jYarskKVgkNJ8Kik9fVeosYnGtLvcrgzdUMghBq3UBBn+Rc1Z7AlkarmVsogvmH+7T
4cZ2bCRJwRgRJ7SMj+w9oGf/wGDr2vd5JYaIlGl3oaoQLxDZVY0ZBLGTnffMUma1E264t+7w5cjH
KKPw8pNw2p4ZzHV4XVdJbQBovn5PSVlf7X8ELPz49W8mXV57pQmW6zDpwIHD+H+8OvljZzCmXb9V
O6WN3WNd1bmONf43R+rJUxo5SL43MU0pEpsuEP4f5n98fQ9+I3cmr6b8DJNF+FqzyJhgAPlJ4f8H
Ddpo7QoJbvcjQu0V/yHwSNWXl2OYBJgeOie3nZShICCkGiBBRIeebHrixIictMfCG4uGfwrfUd5e
5gQsy4DD+YzMU1Z7ofut1Acsnn7hZ6fgeGiHt+ed3hutZr+UkPcUQydegt2yCp/3BuMa2T2A48oJ
OJqpi9KNe6ks9CQsLQ4wI0nMbk1DUMnp2UNKp8CSP6hYA2JQK6Z43ORP59a11eTnpFtotKYod92I
7q54s+oxWPluJB6IGFFfIEkZJnMZHkYzplJ1q7+NWGnq86z5DSbCzjzdY/GTTaVu1oJ83LmWzYKA
/FN9PRCs+Lms/sA+aeE/S/dXmo+eBo3zl0656FesBxnD5ba3uYx7gsgZ/mFleVHjIck2G+/GjhGS
uFNdl6n7GCSvrHTljwJbaFvYOArGf4dwFNh39LhsFZWF59t9r3YFSMIDclWU3xpwJN3d6K4zi9lU
nAKeiNzppYuc2aDEWPT7PGXlQ7bX4GnFpJvSUIug9vKNU2ECsK0TJGt16v8stTAqoXpJJZwF80V+
dJTrxTBPHFEndu2VXrrEmEuGKPYBbKOtYzEDH2Gr3hlKKZh0egeIsu3rLgX9rT16UO6W7qSS+N5L
E/IdFmFgk+nxfeuygI+kEXmq48OSv/ouJFOVDicgcJfPPT64xs2GVRRynSlPGvRodtWYIfJVPiVy
hTW38adrKozwayzFbyy5ssezspeFP6lND4Fmw/jhWNSJT0csQaxNCtv7yYkitufWkTP2dlNJ31dC
brTQNKoJK/mzr5/Y4bDChhyqQ3SSu6zDwiLnQEEUJwoMhWYwQr2x0rwPR9QjOrXzUsJAnzgY6xE8
mu1HMJm/nWdrYRFibEjL/csTWfxDvzBvZRbxHPm7UTskSyJpb3WET32xw5/EUWy24TCGrdrlxIzK
8vf+RYjfPrM8eYrGcRQUZssmI6wJ+ucikFpLV527vQBtYnY2Sy3psutunM1wnffBImjqrNDGsQOS
9hOmGS6ttCV5sZ3kvpCKKtY+kcEhBda/1TteGPMMVx1R++oC2pD67NjUqgpMtRVp2EzRKkNuBgsq
pBeQN94MX54rGXFabxTLCobdRinbU9nUzwwdq5G5cptDz+Bl1v34cTxNYeJ4S4UyC7KiUuEbgqy+
ENn7GAdEIcCU9fHa0lND8Otff8dO3425RDbqGouIC3+PTTvTGugQGtVVy2kN5jBvGY1hk0Ty2HL1
dL+zAoYNfBW8f0N050AatXoHZfKIfCx8xQrVo5E3c7u/LTkqzCFnH/9Ynay1eraE8vzoLUmoTFk3
yhH7qMXg8MGAViII5gZiO8MM6S9lL+NbW9IpJ7vhkF2Mqdn7+aGqxm17aP8GbdrqRThRZhi5hULY
XxshZKHM0xp0Amdtx9or6E5aAtzm9OT8SmwsbBZ0zdDAIO4QBkGK7LkZW8jT2b2pUdCcOdoZNgem
KBvw3moNDAHn16RlZ4e3RBSoMAVWIdSwPx/F/jj9/xRs7Hai/fE49FNl2+woGNqy1o0Uoq86Fq+c
4KSZrI/Pm+jfWBPdJWxpbokl+XC2BR6z0/ltFcHwkwamKgo84Teot0C8ZfWQZ8ehGSJ9auG0Th0v
H7auJyQ8JHaDD+RMrUydsvclNd6YjQXQeger7wZn59VtG9ZR3Y3Ksw4YwwBHAwb6AcynS7Z0wniF
NnG2ZiUEY4WfZaFfoF/wmjyrnnUBJeOw0+ogAu89Ch2+yEPpmHDX8zpaQlRQcKgLKqCZ+EoSoHSo
SVU11OptaJ3exMDPgLT2jza18XlX3WoFBBDEEpC5vi8USIBskOhx8XhASdreSc2W5GARiPJQMfg0
mbc8CBI5I7xEV9jWfE/ZZc0oMa2O6SG7DedA6dVmNsXVVYR62L5504PsXCjlJ4dkjjphbnryBq12
382lUr/ywjfEyAKKLuvbUF0d2ggeE4aFNONsSeEWymusrSgbloPoUTjrMoBeHhdDDsuMz410PKNs
ycTsS5B9xnoqKRK7f3GWFbCwjJj0fiTz0SRAseZATD9shWQTY/GBXXB66oYHELMjxXZy4rXqaI1W
FyLZWTTUCAdGHQ8CMgPl/9FoX7kt5cuGy4tnRTdZLNviDdqFhiIKv092wV1UjQb4sLALSvCMRAus
diAPoglZnURE/iRV4t6lNYtmQtjqawB/Gw4kPOrcjHFongLdWVlbk0DEu3ySpQg0SqYaa3Tw8Teo
lL9oXpAJHmrZOLiSnNCIVtcj5HiFpWB+Y8gSgRJk9MDmT+7dvUTtnVTAZHGursN93DdHYb6f8qzP
44cCq7CBfJdBG+PlNWZWJC0XwKh8FuYh8O4d9QreElgXVfNLut0VCkBOgkmb6Jevmc0mC+j6ujy7
5z0wsGlxJvA453fNQ/Y7yYqsfHt2UHjLZjdyO1YmztgYd/2739Xip9rl0Pv4FY6YIthOEF5FO9jP
Y1iuAU9yJxwq2SnE8SRcrdNftZBzDU48ld11xIjaEoZdQ9wLLeO7Zcqi4SQjgva8SkpNqzDM0j8z
dSTetYShQsP1775PuNtFnHoV6GA5fqRr4kte94xqDwRJJx4QhfJzqbA25OFtX9nD/SdP19tlNYf3
kIt5J1eHkkg21usONa10ItYUZPNSHDBkVIlWOlv6jVXbsCN6gWMtJ8eGK1d9A1ibxj+uk9LsZKu3
0JKgw5+bdMehuIWcnH274YCYI3f/CqvyBQsYCBnmK1VtassOzdjqLfMzXUesWeW5mPzmKpq+yHL5
TDAjyvFSeORcnMxVWlG5RFQMRLgZ1Vb1G6InqUeRdylgb0px2k1p5u9mNcBCJ07meRlZr4zuElum
j/jWiMUe8nLZWzXyDKV9GEwmLuP8kfBQP2vvpEmgAODiLHoTxuDKJpJukg+88NBDDl6LvRZboQ7X
C2QbYPE0u0zyZdi1ho1sNOwkFvcnaMONSrVj7t4hWCS3PYVBcY6ncN8Fc6TPzefg0R99fH24r9BO
fBzJhEjUY39oSkD3WLyS/ggs/m8DS82zjICoweWAQLCVlwjSrRsKTNbCIdkUY3bHSUwZqD3UYuwD
Ua/6oUhjtpvMBd6BR+fi5squsfJ4mSMAu/rYjUFU2KR2x3Et2Ce1LRpg4vEqcELEw+7LpLmH95Gm
ErYyj6vbdEDLyK3fiHiFsL9rpF/ySN+eLoUU4XFf52rESdUfNvOgQMrOi0FbhPId8LoFaa3vsXlp
t11ALLYBTaUURWsZTWkWfA9LjVOiolnZGBJyaADz5iOnyF3g2+2Dteq1NDdV+tCvzvz1RWBEf/Yz
wo0swEPXyV0YpV10h8IMJtZyH+id0XiwBfYMt9IigUzQOkgPbB3E4pUUZlKvL5Au/B/HLh0rP0/o
5UjhDBgRJiHxWY8NkOriu1i/Yrv9PvG52wtU8h93GQGapxi71v9g1HieGoKK9dbVJvDbPof9aJ9o
aBczsSDeJTJw6fUbEIgQXRbjYfmKl9oRLxB7MCDPJWyiR8ZtnejPHn4B4biQW23lOlbGbR0Js5g3
A763+Wwd0nhO/FojaVRtgI7F15jgrf8woJYqe7s7jOxtYEV0JgJfkA45jjSLweNl2Ug7si4rvXGW
sVdjniX/PUpWeoMiCCXysuGggemZG8ap7D9QBAhKaCJgY6zK4U1XrIa3lPuFcbnFD9EbTheObfI6
u8o084pmHgtrm5aEt51OXnM4K1cIzCor8HLPLnCvqvbXr0Z/pe+MztpOjp7GFRYmhROQ+WGSWuyL
GuAp8FB7LZyVCIxhpNGEoKjC+clmSn82tZdV10dV3lhLw42x/hzvbOcBLMnm9fVESQkKDwblFYwH
dEoO67b5Lj4YjCxOE9TaQyKgZWpbhYw5g4k4/MPhKXC9+Rv8G0N39yTtoz44pC57laNqy+VbX6IQ
CkEBHVWClNfEeozEzY9ZWV4d5hn6d2Qo5kGfmyLGs+7q/nPeey2oS30y6biRhD29Kwu1Prt3SBxP
3Ky5p6LYNJVcmYKbY9eo9E4IP7UhcVIE4C/Na44QtGknZYSZy0ATWfVzaH9gBtxKrQ6jI3ffP81V
tYCbYmuvxZZI4k1yVKCcKc6j8+DgrTNZX28pawcdsfL+gKJVc4/EP6NWPx+59ks9gjWcYK3Thqst
4zer/ja5fy7I41kO7+Z5mDydVUYj3BF1Ze48yJulwfkFtWE2qo6TtbprqLm/9puevWoaPVOHtWpQ
mCrAW42kKisC8n8TBYwPt5O3lF7OC5WzrQJMAO6iLz/aMXYqk4jDAdXujgpzRJzR/ETagjm43kmO
fq4CAv6hypywD2vXzX/HFBJbK+RN19WG6sEGFJjuusKJazEslQ6XoqXpzGjOPhxIXplNrtDozcVX
KImkMq4UBMRNvQDWjVmJb6r2aWYFPJ04qNgwVkIvs7X7RXalJoWMHAcUgUuOWNfgcoCYebKZ3eIy
hYIMuWpRra1zi7h9Dnbo95ByR5tCPNzeNnWZoc4acR0v/kgQv8VLgHy2Zjy5h6oMhLaPa8m6sVkf
JN8Ls0224CfqF6UyxUPBENcMtFXYSPUmMWK3dtrw3Nio4u0sH9U+FMIY70HG8RWQ7NJYJ9lmMdUb
kn7VEuwsKAOK61bAyrK1l9Q3+HEVXHPu5ba40/icbOK/cQI5POWKxpKpcr6KI/XlrA5fe6+eufaT
csLl9AJwu8JHZ6m5pTLNy9h25Qb0vNKqHqg38BPV/dUp0tOvRsVWJnML/RQN4IFNdsfnNxprcWRE
V3FIRUQd5cmEjQ5F8AO2WXDXKyNfAu9IETbeVQ0U5W3IZpnQSmDONfbV2yz7daE2FiGU4WRHHqnz
2uXpz17d9QQQA2CMNw1Gk03O2gXkXwXNlzfbJ5MGR8Ds802QYsqVtpCDPT3qQLnSXvaG8xu0ujns
TDjE64LuywJYS6Xc7VxvBT2oJsQ8qp/QLBAE7AgaP45+Zt6UTkOjtYi/6Z+wVzj/dFQVDwdgsKwN
PvGHAspSlG38WfczWqpIQyRfWZg3TuoF9vOSzLoTYc2W5BAVP+gJUaVm/lqllX3+BR0up97R/+Hw
Ok1vzis+z6oCSm8YOTiTZaVn/y8/s5io7xiRyG4XZ1agqNu9CaShS5PsF+qY2OyDVquFwW0CuGiL
fyFX4SujtktPYg+sBtePSZz/ZauRDDSj8CmY06xmLWQDEw62/GWqaemPZwzNP2OmyJ19jMpF8AH8
iIo71wJXgQwsqjBxZnFY+t1fSb4oYBtGmnH3zBB4TTlclwhUNk2fbqh2dp5L9ERFAiSRyTn0s0lN
Nv8MwQSV7Glfl2qpLYHZvOFr3t4soOA+P5kOj3jPyWpnUYw706h8mL5cqW+efp0GcnqvsBUNTAlv
TqtV1cP5yydRpUA2obZoT7FFu2nDayOxeJQIXN8mpVcY0lnjUGb4hmpP+WTd0RN7d0VeRjQ0MLBZ
moXgHEbqVnfrHx/nddxgIAAWcrP7x0UoLVOjlnKk3FFX2PBlNMuFlQqjAirU5FZi8OTSBM34E7iy
SuZx5gGKHrRi0srvWymeOWs3QCF81CvStG+9N/NmMGg0OnHaAYhLomHbMnJlYXbDiRTMam9v6mjA
ugG2pcny2Rf0nC3ka+OAIIxERhchIoJnusuqUP0NiFgYs5a4Pzh1bFATcQGVEmBIrEU3y0LKkXDv
zqD58HiRIzJA/Yq2xEGaUuaJgR793sRz2ThA0tqCIwz0Sud6Sde9U9NREZ9Le+JWhrVFcMxmIsw8
z/tpeUcE+3qnnWy7JHKB38vsZhDbg2n2FRNuW/t405nDzFj6nhGCbKJmTP+UDDeweTuaA4awar1G
mt62hz6e2VKEQGpmSzKRmzX9eHbuCULQ7v1lYRTpWd51covEtTvWUYuPWWUTGL95T9i5rJkyvA+t
149WCR6byH70BR2YWvdx2BYvybatW+qPAmvi8a9iE9MYvFFHGQob4SnM2mTY+n1wq7DAiP9V5DZ8
a9WiL5oxrRlOnqYdnprbiFWy8wYYx1yqqUkrHhxEm2nesigyoch/rWO69/XOd3Nm269CxgF1XZF/
jLXbfuDaNopTM0AAHK3gqC0MnqYGMtNnD7r+OuMXyWDzxP8PnwNxOx4QR3TZgYYeLJaNZdx+sjHf
MzaAPu9HKdUUB1eSfj+n69B9268u419QSPw+ZlRqhOmQfZxFzZQPqrk1zMDUUXudwQNX1Y6G9bBN
wKaUuVLl0x2LUl2nM4wjAkayEA1nll8MyqT/kXFRA4KO/7puKNX4S+idDlTXGO5Q42lh8uxdqMLc
EYVM3J1EK5FwYHq/gu2/n6+DvsTiOr9BziGts2nbk5MQM/tRkLmfS8TT7d3yyVem2qfxnq/Mlow3
pUI+63H3OEqthpq7gDiRr0SXdJ21rPe0JcJVYbNIkKVDNwmSr1PTsQDGu2wqK1/35zUB+HvMnISp
R3AFhwZ/2SAerk+6dVQM8ehShETSLG9nKx1FBg/4bWBQuv+a8Ulx4O0ilzblS56JP0NJAtW25+Vp
tJ0OlwtFZmHhemO0f0Elp17rKE2p4TydcvO/1b9EPRuu1S87hdnvvsFgE9Ik4G7db6jZpQ3L3Cep
SfUPVvomj1wejWV/IhhByyjPZK87avdVzyUF5WnzF5LYYz4MFUys+FOmwMYil5qq9w1nQFPPRjPz
1s3L73Cn4rxLeskbCubEZHqpgKTStmxxEq/N6osDwoJUUryq5ne+DyAb3okfLr6fdxrYjl1ZO/Rx
M8UxUq+vAs/ItMNbBO2Kl9BOXbOpy22vn/fvBkIcY5E5rxDUYznpNfHf3hG9QUsV/Mj8coRy1Tlb
5MnzV5UOJeYk30vYWU6dXFc+noouqbWXVkRFi5Wbi0EmPHTvZUyooyQkxwR6qd6Mah3u2hHtAY4O
muRitIGYopKQJeuQ6AgEEnFzgrp1B9YVnz+iQc01eXg4E1onynPBoDozM9qGwhiFTGjpfRodWxQd
l3zrpwssBtfIdI83eWj/+bvIO++Ei4tV2/PLv70xme9keo983tyrCtVcXf9AmVItKa6ROfp9+bLg
XterADaeScfdsEAiw9ER5bnBJmmifI41i0eEaU8Ufo/CirbzTEQJ74siXX6WummrL9NdkT29s24H
SlaerKmwWkWDQ024d4mUM8h5ip2t7Y01E7dHQJ3XwBbu/tVwtoix0svAyTh1ZOMp2fyWnD81WjUU
87ghWZSEtSZqJfQT0gOY6W7baxqC7p8KnSoMgbUWXJs+djLIet1nk++ghErDsVYj4WatXDMG+aZh
RRvuruSNtNJJCORCiF5OQgLpBDtI5F4Dv6q5EMN6Mv0Ya5ZOE3/BZ2ABoPWqSJpvxOeHgQMawcXU
JUYv3lO8w64aMlSgAiMY9WPHtERBgd/bOVfVtGlZk56qTd85z989QYMhMcLAfh+t+61nzY+LxpJ0
PLzYeC6gmjSR3bCvcq6DKcdNMPu/tW4F7tBSpO2zuzsbJyrFoWfrAUIk6X8llyKeVMsjpW5zmRYm
/Zikith31G2P3Z7vJclgy1KpulHhIS3Da6ryYYhVA2Lb6tjprLLmQyBBH1XTr7R/80QDpe7oTN3t
3PBaIs3Ao+6C+qR+5Fy57/DkRsZB9dyytVaFL0rsUMwotEvKi8fUZLRM6ZiYHvLzZdmrS2AjhB14
BFlskwjTa5CjGX54Kdw7aK4ecl3AAqaZ0N5IhFDF/eLeKXQs45kY/2SLfhMebrs6W9uIzgeuMfud
ZhykDKVsh9E4PvMcOmZbNR5AzPr3ib4ENu6hmXAAZo1D802uQmZo34pRkxDkJ2CfCiF5o9L8HiWx
fqtIcstiaw/DsKa9W8wZgndYVd/5gT9Fv/auAMx0u58w2GqbgewMqJEKHRrJEgY7VbK6nRHKi4zy
H+dCFEPm1XaYATSs/IGyAZoh+uRBKhU4aJSQ+QPWExvIAgwhZWzvndLT7b9OLKNUxA6PR59oHxXZ
ObgSRPsoT4RmyZDYBa2DAEKVavBkXCaApz0e47WwTnS/e5xnrvWnB4XQXi8rJDnyaISBdLAQf3Yl
Ck76ZybgtFCQNQ2IOzFsovyv6gMF1wiu61iotrT2Yoic18attnyJrviIkglRfNIq1hXQCvEaz/+I
sOhEB6yH7dCxoIMtCRrkFmUytT6kI2XyAFW5fkYbZpb9LAcpTUZlT2dWEgmEc3q/jeSUo61zrQxc
cqS5eStvXkt5TParUDTntDn1zFfbatw12VvEXp629CDn/9zAs7QCYwu6jf3q2L6zUIvkGSR12tj5
tXbC5DEa1LXZKfkxE67d4jzxkSRwrrAuMzRKcAEjHO+4xx9VqfQTDPcFa6i7gkY2Yla/p04XQYZA
6/2esRpoAPRhknqbKYQuN963EcnPasePb6PgCD0oPMg/hqb8o5MkuZsq9KNdVM+oSDNGBGBzWOju
ANMymjg2bv9As/jeIH/eUJSNVGi2GtnX5LVdNoeAvqF8DMk1S0Er0NYpEDD2X2hcXGnvJJ/Gb1Bp
iAO3jDKXiogD8glx3//ObJFkkIff9uE+GohlIejwfIGT/K0WShLZ6PD5r+xHkDUQNUw2m+ZgE1Cx
L3+IR7N/SIofAav2ASayg2Yjl8jWNekYzs4AEvQxz5aWtxY3VRboe3ErpTYeX8UoPiOXkc6khPA0
kkZCE0sfJrBazPANVldwd6n80mxY+LiEZXWPuydQweBXxpwjjAjWvJIWPEImlIQ9ymAqdeerC2yN
5d6qcDJ2ZfGgtkxvk1mR2ZJhath1I2vlgtFt4p012UoNAH5OVqz6TV1Fv7D40JMaak/Oq5GVDqt4
6CQjVge3bvc4JgQ5BsXN2i/GhqOp/fnlz4CaE03FcEPdQOxgOO1BDhLycolYJKa77c7TAeHsGT+F
VhLZzFnfQZIvZg95JwEUt/UowBQPAxBC2lV/7zS+YdufimQWL0O3fQiG5+m8fPpWnULKxT9A49+j
h3aOolIW/RcnGNrHPRgH1DLqAtCx9Ike5jGLlGFfhh+Yrm32PYbr+4WBs3gJSkueH0f9oFK1ZTuh
v0fYOU34x5ikd/0Q2FuY7geROLq0M5ilBvY9PLv+67ydL0RIuwms2HjJJEAUjIkk5tJV3IZnFvxX
L4UoTUytviDxYl89qFNFMAkz/JeuZKd12l1wnQ08mesFKcbJ6frIOOIN6CQh7iH34NV8uYoyFpzU
qFAjAJfAacHpUrkbCw0nJJRg9uY8sS9X29yaa2IVhTpSrtXV9PgSJGlj8ljwcfdyULo0NUTdNlJ4
ZH32HrNN9jJ5ZaaL0lq0yS6GBDf/G1EsRK+nN4dO6uoFCpmgV/P6NB7sQuZK7ePabWKImwm68WSI
wdZnBQy0fULDD31Gqv0/RL3/8nPAxDzEO2e7g1IVF6uzb4sPkr1xFWA1M8NcuJvPmwrFN5Hji896
rfCqJDv56E2RgtcxUralq9+bhWvYe8zPCFNfg3ptwJylLPLMMZ2dMUbfeZy9Fau/3pqJBCpkl798
DLOhqkzMFwFTAb0zh9bdMyU3kZ2MU5q2EcK5HNE8GUkYhSVmCneUkFIlzgTCIq9XsQhwtBX+MFi8
4WW26DDZAGDOozWxGU+I6zPrt4chqypCnxr1vYYFHTQOwopYD761IJnWCZxsXew8+diJWU+OpR1b
xhznYVDFj1KIp7vusoHUkCR8SM4322sSKOkgsyKBWQBLjyaqROK02zmDvApHoT3cUKS7Pptdf1fv
y71D3OqIAgwyKIQke+De8GEw8+E1QSKljDNBAd5CfLHWQYZAfXkEakabtf04oaa+Qo8U0pu8+q08
xxEgi6iVK19eF77puyNu5inD8//gIgixsfkRsqXBkA3MwaDHFT1XGdEZ6aL2/odPolwcN+Dqv2Yq
aAIt+7vSXILEcfVV1H58NG6JswRsZCGEvQCPVrg1zALv7lb/541YsrEK0ujkU6prD9mCcqRByUL7
uBNLqFH4WlKSyscqX7zmE4twxGI5r9FUfPYfanMP5Yqk9K9pcp41xaPDof9zkUaY12qSerpknter
iezslWe21+cveTDon67PZ8NulKpTYmQmT9BcD5NN0zOcIa7LRoY1AO2rCKugYM/8bjCplOMZGvLR
KE3iGD3rYyfRf1w/m1bdv9e2xBi8UTBvZ0oHC0VxqDzEsEO1id5p9crhITJznyzfWXY0JB435azb
bTECIgrbUtHyP1i/EULGItRxH3WG0GLso7DlCj8k4foj4rkxWluHzdIIuEWvV3376bcbUYeWkH7h
fhUNETzBMZigQXUca3pIbL17g03niwvA5SKO21LzNclYKSjpCYlB5G7FmMB2bTTjPRMhHoZqZjg/
z0WYUyqLEktpPfpspqo8cw/IrtA25s9Kda5BgGiGZRyAlkNCeTnlUe8K8Swz7xU8qp1eE9GH/JZD
u6myCEsA+ZATB7gEl9mPNYpbJ6n7Oq+l20HPg3rZzAlBqsrJ89cao8DAQL9olkeV8kxTQ9ciwa3x
+c1O/+SpjdIqf4nR7Y4cYVejAMrYFMSl24LmK6kGsbRlDnBg7jf/4cxh6kGN6iSzlhb6urGvu5Aj
BWc+CTm0DU9u4kcaoTgR26aLxf+lmgUR+hZnPVH/jSYnhqhzLFFxBsv5wles5I/qXOTGv4rP2k3u
OBeZHHB9yVg/bvKWyvpjfw3sMlU1ulAlM4yXv78sYqiNqop0ANrcRb7snIeQHrWxECuVApbwFt40
XTj4WVfjj86Wxt+Xyi0Kl4VbsJoaHtJ33F/0NrZE4pZH38yalOGK3W0xB9tQ7MD5/wSGfM0DgW5c
Fp9bPphNkOhqVU9nA8e62ghaxahSccRKCYDNttSk46iX7Q6kCjHab0/7NdFDtIKMR1mrRROoT1Sb
FQp9Ss3EtFQnlo/kbA4TWw7VTeuvPO5O+80jQjHdo9LLh67E46q8OVGz+b2hHX4PneREnlruLN/j
4n7KfQDgni7M8xqYhrgj6ZNkclisnjglD7LGwXyDWrciEC0q4vIMgFG3hxAdzIuj6yCdLLjsqi8n
Rnbz4towePSLgJyikVPtlzlnhFvqBFEht+sqjB9WbLZoGjRzvOJnceXnQPLAmhrbhhTTSOPbx8qo
v/W7M7GL/A87vd7TrHv5QE3YKgDkkTM2szlufiaBl3F6D78sNYZuZ6JqyC+OJ1PUy4/Hq18BFuwq
kf25ln+ObXuTM4MpaOrImVcOA+MvZd0bGzt6MDeIpKnuyysFBftuhjYCZSmmQpxeKPfePHkAprIE
i0p/mqyDN/hT8CnMgfnbAonfwl70SlTLO4M9KhFO2jVitTl7B+qc1C2aUjsAzc+XKJOAFoI+SBuE
rsZIxcrq2f0159bTRSmGOlCiUyxJIfqRwab5diE1t7MreOZV6g1ymw192nMWf1kIOZe9afGEtaxl
h8zeNhLOvtoMLurG5e6vd32D18jmCHvmcEeS0YcpFucqXdTZf0lnUmF7QYaqnGunu3nllqubHxQ/
t3/dhPqTt5MVevZ0OfZr1UeL39G35OphDhqBYe7Y7DTm7hbytFnPOhvfsBrStRYkzwJE5N/P/T/8
k9b2X2CXbJ4lbd+EYx3aYRDylP5p6Gs6qaLj2cCkCcdu+Ah/wkIygt2mSmP+8H+haKfUxLT4FyBU
bJwagR7ebvbgGu65ekp4h6qPqwqaJATy3/518tkja8JxwaM2wq9NxhjyIdOAP7bYKLL/QXQwFpqH
0vUNMHALgR48On0EtA+W57l/aQXfLJf0+i/nRFLWNQJEpfm3z4eA/KG4U7bo5P7PhqG2Ok1uLiUa
lzsN5COo7PyrEZLbjM7O6cTP3eqSYfLR5BnXvTk/w7yf57CIzzIy8DFwHFyECynK5v1UNcH+M3qA
m6NLEyM9gNPzZu+/HV5jznQlgJKuJt4isYoe5udFxuSDiVnSRbMGcStwaq31CFgpgr8gikOfg0a5
cwbLfbSaopyI4DK3TPJ9qzMkyMYQEuk8Z4VEGf8IqL2//yHShYjPKr9uh70TKng3GtjPCsr2RVLS
VA5/duM98G/I5juWsugQrlaNNVVWzHgg+aarhpTxYWEI/Bbtit0kUThn/nO6rS5V0ryB6FPILUlm
DC65Fc3tIm9RZ1nWVDHPxkt67nDco8BHnNA5s4dwStnyqTkzNpeMKxPNA1XjVkeEAs9SuBFq425K
Lu6O16zFAg+UqDv9P8S9IMCtID0rXFTseE0QkXbD3rFXw6QFEUGqiVQGW5DoNMocewUSzyZ2Sy7g
yOTOvt8ahqLKfeFaAk8s0YCA3kDVuMqIv2CbnWppDTSZnqR369V8XNuh0+Ucv+ejQ7EOm4YfBRXY
4NP0liHJnmQ8C/f1MPFUl9lHRMgAoxrMpeCdk0VHG/upaE607qOd7cmNCTM5vsp5Aq3qx7406Kk6
8bIKFSwl/HzNVwk2A6Q/GcjeCD0+r73+YsQyxcpPvjMWJzWBAkR17OzzDPjKtKkHsFHpQ9+4hgZq
f5RjzKJSU0zbHqobU1kj9cgJefyGUGBmxdNmIgM0X5L+tY6BSacEtpgrDuXjgglNx0DFlroSQxL7
7JRt6AGlWrp203joC+Dgon+xEFO1yLXeZ4biStKvo6quJaoE1zbpGK2Cv0Q1AY5AqvyzXcQKGJTN
MOO2VGth02H1qJILRUSAnEreppRNrpAkv5TVGcK8N2LIvgWLe33MKm/10jx93P1MLINqkncjUrcj
4a7FK9WypmCSHZBIhfvCAd6EYUvz/zdGXVA57kjdgpaAQKvppARarZUQFEoYgzg6bNsALhFadumd
7SiOxqHWKNtrXk+nu8ie03OZvH0BYdZC/M1JrO0TTFUxSBNPZ9PMpxmV1Jpz936DP9J8zWirhDKS
S85RAxgqvs3VT7efKo+77URw1s1wTd41gT8Fy6qQijJ+40gIjyPmsvJq66utoNpy8LXUuwNLAHDL
v4Zvx2/V63eomclLWdm2mt3rD0luXoyfi37zSs4ZVYl7DuGYXa05FX+XONfbwnZn9gAAemFy5Gzv
LCdhgz6D6N4KtwBF+I3BkJrO01TaUqySl0/mo3QH9sTf7+KiGcClXxwHOJFCwqR++PlqBPwTolHa
9knMJG4p2xaJ/ypbubtFWPNjVyLCUVYCP5JLSWxo6o6MtFz7n159S82hQkn4+RJvhC2VvAk0P7zV
BLrdQP0cniZ742UB/fuBroS2vLTzRkPyBu3MqWJ/gdleao3MQivd6DMWakhPl88d7oYS7/VSi13d
DFD8D4558aacYoHUeloYKho2tdWmTTpqmFoHLpaOgdyQmNrHW/zDQpNepThNjooUousSIamOfDhL
lcIJGc+AZQWLkDvSx9YL6XSoOLQJUh++7ppJwKFXKIJTvxyTQ5Mcd1CicRnK4rMq7j6qhsV26G6k
QH9PweVtqiD/TODSRNfODlGvjWm5D9J1PnMJR0mQoqooJU980p0YBV4tQWMjMXBYCQRBX30ZBknx
Dku4jJV78HHAZ2xJJcazi8hNtpuYvepBv8a9blBPeax9S33WGCX/KyaCnSjlR7TBveW8MkZP+ihL
JToZRBNp/+vfRLw4ij0XpCaIH5COwXKgqHwedx6ysO6bX0I2jkG3ErfMJrPt6nMAIHk8qU59KQDp
hHMNe9eCrF6buAWpBs5vaP+5FUgmSpyy53GwNkXg9EjsImqgcn9sLsoqJnE4WbuD0rnBAM+5aP4h
9fFYSfK1mTKwnzyrFGtGBgN/E1xrOrwt9+N9abZWex4Cm/bLqUkYqRJ7+GJFQicgzV7nArV+zT2O
FtrtzplPXseU5jfLDmKWzDFy0whbvXNqXxZYGBLjJCErVAHnqg2aucz776ko41o13SbCv6DK99lt
aHPh9kipnUo9MFX4k/QFqW2QlskuUxaL7hQ9Entg1idMcCrT1fHk3L3ZIykd7eBixuAyMcR0tDEm
W/0WuwY2a3XpvhGBZpj0jqLpMn97w8RX33LIRS0djjC0GbplnLi+pFR9VXUl1DkAlMJcCyo8vRqk
p3qx6L2BWAfI8574O4zGqId/P8q92cMYBsqpNo+J16AAxCYJVaM8v36aBpBT5va9R/vMt5xZvVXh
TZxD7oIdPtstMDIe5GltmzLOjxd5h5zJWX4K9K0aJhnfaAwi25c64594elRhvG3dZuv4i7q/nNCC
zUsSGZRBtfAWVZ67Gu9sgkcVJ593MNxRukmS/nOgm6HB9w9/yrndeHoAy+opSjiFTzcIWjbOMAhy
IDCp8jPncoejbAupXlKosyNDbmg++DYfB2O8+5j5FPKT0b3ZrmLa5c6diSpdeoH1noKtjoxIJP/0
zFSqOYWBdZNnaQAeMYjeW4ljMtjwZZlCrbajKSS/QahEVmt6n1Hbg7FF4nvjQCapWAiFZ0v303Mm
sKSFXbXL/VUiRD6dzq0duDoc+V87VllGHbBcMEgB+RjmduGIpG+0h3yIIapFYhLRQzj0X+tEAaRF
g8igSQoGwsTnyrbZ5f3AG16Y/XD2u/sQdPXbJq/UBq512RnoG2Cv7bgL78tdOmtj+jadDtQj9+Hl
/SoaQhGd42ro4/8sUJvZoUK9IKLLdaN3qZ0PcMWbU65v1M/7OkmRqkhgg/W0YQ8+Z5vg8jtwIj29
BumoH4ulG9mY1lcWSzcYm1glnK0TulnrMlydYd36lonvqrljPr8vLYlGjEOmu9bWLH8XDa54uM5K
gJ9Hbvi0DKSOFRzs1Cgak3cqyWm+QtLpgKtjSQDBBBEM83j+Asj1RAxl5xwIdYzJXXhWlbaN5sTX
4AcqFeJ/83q6S6c5QYBNRFVsOqKKRq4e+NjGIiJJJApZ82nKang3KZPFxXHmGBkn8XEIM962DEoW
jLUcePyyC6Z8r3LgNvCduN/0FNZDAlyQdebLAEgpcPswW64CcZYweyH1nPjMCZ2ROyZWLAGWVltP
/VwsNBeP4MT1av91b62H+FIIPL6h6ISEelnnsW854YYLDLCl8PdkdtrauUmfHGv6PG/ryrDmaWO7
vkt7MkEDW5KHdLMk+LqfPgFOvKiP6pUmIvRJWg4qtAlfCPkQYNj/7BYH8TIbpiu+0xTt7emuSYMR
mWEaUDegLf4gkz64hxuh8/xMRBlCQbRXRJwL8kl2YdFPfhCUDnoU/F9FxEQJU5a2ia83wTfoBiv1
Zgi/HFJ6AE0Zjty8KM8f8mNiCjG1IGmsI7qlr6bnRGaxkfR0witldeXnCqi7vbSbRUI+2vlcyPtW
+dmRcJ1a2/Jbsqb3r76L01VJSRSZHRGk7xdYQCAyMXjmBkEynAqEewSaQ/bIipxk8teUuZOMfb7p
Tm9boG5HoyYDyOKbv0qzDPAPK7Howe1yfAVQb/3hRnznl1ESEgYxHMnYpmwaPF9NUADhJMV7AQ3E
DAjlFe+RSLeLjtUSGvxj8uY9SVKiAronikn0EAvRg3kfE0h/zmonae8h17dzl9r2KmGruEPdbwgo
XXB9pUv7wrzAvE7KLci7S7p+UCSjh0MYQLZcmqZlcQ9Qp8IFtflrjvoOsCFxYvSWKiUI15bDSfE8
Hsm5pDkk0YtIjuioLxbqkjOIgk4zHY+LQ8/SE/feZzsHEI+41LLPontAiqymCSlxBZyH0e3VFAJR
393oraGkfUPb3QCEPlUa2wYYWOmvX8ZWl193kkDXkvGUpQ0S1iFo0iitodSzCFSDF1zx7TUBt7gG
hG+HqGo64IEt+HbEAqRjtrTJVxPjIKtqL9JgalE3zjP5+KdvkXwm1RAdbx9QRYNk4oeLZIFlt6IA
WJ6bWhlvj8LFElNyVGPggfbp81cJGkgiivrrVm8PbnxW1uFPazKnS9APC08jfEELUbcKbZfYgftp
UVDczhnsLlacoLTmY14Gedm4cTGb7f1sprmKsSIX5a7vDPdn+q3USExo0UrBT6Ku0KQcpE6kJivY
98mWrNxabAVgPIta1bZpZ0KN+10JXZ0zKRt9KMUD8FAP6Hrz5nQa8PqhqPo/rtvYDsIicXO2hiKf
jb1018uf7Z2feMK7bfInSinuPwyMhoN0s//dLgI3NbWjZTn+q/J9nrUFz29kv0LcQ7y+G9BX/HM6
8gVC87i4EOJZoCZgrdP4ZQDkH6DbWlUl8dBIR9vFaGMiX/uJ7afq2HzuzSOL/uQaYzABXwvp56hb
mw17hMtgN8JG3HUEu4PZ+VmLs9i2YK4UkWg+yMFcK69vmw2DX71LTHW+1ZSS1hFproO2xtrsS6qu
xqj5PQ2BBhDwUvQg8Es/iVwOwEqLbYsc1QyxKiz+FfBKMA1ZAkODe6uNChskJZy4bAFwJmjt3Q1A
hi3BvgQXCd2bcp2Yx9koWPMRLIOPxgkfPlhRUhLg/yx0S7irBmPjZqannLKjnYPjNI87u4XJDckq
As3/L7V7ff8lFX/HdS4nDrfjNVuE4d9Et/I/9DX1nldxM/3tJ4uaLlT+6f3erw7Of2zU5GMkgRBT
hBxJ4JqZTilwoAr2pDJu3cw35ivJu8UMW/Ln0aC6qfBJuQpMMJJgehVbouPkDB534A9AyWWaUt8z
jJtrRAC1iJb16E3zZLx43osofe5V7GWy9sjqyr5zkXNiT7f4hiEcUxMOGFa209B8Euz6v/1ISyb6
YsgBp+J4gR4/nbM4THi2uA0+7xf+8YrWGNsZavcvof9q1883V2cAl3HSSvBaz6uK9S5eGGilIXyq
0VxYCW9ZJGrSG8KRojl057wQDtzMp+4fCAnU0bFZsQ07u0EMe9ypzo3caijjHXkQvyFUMyiKiNH4
faYU1FCTgdW+6D9yGP/B+zjy1a/VcGZ632HKCMdyt3qTawUHIOCVaJYq5YF6oP9JQo/MtClTI9tK
OjMpoZivK7BZV5w8yn94jpoF4L6zOyqZ4XqYfRkLtIB9jc0xv2weHy4xPftGeZqTc1jdP5d9Pxne
dUY0wNyIGg4CRdVIiqw8rfEF10WnbV/M3yA+cJqfU1Ag/H7pgkL5ovneG2ObB46v0ehKDGatqe5B
MLUXxe1YszwrrdIfybphStaPQ2BFSlowmzkrfX04A9vQEWpMmfF0OHA2V/sxip2O8EJ5zQHdkeq1
e6oOKY5u8rjRsg+XZxeo297I9dbDNdH58L7TTPJSud6YAeK71ZY/SXPQqZV5Rb1zRoTqEpvtD546
W2cD6yfRh9RX0HqUhABf6C1KG1e7IwnV60nNuWGBCNmhGf+XeM0LiOnxQbUpKoWGBPyhhPniFFuv
KEf1hztWa25zLyd8gFw6vWymfO2fbpO5OyQuF8iZKiGJ5QLZIpwCx3eWheMxtDJ9vL2qmZay70HG
NzJk92/0WXSCGhfRgm1ONt22bQWIHA6SmnaVJ6Nzmln9qQc6TNT5q/Z8FGVobGRatG75VPm+be6D
uIeamc9iltN2yJlFKPkfJZ+48r2cVSj8m3CnDie2KWPuOW+GCRacY0Liq5+7I1ikwXTbr15h6em2
SrsKRc8gpMv9FAWgzW7C+xTAv4ZzUWcI1rOdjp7dagJKl3Pj34c+Nk2MPMN0x7QOumpFZ+ewO6Jl
noRzx2tJ8ZII/AjIDKZN3Plm6kLy33wUNzHNAJvjl2kR36ZduVxVV0866zMoya4hdXcmCAeZXhhW
IzqzdJtEJBqfohk7/VAsi/k7xfUE9Tli8y8gBCQCAEOaOc5m5RzlbrhTqnEvO+dMxwB1H3uEvmPk
d2iuTYi6/3pqiXUfVCaAXv45CzQzNQyPuJ7BBHyCEtt0fZtqmw2OCApJhI4g8p0XIaI98xDvYfLx
8Qk63GJ7+z4z4a6La0/qA6zf7Kk7u6tASZro9QDaQUP7pwYUGQneXSOg3B7B8qUW9cVDjjYXXQPR
WzinfIGVadE3G6A2nQKw4gv6a65HCBlq3eFIS6JpbH5wZrZsL+R5Qxv/fW5CYG6f1GKxFo2F7zkF
6LCLBbyVESWitJmdwhbYZffIqcaOMvOCmEPUk8T3ECg1q9nNPWvcqTINuvKJBn1gs2J/TQLANJA7
odpgzFoqBZcLeCzjgNqdJjWvkdM//B5Se+MptvII2jnxHnjFmCMIi+tSZMT90+1/9FD3ZoODlS4J
P0Ouk/EH26TD413tNw628WHMiK0NAoJE6QoJDEY1jzKPHJwyTOyEqFKb1LWlaJ3DoTOcMBR2VLeb
WuRgMHwIT4SYnZJe75LQAPEpl4Rb+miF8+6QCYbqeKYXC5bDOcdFNN3fOh7NlEKwaH4Z0/4ZwW9r
AP+g+d1CGjRfaToGFZeW7/zCBL1Migh7YdKz/5Vs4qJLLziHEh2FGioss9DQmYAxc2BcerHIW5UR
6yVKUlEQ5N8Ye+sNSdzeX9lg48/GDCPSs4Yd1weOaIiyurtFN5cy9+LKAHVwrxculqdLOXlCBt/Q
kfP3YWvefoLNrj7dxgsiyEK28TM5B3vPNjB/1UjCUibyvL01JH5/Z3/UsniRr7j9+uDkgDqbpk2R
5FPBCpnCchzEnCn+958PiNIHB39nYUzPHaxH/coidSImGCEM9h+LIU5ucpzE1hZ2cbBoD5FGheCL
yE6arbuH+JXlgT7IJxDcNYyhOBIuy8Jran9g1/O/AUAsDNFa2f4A1DWdavxkW2IWrUEX1EOK6dky
ObKtEeY9BBQEUAxDbNRpVCZGJUTW6gp+OCKz0smGLHuWFL0nd1v2QnA06bGwCNoJljZksasFDCU2
5i3JrEwkTOxKe6ypDrcvSdD48CIBZvaWasH8gIYVIKp/XnZ7AZarYsMr4IGSXHcUdy4pnIrDPMqr
fF+eJ5PvqazhPD2yiI8niU0J57J9RQxcmjFaZ/j9uWKFeToEQxHGCemov2BUI/meOt9EGicR7pWC
GwMhHQ9WYETyX9rF/2kIcBgE7DiyFhPq2h4fpYj1I57bejYJ7yEuWBx5fs9w06bqL/I1Mbobk2Vi
bEsEEbLX7LnRLRX3AyFR+c7mRD8xWlmvmWhWcxBGX3TGfHFwgnPwqMKlKmOTveaeQrkP87A8lix6
/VfPa1Ye1BZTrBfh1mFKmGKRzaQLBcXRES3KQWwL7eXq9ndCxZ9A9icDfGbXRCcv1j3mUiIPcJT/
4vrdrjcxRQsnJWN7g5cQ1DyehCmLxh1mmrQ1cu2cdMyc+DOMRIr54/v7UrYHwfvMTgoIQQ8l/9q0
ASLDT6drgbhG7EMVDvNo8E2joFxChWiJlnoJvtkUKUmfw/4s4x5bT44JtKn8F/RlcG1eH0e4Jue2
3UtjmIuZWg60lnikOqJQLPDKb+6pe6lH3QQ1ONm0aOrhIzg/tOalXCAAVkrYC6hufp+n8u9kT00E
nt8CbyhXxQg5YEbdQhmkR6yjQUiqk00l81Hz0qnBzm4xccUeoNL5Hgn6H0QPT8TeHwVra2cSYlc3
nwiCF2eWb+26AWhekbeEsIqHN7Y7K5kKpfdrRVqPCWBWW0APQdXC2DMzoyLPmHed79QTJTSez82D
OT/g1gyHb5WFUnr7+LyJGAKI42Hpm7XR9wPpgBxMxfrYqZFZnJ/PdOdJ5CvfxmH8kOBuOfaEij7r
abKgiNYrqKKMdMtDzMlAJqD6imK+biqNeAt76tDvdFyxZhqdFzYMJi+FfYyGgE+GSsozKpw1NUW2
bHP6G8B0EGdqRzoB/9wEKYKqtSr813NtyqD15aC8xllv1UzrbPb55GK5AMJPN327R3MMvkQWHZqr
CX8St3jD6owWiiPfdC8W00Q6rehkA6CBsRWYVN2ghYsFAzU/JNuhvdw2MKA3i6J4CE1QQxmb+stG
kvy2Gn8uW4Ubei1DYgn8zYr1Z82YEwxqGODbT2112/ueIFuYscaP5i9Y3DwCasXjgXhFUnc2c3Pz
mw7HCVxnChhtuv+tcFl7Ez+dUkgHuMGvNkboRsxmH97R5tixip43NYzn4VqvWEFyR627QVTEPn1p
npvAIlcVGYfdCV14NhE9YKLWPMGjpVxbhY05xjCHmw5eX0HmI9chHme451CoAaUMOH+eIOibSHqv
X+/gsYC+oHAqxHV2t+Dpu10nw2InzdVpZmREaQvLX5duW9i+q8SYVJzv/shT3vpTh/IY7RB572aI
9pV5/OXLlQgt1mkPUYsBG4HKRA4CQey+Tr4yuf89FleQp7nV/FO3LV7liLd1CAsZB4BwPn9RezK+
4eNTBZyPKvNsWvxUmVV7uWKvDl3Il23mOAV/JFoTGrKLlhl7D4ESkn4c1gpW7+vda5ADOp1slsjh
V8FBP5IRKebQ5Q+ucsf8TrnKH+3HxMPn5Vt/Qx0SxK69RW1+cz1Kv+oZzD+zi/2yEmTuHVy0qZqW
6AuM14wroSTNYcAmEJl5KHA7k1nJnPwEUWseRRdVuuUvT/Aj3cpA4HXOhfeSdTiqjuKlJMgt24q5
dO0CMVjHCm+Kmtz51mHMfBsbzyMu6OYF+QqeD1ujRozNB0eitthYJURzOltPRi3/aiOdtjXiRuqc
oWOfAThbxUPwjcL/U18uREUwn7x/qBEuQ26n3jJ5fnV1Q3Es0PwIbekZYochFIfkNlbjEjs92Rgb
Y5PcsiDlW6vNMuOaKGJ2AwK/hAdFgzxkqPoU26ZdOCagZCzt9YsV53/3oue2lCRP1rnkTAKxsinQ
b9QRLZutgDIuSWQKi+2iDNhItdtHBfyy/x7nexA/r3GDboGvnrRAk1WTpD6M2DIM5dhQAHwQCBH/
cHiVx4bvFxdx6G0eZjbG9q8ITcuCvboHSqcweWk57OQQrfrc7Z9MrhMtzAkQrhR19Ji2Fk4HOS1Q
4+rZsXZX48xfrro8DWETLMEn7kItofSP8wjC0cOPSJ7aDvA0DyY4kO/OPWJhOAgkxtz7CXpYbfOi
Uk+/sxMih7KWAuS2xBTzLXxCHyXz9ter3dMI/lwYKKBqPD35gKllS0VzefJIvLHPSOsTcXnTzpd7
BOuWxubSUltBj4mORXCI1pnrtFTLKmc95mL4k24fcCjYt5HqmZgI6ZOINj90P7TzM5B2b9U/VkND
1iPb/F51Lu8WBfxpiuEcCb3WXgPMctvsF/gcd4VV+QCU7Flh7qK350oZhzXsi8DlL6vvYon/MKNQ
lU9Nt0lUUCWKhUXVSF7MsZ4nZR/oRFg6EN28vbVQBbVFTEBy99rz3iCukLWXyQ/EfZzZ/Mms1A8H
aU/ATJ6Vl/nJAzjKd4jXukOK5guCjgBkvfzK16sNFkTYuiTgYB/8+GgzC58Uu/04rGDlsPdaU/WE
R19vv8KOSnyNCdVgK4hQGGRVln6MVjzv1wwCgyXVUOPSXBnST9BXjPoKClhkgFyuMQI93k1/Xi4h
Xs+b3cWu5Uo8VGLmnkdewEPPh59A28ic7aM+uI1jImDXFMQAkcczsrlA5EIl1GOm22VL2wjtWoTO
Rg5K41yKpGmjtW/vFZlIrMuOfxyB5vZs/YzYplmFKX+PelbUT0n0F3/2InPQXRTZlxsehC/0pziQ
mKOciE8njlMd4MlL2xF6bbiLvS+I8FT2+coCrUX8GtmtpTv7fOp2TGyfcK9DX9ZznxgDVmaEYjzU
qYDgfE71wRj7GSRy0gh0Kuh1Hr1PwRwrJpFf0bU3+114u7g8xxMZTzE+MAgX6FoewJisgz2LM/6+
eajodT1h9ZAFa3Oj155DC2AcHaLot2ytNVTQk5/kKFActbfD2pCm7aZnqmB4n93i0ETYXUSHsmhh
gpu7tuBA58BEwgaPDlqibPTqC/yuBYzotzvAy35SZUSx4HNNPG0czteioyUN+p4J8QQQtBcJFYsl
jTCkaejKA7odBiCrH3y61SKzO0OBf6/8/Dh+QnzPnYE9C4z5ZEibH8BHGoyngdn27l5pqcTA7b9y
MPTYsuOHlsJ7wKTeK3KMWVcuIcjDWsTQc6968l37W8doDD71vf9IEcleBnx8rH6V7/CCCWX7hWBU
+YTIs7p6JTyAJWrz6v8cpXnONlcKcQFR8NhHQTCBeQpI2wifEbB/kq1ZahXtV37t9mRyXLN2CIbG
5J7eGVtM5PdbfVU2+8b4fUKnq2J19/GxlBTI1Vh4CJwiwQtkDDyKgicR+/XJOs0xrviK6oD4XKYw
VY/mW4IUtflQfPpvzIViMhJlieOeIpUDpUfLgAmzlWKI9DdZ8HSLRRj3SbxscLFVLQANtloywHnf
2whj206ii5b8tEQLUN8vzd6Oh7NTwTZXZ6GN+0kpUfvWPfmwHq1IkmUmitgTUmPh4SjuWmNzkK8B
5KQ9pYdFAxOpCkMlS//JQ9hdAQVexn139N3+3RiYfGPXPeO2eZTCQkaBuyI2KjD7Zk/zUoSB53qq
JLgBMvciLYnajZjWVmet3Z0FoMeGSz30sOnGqx+cl98rD7HUkQcLZgy1a6rm2mhmjaz9q2XNrrxC
jXHnjmUi52T6diZSjDuuxPQWXSbDn9fX0eY6bNfx4Gkmq+149SFD1soYMXFrgd23eDJqavA2c+SG
Z33box2bfhc1dJVrktwRMD2YhqKf880z795ZvQ7ckGmQ0azdO3mPxZtsgpRsFy6ImKaFv1w9+fFE
+PjF2noZw6IRnm+LY3ZTACSvhouJ5ttfJPC4iylbUfu4umVJzAwLbAM58U0uuV8qYsThqmemryXT
jHsOFejyd9FXdqiKquXYCY36Ys9X/u7NiqlKpoU8x8NO8lhvEZ5AQON2Eqxpr8s72BD7e/lugd6P
RYJZ1Q8Fj3X0ZYCc9xm8B8ZPk/mkF+NLxLDmN+3U2NOeaYYP7Lr9y+3UwebUSlOVmRcha/J23Wir
Cx2+bRm2jY9TofWgTRUw1jj71yS9B3KfMO1yWEhDoYUpnaLmV/przxIghVLF3ORMBOfJPHC8wY52
a8cLoDWR+La79rDU0lvDQM+a97QGN063/aQxke8zw9HToN/T8gIyZ+22M69vhzlN92n6netVnsYg
lYPDGkAqu2etjlUuwYyHSF0zq4MZeYaRRlMoqEUtMQwrYo0rFsmXjFMjtc/QQX4JHwSl7b6kaPVr
WqfSib2zZ/kPFzvDBf0ET2ktbjhsmy54fUPtwKPaqBonXf2hehvu1EOvqHhAF0jRjFfXz7LSJXeo
g6oOitv64z+KCYUNhDk/YHEp+/P6NcAi8SUg04N22Z2iBYKNwmuuFJEtv/53w0hpME9n3KXFnLPL
kT8/clvi8V7SVhqfkdhqOgV+CpCAg4TdTKNbgs+54I5fceTUDYa/oBlusZ9dFpsHehFNNbMBLQhP
rPNX80IdAO93Lx2DLtAeMJOColm8A9GhIFgzkdmTkZm2gVkVJaYMdD3IG0maqup1OW7XSOROCztc
oxuc96RKpiSa+Ue6R3gxXOHl5U0L8ej8x9dfDY1W5hS73WJ/5wGa2waNXLp6eL5rQiD89SbVMdj4
NPEca1L0jUHTDOf9zQH3DbmSIxb7NlMytHOe1ebYz8us8ru+D0UmRCwh8LRPDNCP6wAmMQz0UdPZ
Z66ilGnQCnf0zQI0Y5mz+j889xbPkX0XoG+EouXXu/2vgkwWaHvMEOQQcrSyJRCSgqdMdsyUGSok
pRyEfvhJzHGyvyfnY1BaYPAngmjniDh8Pl3bbU8rZ6TkGKEdpbrgiAAZm/ggbpeVM/VY0RC31Gu9
0pi2DTa/2cYeuqSn4dMC3UA/t6tG8SFy36JZMelkhqId45z7Jta6oOGvxxoaPyxEJuXU01unVjmk
krt7PKn/ktneUqkfTjEapNGeH4ebzyzHv4TRYGHsGH4tmwXs0/MtFz27EELxs8/tfKhqdnxhPQg5
0tQ/q8CO1VPAHefrFh3XvIwy2ky4vqu1UN2azx0CrKJb5R+MrR2QPBg78PRRGe103gf5bGSJQLmn
Ggg/T4GhvjIqSrSQWlRJ+BVIF4C9vC9r/PIuCm6m93K6Jn1bI/VVAECnvEsQCeY2upchMDIHC12W
rd+6gPzCmWJiCcFzpvKuhUa2RLglXvWjyL7r6sdfRyy/8AVkh1xI6widnFSFf7Eit1evOPMkwAoR
bzkGOG7h1b/Fpnk4oRPdZBHg5+lMGQW/CnqExSorFAcoCJdVJLFM7A56UDkA4kDvTmwCjbpHUQ6c
CtJVrkokXJRb8i/n81hygJEIc2o5/xu5qEkOEkIoaS+uy42iIRHu358UYldHkWMJkfgciWujSG21
lZCZUh45HHXb1IxiBETk+wPAPAu02xdkIvrwHWoTI01gUOQRscjp7szRMyTLeQbUbBGWKaRwwAXX
HJ/96LHMjAiNmZLgeRynaszSZE6iECiUz/IKc+APjNFvqb6ABeT2Bu6KuEi3NBfGaw6lSdw/B6Pu
O4mOW4k/Uzq3xwAnuu5yJKE5puTStgOUMs7QJIKmW6qnpDb66qMPIohSzvaXuI+QHhav44TZ7k/T
9Z1EcWysWaHawDsnLfBY8E1DFJlMho3HytwIN4eeNOge/on8e1nX6vcQ5L/cLQv3vgdvMA6NCvsn
ay+u/tJc5N1ez1jgvqjtnkB9kcMWX7k3s4cQWSnQl+Bl2OuLPTGbprl5+eHC7Ys8JYQcxrXrnCsm
aEjP1YJXbcD3O135oWtDXsBThKN8OJtHg3Vcjm6YeWwvXJEQkhlXmgWFdfFGSAA61UBBhfj8zmUr
IMlCellKdCAIT/ZzY8hDqvZOzCqWO3DxXGhQAzws5LlXX5Jp2jdKM8ePgfRsj3J+gbUmPCqLesoU
eUCDBFl4x2DqJt2An9BI13ZZ7YiUEOTxKBVfIcTsmVm3/XIIGMviYtVWSHPRGAvZ3b2CyFOtrgKd
5JEYM0lKt4Tvzu/blZWNaEtcuYLtOUf4EJgmb9jYXjdV1iYnIRL8AM0UjJ9VRL8pnFbIbjnbnhxD
THLh9SYrRd+t2yce9icbgQwl2cEHq1akoiNSsPcfhTIHer65jW5LL6MHlWyse9a0h2cSB/EAKYal
Oqq1XjtCH7uSWhiequ3Q/lf4WnB4KZPQJR9YFfeuXeStcyXlFa1ANAWNWB+ht5SDF9QMoVzrvNqE
6Of5hhtJhkUWGSo8NXl+vVeXfS5FpJm8vpnFWJVXjdTJ4nLaqP9Yx///y1C6EgwwRMwLCm4XES8r
WuhE6cZUK1aqHSgaU3jyZZfStZG5NbcB9tDwuHANkZyrsn39vuMRTvlBSn9+sBJd8zJKCE2sve4s
TVRdDrBmo1Bugs4vzZw51JR4UMXy/QqMveDEO93e1uHJShIA06sfwcHHW+T1mMXJt3DWVk4WmUqq
pAYd0zzjpJENc9R50aVcQ+5NIqEWaIs8obwdrk8otvKZfskIgai6LrsC3JBvu7/I36A8EEA7eFzX
aS5/aOrjP3hTwpSoa0uhCer3RgCQX1PmU3qvN9NWbjXCq6b6CMUpb6AQDV37e2E0NNkvQIKO6u6D
oZ7iJ/dkjzM1eZUYL+uQXCZN9w9oxz3pEobzsSTALI00Qodhf+rkyvH7Bpm411SuclIgBDwsGOA+
L1I/7ey9uCQhYUu8Zo02ELA9Rx7A9F436uIrLHuLdoNDuStKG8rK2GEYaHlIgip00mqBS9l5+KEF
JvrhhmnnkaUgTc03ofe19hdDN/8jaqrn+NUIwbaU1CtrZzOvpQB394PRvAhPZWCDXFFSld7s+Ju6
AoZyP5hkPQoBJeCIhgX2ClLBSwv/WK6UDXqL9s97aMaoKTvGPinAkLhHBLhjxe8JkEDNPM6RORTZ
y2X0M9wIW1kt0SQkd15EbflRJdqGI4VTqk2V89DgPNnjoKY0cca2K1ipYE1X4nLk+rbtxIRpsCWh
a0hRz59XtiV/Yc8D/Q/uonYvp3hjjF+1mSc5Br0gGt8NEQO09zh79dUEbZ5mqf1Us40HL9hp6I/R
Wnnn6Mrvb+eLCt+J9+CU+w8KrpManIEVjODbI0VQrHIvw7SU5JLM3qhaqqvahquYUTi6VYXSZfuQ
+145X092OZP2zTZM6hXUdVOTT8EJfzm6n6XB9b9bAJXqlw1u+FHSraYVS4b9lXwSi+wZavhJoXmX
dGyeH2JfTpJeQ3l0KRKVoAIsMqOthEeJBrN8mTqW4AqL2L38t6fSBHPeyYEtAGWrCyftDTHzgyKh
ue2DUGAXEB0xmDIlDYEpxpExDufVu1sDSx10tCPEpLy1rkdWiCWthKvhfuKH8gg65MLf1wQWDXiy
gKtw7eRP0rZEaonM43Xq01d1DBgah6ZebP5kGgp33CeAqS3YdFZKvVbB2V8g47U/LPv5KPBWCMpZ
EQE+MPNctFdRyN7IR+HSIrflZl3ef9u8lnuSVBun0U74LCi7xZ7geLwKSnjBTldTz8hm7nNnTtBO
vaJo5+Gn3+w83AY5F9168xmobqfAKzXkt5v67Fk4f9KxoKR/QqlV0q1RtOklzE1L84VCzyPbimOl
+ReaxEyG45ICjsYe4RLSsJ7/6hybTxQT5oTQ1T2qSok7v5g/f2a/wplUGoCsoRGazg6PEjHsXWNQ
gRKVxfgVg/DAeSvxFzQ5KM+PP/oOVh5yGA76DOmEUbimnq3mno5k7TRIm3bhZPukOK35aXmcyNwp
3HTRHNWHqff7eeZ+Fg96S8ZottQIIUOdi42FTWb+XlH/60kolL2ESSDjFz3EH9brTHiUCfxlXKqW
vSRapGdS72lzRejJyCz/GMFloWn85QV1b80YysoQTDoPGdNfBlX7hpsG4A067A4vDN7yjZUWpwSd
UjPy6uGfAAdfg7mxnsEiD1B+dPKzhNDLY53as93328C/BeaqTblwB/6YdiG4GXA0JQLK8p8Jn8Fw
cQU1U8zipuI9MpEUe9zZXh9XJCwVfwleHluZPz2Jrrj6M0G2Rq0g5Md2CcXTaOICs7zK0yktpaAz
VgHHAV7SC86Cwi/6CYo9Ew6FX9YLU0lrewETBCyc/N/TNX3uxVOhyGrWIrypAVTY3La6H+1f0BFJ
D49OYOe3yly/jW9qoS1upYSoUXuDspvUylWJfNnN3s2SSul9pwLEmM/o53Exus3ktuzI1JZND9PF
4ZESmeLEyZ6hMHbF7KMvp9eqhSD070G5sFZRIh2Ydha+sPxH7zh4GIWcNEqs7aneickD5Z/CUtXP
L49JGRv8gqW3IeqE4CVljhQSXuGbRF34+GG4o+ipM4lT+t8dr8W5mysyOzXFG+FHN9SqlfTXSN4w
gTdJgMEWZGVeErcLG87HOuyLz1Lt/MEK6lIbxp3vTYUr/OHxWniYfKcETYw/NzcPtfdvvL2yo+dz
Hj2GknGhfBz0PNk7FBb05MLBtjUuWpNv+d3gu5BHKhaeo42aZ0+uda3R7owf7maIg8C7ywuj1Nt3
MNv41hsCvrlS6pfwVI1GRWuZjLoKDQX5dkBBDlVKAXG6vlu7HbjJoFFrOvdgQ+twV2nk2l3YzQCJ
gs7+FM5MXpnLuJWbbxLxM5jOY3yxO5v1OeUFBZCr++W2QlXd1iUIIY6PajTQkYUwd4bT9Dr7Mn1u
qW10r9lHIOV0UAba2kOSrKMtqzeWw6ObpCSfK0HAwaljHhxVwC0ZnwgEzBCK4ETFBsOpy8QL9qgT
9QV05b+ex9nfMgiB2dPNLgnSW5hINUMzKvGMAk3fF8NahhbZ9uFRswCfaF5sVd1/uqsJI3o9WbSd
PoDvLo6pDfEtsbRaus2O0cEfhfjnYkQjoSbWF/0kreV1vLXQ5r5P1PMscJb/ZcSXlv87WP/GV0ZM
JebXbN+j7OAsXS4/Bs96tv82Qm+749aIFtDB9yaX1ZlQrfUnpU0cErzvQ/iiwWWu6la3H3F61MS9
aJrpFkTsQbNbEU0CgzI6WnlEnMrhlD/Pb/CbgL61cxkj5G7GNEp6EI2honCq9AvYPBkuidkT23JV
dcp//bN5/TdX/HiWszdXz9kS8V6D4UEn/M97y9nmUkN2KcVUP1pEZUyQlvn3oX0qGgVzk0Qt6F5G
hNFGDysbEgpneDlrKTHIC8TqYk2r7fyxw0oDHs8dpycl8+CyOUl/5//Unyi6yS7Ptezvrt6XxopT
Wk1kbAzUAJ5OlkYQRpWoQxFFhjZUBXCBy6X2UvKkJw8N5kAeOsXZXzjDnBTd1CZ/n3xdUSPLOW3F
8MqzR6ce1H97r/TtF/32Mr3ynjTwLJjOdVhW7eBzdJFpfli/JY52YhHs/k3QijL4G6zj6cv0jCrK
NUS0P1Vn31+RogLuKSOdMZd+cfAxso7tBcMq+8Mm1sP1jebvhebC4vAClkA+q1aTrd+2LBv5WyKe
RFwZZa+0XRmfdYxx06WvVBtgsSPZtKR/YwISRpMcSIauT6KQ6w1zt3ZESg2G9Ee9SqZxi/Az7fI0
+Av4VzMVHHX447khVTJk2lIDBOZex5FGD6KJrYbxXLJjcnTablkBwqtRpTUP9R+bjjjGYamwuJlV
FE7RGXe0mAFuajn7DqjmSTsFR8K3eDGDIpDqAiod/wrDpjdOl1IBj7s9qbIlCAeFRO8TcaQVK68X
bM6BVt1XkYnNgEkyuuKmn1DMymyf7ec9xY3+bDY9RySb7CFYM5QynSiak2xVOxKp2nBLJZ/RkSYE
WtNAAtYOyfXpu+lwL6GO0czPCIw5KRRztzE3B+E1xhZAlSGp+qwWvBYwCl10jOt863K7r5dYgt/h
3u0sU5TnED82PPKV9BM+ZsLHa7sVPM8Gy9hGKqY6luv5p01V3oLqdtMYJ2Nw9vSAKfrusG+qJEQa
T3L2KvJ2VRwCu2GhtjKK2GjjQa2Nr28bhcDfj33+Mtf8P8KEztq6REb7PbmqvFJvhz/zuTywHwgk
F+QD38kOVRe8p74wxmLUSnLa/xfrnuIcYKgKuYGqzU7jUloZmz5oMTkZePib/F3G2Ju8Y3NRemhu
nWI9Nc+OmJRgsjrxKudc6Gj+bUvvmMQXySDTgk9VgJgBvxmF7Q7aUHFgFGcDlfVM1ePm7nXEvsGg
hHFObyU2DYtdjNWr5ogNslsHsuyLK4hRAIS2fv2uQJ6mFwvJEyHupXflTDeVaHTNLDggSiQsRKJA
dNjcMIIsKoQsIhNAfDeKPWUp0EQRmQDY5ZSq0LtdHh4Jm1Gr6yFrT4WolZ8rekhlq5SwSDwsON7T
yt1qeKBi5kJo/1M3fkJjAIUoBJBdDf8MePzrQaIPPHsG1S2rWPseTn2rC0oRSdtu0jBNRFeW5WeE
qVyOeF2QihAW6G2esmII8LQRfGevwb3EqWGpqO78Y8KBgjv2i7jeOyBnJtKZF78GgyAm3tdUItO/
erQV45A00RMCKm9eGbFmoxaIb/UscRs2Ys6LuHknXcp8hp9B+u9I5mMhObNg+2GVchmQB+ZhDMug
g9QwbAuEaqjyoNAeM5GHj5l/xBCoLpMig1811hNFgxAWMuspmBp28vTpmYVZpWpAgggeU685gjGk
6/74yCBKbZordzA6MARCIpu8FDMjiaJ/dk/NVFXZQDUhpMs8+6WSjr9VEiGhjoXFeWv5LAVv8//1
9a7ES3kfrlijoD577IrZfX4Aj/5jU/PTGptvqvR0PZxPx37EZpDHRdhCisBGIRxdxT3+CBqopgE4
yVZv7kNAjBPNTmL/0kzHSYQ8patnFUNCbxGj5WZgJRm2lhIbwHWsFJilBMkbUK9aeKLyJFqKccVO
MmBgLXweyPrWv1Ru7dqJIS+VyWneYFaDt20lZa+fJVDF2egvJK9LnF24Xg6m24zxbRjhUnpzjbcg
OC0R5EqtESN8VXnnqWoKbLm0EoIE5izhHVZvgmmifGnWnnaK70/YKvp/RHrJZG/OKiPasLw0RtNC
5dxug0cOmopcGoosm1pDeAWM+t2YM4spwGjK5tWsspAIMJUfco3Zk3gr/V42tMubr3FddbWf3LfS
ezFZqMuNYzfRb4DcefLVJOTtYoWheYtTiER1w+bTJ90fGhd+Y+m9LBOieq2zVd7O7etZ+lqJM48T
F44CifkStjJxpTNbx4x599GgyqDGJx9ycUHPhoewdiPG2P3kQMUklYyXonBVXoZFkZCcxV4DEcCG
wznBxRNLR59Nz1dMrveCFN/9jtCfsqDLQcduh3Y/RMPA2BiYMIT5ukPyPXyI9uEMM1oZhlvOVjD+
miWgltfDVWLdrZwR6Z5FmIXTtbPwxBBuPH6JXEOCx1MHEYOxe7IMCVL1oemJi4EPGlszVUSnladT
CdT4cJ3RLXL5hTJXgI5ecRGYMIssT3WheAYMR5xtNERPEQCuRK9nhXINXa1xal1AAygBppsj66+3
GBQNbakqmy6thPJMiGheAZ8ZFsbY/yf5hGf/xQA2Vl17HpV4+cisJChmWq72W+zXTNagM9r7hOqT
7+I7EHqNbWLWrdBdsMPR3cbNPCqjeuq1UhF1Eiu8Ia/fIPwQyTx5+KBgteZA1gLliMEhtm6hCzyX
fqVm/qLXH0mW4NDCh7D2ztYRD7aCBcio0Lgz3QYhqxC1CvDiWLy07gUdOZlmDvaNfve2qAw95tGN
63b4ErJqHRd3C7FGuntNNyIh2Wws2c9rm0F2gQFbE6pbckK1ju2btTRqcuIOh1pxcmj/xRL6DbqU
Z5NaVsz3oqGuRii3REMQ3aoEYD9jfXk+yq1flnIL3KWshztuivwQ+MIisSio3KW7Crm37Ema9cb2
TjKbO7QH2wRoXTPo9HGVvWbNKH/nfmjqfmb2w9TZB5qxg6BI0JuAsjNvC6Qp13a7TwrDEVjG7gp5
aCc6F1tju/5qgXNdD3WRLw9g9rKg8zUy+tW8/hzMr0/+D1hnjGDU8RxeopFWvQUuIqsbB+FDgisW
6SSyGQJV9LOJPBw55ghKRhHG0MYFXJ+Kb8y5ZPlk/NA1Sb3oi1F8YbCXii4XrBa67ZB9MJNqmM9P
xMeJr3lIxP49X5HHtVP5m30ZpitwhmXoA40rT4FtRioLeYSVVpSSAGjFl/+6P0Zy7u3pupogRyHy
kyiIuZ158irvAuzsiqsA4G/yTQuo7q1x7QnNWFRN3JAzek2DvD4m7gc/q95k/ZADrputX7D5wLx/
qO04e9DwxvDaS9U9QSVjix/+77pSRrPxGWE2xygON7dkmbDTmXbJkSRFIvi2h3JEF5X/TZOLqeQk
ZhEMn10YumL97zf3tIIR01W0upd1WOLwkHmx/1tGiplNHhTMVTuCDC4J3iA4TXLNZ9Y194eTsVFL
zsqD2qNBAhVkc/S86aIMCCqI5H3eS01nt68O3hYWDq3NyqgAhGH3u6RNsw8HhbOG+sFRMPytpIW1
ES0SslK9W48XGXzG0PoQm1k3QJrsUGSMrcHJiAAYy+INq/ghUBUX8I9PYDko9zDgR6TPR68d7RxR
eyx7EHWEnDj+ZcQH4bXHTC1QDl2eItlubP6uGWv7+LFWqIfa+PHhv47k/cadXcjHL0E1kDHCwKC0
8L42kQA29A5SRatL03s7MShrMjK5nP0UjR2SFl2kd5U5Sgci2FCfkGRdtsTpbQ06Hjshx0GSYa9s
Oy6FkdNWRfLS49rDI/A9LqyrDKRAlr1kSZ1w5ySMfoMzYDm38W2KXD/OL+29nvnGxsVwKxaZr2SA
2ugCb5hcnEVqvv01iNJkkOz7XSJYhOvsiWRtqpTuTGTHlflUII11sjZ2zdlc3qPBlt/c03IKFdIT
GuybQzvW9WTO20LGrCg9h/ZZYFH75L8nB9mE8Km85pqJe5EhRl+8z4ISkInOm0kg4AwM8SgST+nF
P9MMsJAhs6WJ7MsiFB17S6zoUa32QzJsArtvPrjXPxe2I699GiKMak6w02z8ULGhtj6gLCCvSLYV
Q5HgXjdZuPElFnJLInHVVzMpOBuuXF6Zxt8Lmgb91q4AJrSJviE3OHNNLZ0flbnckG93SYEH130s
EUH03kAbucfAlqmGMezJTbTYQjU7I97Pd/hC10NPinFnfk/ILKUyjtWrMSdsH13cXu7nptv4BrWP
XnHD+8olvEYn8maWtykRoT5o7X2UgBAU+P11AD16e/FZOdWvvh6o+HxgFlZqaLGc12ItkLzIFz8x
h/JgCMJo0kEBvhpMQMK2HDOgYdgWm4ZBIvMun5omZcwHevRQr0xrySfShj9C634iB57uK6zVvuEC
W/eOElmSjFqKKE2BiIiNV2kg6KX31rvOFDSsGox9bsBnvK4h5Yfasm1aqsPJ0vf8qo0acCQfty3O
Re0aR5BHrvGFaC6nlJmdAdoH/znIykjg+EoOvgNqkVEKgui4uNIzafbl+31eOyEA5J2QZXaxXmv7
J0+D7ZSsBOwq85RRbS/GmoSdTgNBoYDFqd1ejSY7C1PPPzu8LTxdLK9YR1kUy5R4xPZdg1pVd58c
66cQ2OZzaHag6CcI22/gMmQB6/eYX+gt/wHoa1WMnErFirtzy+TN3MzksElEL38eDyCB0GNNLXKk
eFFbFdp/n7MmfWKBGjI0TekPszS3ef+lRYdGU6ROPZTAOuhfZ1iF0SFNd39vnop2GSegrnBA1CIc
ID8HgFy1UnL97SBCZa293TiSbxaroMMgxctrTfMXUNDtskgp2FPTKIBKrVmAv0Ki12nHJAM8RFxh
kDG0zdHqFZ6zXfeUQ59QYCIDVsnRkNNlU4LveQI9wFxGA43B/XKNgFI6rWrh7KoGD7CCZ8R7Ug2m
IxT+u3ShFjecWkLdRdSo/WGyDRlBKM3sciK7DnUDxiSbo6nzyCIw31xxZj2XpfGyAPG8Z/V4B9aX
D/tjyXc7TFeke1wbpEr4wBhDJ240j7Eu9j9NTUaBAeEzLHzx8/Ah1wjA5sZKmfiE4sevmhBB6vCA
laR+Tl5Zoj5HTX05wsTvw9MAh9FMDmbOrZlQaKqPlhIHNqFZH7ybF/ashgDl5sP6MGwKm9zVkBKt
UFtNh55gxLU/q6MWDEKXCAlfiJJGEUyOQHePEi3py8/5Qn4Qd4XdrcKckplUrk6ecIZ7jSp/+HoD
5e8majMyCnh1HthV+09WgpEZk/E1pfXtlkkmkuM4ROG/ZGZAOiM18Lb4lFBc8Ki8nGsgJZjIAtkk
hJBTYSInKO0n5oPVStJ53U6bh7sS0Q2TWgjfKgj15c2Gbr0lGqFKJvvRmKUnwp899or0+r/h5zHS
gef2lmoIovHt1f+SL1Ear0Xpynbbt/E2ojz9dxqjsXT7L0kGJk6EPzG1xWgXrxKd+z8CgJGogSJ0
xoJ9jv7uVTT6lndBUD1WjvIDeKnZRf1ai0peI2lpceSE+QWVNq54Nttuv1tZ+zTZ9o6bSNRyq4/u
wiokVkIBo22mMjs8re8AifIvtLPAvt7obv6KORyC9nnOlHjeSfeqnQvhOHpCw6MKCtvR+nHJtYOZ
xTxGfakXmbPgBqY5QcpjHXWqomoyjOEhrmt9NH5Vwwnk7+IHEei23ynNuG7fvY50avoZRKCBS5+Z
VtAIKIEX5KU2nk8PRe1K+Ae0We+h+bofiwYVO8b5uhlq9zdlgEE3svwsLzWVdGiMfPy5Tn7mh/mi
eYcfmY6cBljJnFayMAzCKUrcD+YD1HjSi1faxHezKJC7zgPU8zbpx8XIGLRh3ZZd2q/Qv9LKIQ8M
ulKThM7kwomKsiWBKzo+UUM7yH4rVHqyI1spwlxt4iUYN7ZbNVvV6+hWZ/dhhyGhIQJS2vBPOxV/
ArjHVIY6Sz0gpc78UWk7vGqkW8YuTEcyM56EtbJZcBu8VvdkHSsz7oXhS8z5510Uym1AbuU9Y8G6
X6SdNvfHAuFCps/JgYSSyTy0m5+wjKl1aNKW2UOuM3j4T2fnwyJPIQdWgZ34u1rG5v2HUillQila
SVptxGyLfcRj8VnS6TKu9FqSjuVnE+rTzCRUj3UYLD+6e7VBGxe3DKv5149x9sJ+zhNDa+dpQmKV
gI+zIzaWWPvYT51N8mpXIYrY02W+Qlo3NCZkI9l5+un7rXONgQrkXkFjFsOdsXTvT5Q7sg93XVbv
ussS/NdHr2STBEZL/HL1K9zVvXDCx4Druj9nDjQerUv/5WdkXXxw+y+iW8zPw+nHk+owkKP8Dt30
4fag6h9pPCx71N9n2f7E3npqiKXnhrt8n6BXjEYVzNkYKOSnr27+YZFPd+i00kt401X8+5QplZIB
DPLxKlPWbpor0Vtc/mXj+WsZe/wrerdavmjZKqpfV169nAMj10l4slRYIPkAY6khEe1UWyhu7sob
9eZvwy1a21rMGyunGgIQih/ZaHsZUw72UE4CNF94BmYsB0BtkUIfsqd1h7DdbOTiAcKkMYTclFas
0lvvQ9WNxjLjm566I5hdIq3GFDvRkvUvahT4KYaIf/Epnm81YgJxL5nKdI2iqjLW21PCHOErXN3G
dNr4FRNTxFUonFnkCNd5vPEcnWddzkcBc0roRzfjQ2WmHLvPA/p44tgq/BpsY9sMOdd5HxbHc/az
Uy7vo+RV0ZBmT0gfzwpoTWcK9z+aRy3TuF4mOcjDQspTNaxo67ItP9kesb4T7S6z1SpG4/kZ4sWF
a75nmJIyNPJodqvG6J0iQX6S+IQ/qaoHIOG244PwZ6pwHakCKRc/2Cdx70iyf7fwXkbq/IuTBybg
5OvMcFEHkNESKtJIqzeDpi+KHOVp8gGo3yOUTBk696iPTI0LOG7XqRbRzYuo10j4GDWWigkaCuH9
sjWod0A/m1Nv2qrc9nzpteRxWT5ACaAb5YOfGCLq/X7b/OY4DmvXzeKHSCzUty2VTqziUqpYL3kO
1Yd2ZHN7PvDc97u5kQRcMlrPcTdtAdZ6JsaudU2yDp4w2EsTUIE8g8I8GyMgRhB7oXENEqACx2TB
OYtjU50aITpKn/wMKPIFIukQJwGIaPI5HpYyU9gu1PNZgvb1h/mjDSU2aaxGrec+9lhSjqXv9i0h
3RhYXGVGXthOnLhZTbTe2cb2+gZKIvhlMkKQsL9OKXyvoVMC3DUVguOM0PGSDQkZSFsZwYx9vwKi
yH+eIpM9B5+a3xbM5IU7dacorW6bZlHAw5uDM/zDG79CFy29kzohR1CSzw3rrT7tax4K7tLJf6Xp
/sYdd6SLwwmqjf0juE3XQntU8nrsKvm/dyztRuypvYyDh+WLhQYhA+SSRdp7RprBX0m58M9mCa/t
AXb80hZ4oOXEwX1E3yc7iQrG1LzNbsEuRjVal9Lq/G1oqimHk4hRXktCp9xhTqZbc3QHeEnDJDw0
VFE2QNv0+bi+HFZpcTIrtQQkU8gHX+cFDJwr1X9/tYE/sQTBhnvE5Z9CKo1KcAPj8iWr+CGqqy0J
dfhKPOz0kuUN3PwoY0eZDNsmCH8o1fVrc0v//lXVUhYCS05jgmKdhpwba68dvvHxClwmU7MHhw8+
9CmID4+V7o5I7bPaeaCF0RbJFHT+PYqJeiscqYPk+BjhCHYMzTajD/3f2H64b0jOQTJbF5yfohRN
poappyeBBWqbuUJK5dz3elVSeLTIQg5NjihyE7oQzG3fmu/oIaGUNiVBEuMki/ulg48K3EXZ2Ru0
GguVC9RRoGVCRWo1z2NzYpismuzgtWQW1+cijgFr2RWIDW9kWkecn4f1uHflKnM67Dml9t0WfN4C
+6D4EiPoIkvXNDRUOyNhhNLSHzQue0rB1IA+CCwvXSAPlDhIWV2Wl3OOujIYqsBsDONqVrjZWKZ+
QA/XH4xAcz1BEcmhs7Qf21o7ZOzva2cotBXr1wzuFEXDHLZqxt/qIYQWFu1uFzfmko51JQ0++9he
5OgCSyqWGmfdLtP1oCAUxEneW643fhsjlobeKJywrIa1F4YEb64zXhONJpy83VyzsY6u6L5woXAL
DCnqr1jY4L7dtektlEmKjuXWYLWK5gbWrvKmJKP19d4IPFJmW1KgTU26jkzJPSaByr1B7dZKADKC
iv3zC5x4up072ozbVqWR0iXE+tJhoiqFAaiIi++6wvxUTsIdb8NUkAFypwTo6KjmoMs0QboaTfVv
3npqyV4JsaOcGSwMD6kvSyYoST8vd5O04YRHtyd/ew1NfV2JRNJlzOBenyYED3/QqJ0/PNjh9y+b
YVvVm3QTNgVQRHMO4Hg8CwXyM/jS/YE18Rt2E8ZOiaKnCcSLEGEevQTb9gzak6YtqhNkl5gcc5MW
PvBp5v4fjX4cO/p6bl5WMnN6DLlqojmM4gkWPOIF2W5c5wiZuO2Lu2HBcoV/v3rM+B6uCgjK1bBl
9Efo7LntzhrZqEhRfsxw+3RF0tWDwVKKW5wJwfO8bxqoP9FbQFiz4URi3EuX0Pa+6rE5TrpcVKRl
jGGEDQS4Hq00WU4CU8Sd9tVXcTzhTLM0Xd1jkw8WTgwYzi1GG8Fbyin8/TXJkATdH0VARe3Bat0r
wqV+5UMJMeA01nt6SvubGZuJsNs0XHBMwrtmMWtyXFOnRHkgIsJi3VP0EMoRX2ExONlCAZOsMsFm
zynmLYBdHeDWZQjNbfLnfb3KCPZ+gNz1EoNHrlPGBpTOsrUzjMCvNzIbgSIRJwr/QCVBppQk/H3R
TYZcGMs5SL6Fa39GbwfU9czCzKCUcDtusl2VQBbI2b7cBNSdUUxDoDzrmucBEhHvDoCId+w2H4jM
T6dXtNVizpBL0zywRQFlrIHeSr9v/Wvp9udb9jy+XULJnw6/UUhLgoFyapO6bdAAPP8CWyYFRQU/
+5uOUbhwPIMLplUM0ACPDE7jlhUWIoO4begJGaTrmYOItnoSANkZBAkKTuVL7eciQtbPD8etGi2G
cEcurX1QdjhWhsnxjvhCg8G3GzL6qjfqmpAVJowqGxY1UpQstHdJ6DzkZnASoKRmXn+RduoYCixE
Xj+QdrtrDxnOK1ZasE+/81oFI8mi7OEMyyNTMFcIIaM33BWsN7KphtEHkgWvJUFNr1Yc1XRW/Aic
TtPpb+fzN3O1Tn+o92n80S1RVA03bXsvQnoL6eb3wYO0ZWksbm82QkJgiOTGhGGMWslhCLREWD+7
D/vLonUXaI8KF8ubZxVjulRNp9RD+wVljw14cOgMofKwwHGcEZM7wJBAK3lRabvhxh1ZslJxYXLF
ZpDVk15bb57FM71/zUrTbRDvaWCEtQq97c+T100IjqJBaxjcwqSSZC/irE7vAwj56ts6Gbga3PX+
mA/6XY6fWwmzPaDto203/p1Rbevubl0ml2kRqYKgwtQa7tA81CIESxuqTsngR2+/J5ZnYY3pWmwR
+7+WHbMyGhKbiVHxdVZpql6oupSpc6et62hZkENIirs5607Fmg5CuowpBVjW/Ev1c8L34Dp1FVtC
BvbT5Fk+WFGt5QrS2luqzzgmG2GgtOig3ymdprfo3opDYhlll4Ot10Q+9VRuRdOpZgr9EUXfRJmH
vR7HLqbUDuzgoFbUOx7/wkk9Tkv/5p4SpNtCiIOJbuatppfLZyvkMW0kVDdcQisPpf+/wgXccuFy
RSz+YWqCvqxlcBdAkRFiEzjE2yYxciZQsFaq9NgmVZaJYWrtDjjnK+h4TJJUq/laRa/EXpjmMU8j
4MwL6suYvFe2Cyn06sDOI8Y9StebNJX3TzYie9BaEY1MPMgBIN/bZvI7MooRVnsODp9SbgTlSA6T
/3Kk6QjrYQL91EETVsyqwjV1CGequ7FLHkMyGPZRIRqJYLNkJkfxWH9/QnGXHseFYGoK5VSk00Qs
lUfMRNJKf7y0FksJrhNQKQiMeDmcdStOnm1HT8ltz2+Tw6TfV++XhEmsMhHzWKtrN0tNkFmgUhMh
HWkc+CWUsDMC13wD4Doatx2iJNuAV0Nfj97FqbZFIidvlmLBOywUop5bkWkkw0wEMAsbI3AMYz+q
ohUjXXenl0t4D7yuRO87CjS4++Y/E/0xrN2kA3R8QuX3YeyVPRS426YO/8X5A7nANx9UTkoCBbAF
NPGeqoe4c4ARjDaFhRc94Tv5l4a1LGMG44xLxTBBzNW85keRI0Bq89oUUIjLtIn343imEvlPzKcZ
7kfqL6p3+aNHH8Kova+d2JScfeqt+RRg+l3GQJcut+hI35Ue2O3eDKhn1v+yGhdGFTEGQ74ODwL5
jL56ydAU3yi8rHcqNkHvd4DWxXm2bAAjO+56RgJQScywRmMeuVQRdKYotXgh/+Zojj9QHsZWM7Rj
ak/cdAp6BlsACb0bLxByAOazt7SGnnSMwwu+AF1IN1smp/VtaoMe9HwnDLlyPzswZC/BIYq0IUl8
lj+A6hmY0jnBqktY6b8iypOSYSpK0HDoXOf5a4Y9UJ1TKoxktKOPcTJ2FlafFFRrzgRviMaNk7YQ
ghoXri+CsTGmS75Fj8tgs+ZMQH90vKgDQ8XV7KX8JN+I4tZ0/F6tKbG0g4bIJ73lXT/a6NT3JJkC
X9biX9TPTGFALb3rpz+R1btbbUi+dt/SnsYzzjTPc198TMEGYmQyCB0DMcx03UHK2eCnUYsx4sDs
zsh7PIpxXQyZPFKIi2vuTKBbhopEr2l0RUQDACH5dqOfi9zjRdcLpuOYb73FqctLPXhUBwKiGIBC
bFJWQR3Hddy1PoeeEhGcdY9llkbjX7tXMDIaL7I/chFl8lhsJpn5RhhdH6X9951GuTzJ61BVU3NV
kkgmBgYvw6+zFHH9/rNYNqEu5Bn6Egi/O5XVpMSzokjpVywT/8ebn6Hv8KMtlF1ygSSy7hIGr6tY
/8AUFR0UkDXLrkyk7y4seP3/cxk54Vxdw4mNlZ4+XnXnmdR1HV/wmAJcYPdPBgFrdBsxZNhgFdUy
JYDgVLZ/Fsyig8s7K/Z9NRB9NoskZNFjwSi+tbcvVPlo7Ddigrw/Mpp+HUlbS6fQHNjd5JHJms5D
KUdmk9ePNAyJileSKQQb3RIrK50SsuGXROjz9nLIMQIkJSYdy69kn3/BbraavpFpkzK5QfgbhUI3
wBTx7a+dY8c6kpU+H0zz+PF0J3Ls1FCtd6pwen9ATlBJcVEUxOExhAXDxzTMN85XOLjVnQ71Se0T
QRnSz++K0B8Z+j2DjFx+kQ7MUfjs51UltoAs6g5NkC9WI5bsuqr7iUpW8+PfVtheCTpf2dG9fwb7
c6Kr9NqpvTPF0j/9LE73zRcBv8ID2wyqNXLPpGGxU75AQAK73hZnm7WJ8ES/JzVgJoI+JkZQfG7+
eSiJfe4+xVchZBEtZiFYckSmv+Er292rbBjEBKfzC8gKZJRsjKL7tvUpTuL9x+8zJxPtASzS1FmF
CGLfH9fpfixRue+nOKY4/XsvJCyCskhTEEDaxNdU5GZrs0vOOLGgzg+0QQbkm0fTEGummyMxjfWR
QplRT2NbUbdpcIiU+vewOr1ZQvpciGMmcOFPQmTV9sw34m8reisZmHvmNbp6AVl1Cx/QCcc7Fbbz
OH1cTQoi+EHr0Sf9asoPY3+FPCqdlV2narGHaaCiQqUC91Tz46nERkPYvRSlCSPPO1jBsd/5ojcm
HWSXcgRi/Iq69QcuObRA0hV47uS9wRhDP0itYJYFU5dkngt+OfiM3wvxAeaioKVVufO2IyJ62Yoj
T3T4lCRuyj0rkrE2h1/MLacbw/5cWc243u3n+b2Mn9qJufx5bt7zMVhTHLTxM8QzrVY/JPDIIQ5r
wOxCXZ3zyR9smQ/BJ3rLneBW6/6yE4H7OuGaq7j49v869wnHbaRuoKeMQ5wfBkSAg8oW2WNJ9pHT
DNoF0iN509nEm7O7NnV2/4UWhbDBrIqK5IpK3X6g1RYn6WLJ3k2fuHLwLnj79XU0L74luQFoLaCU
Is9BeUuW+VFdHzolYUtfPGxagisvAVaFfFKNYY1Iq5HIURGf2R2LvILdxC9Zh6gjGE0J6Vy2WafJ
OhkW+9OEeBOuoNEIU1/6vNj8SMwfxpfQMz6ci49rqxsJaLG1QMIQlBVnrVtSpoBvovGYIGyFDGFx
IsWjtiv/3YsJZoryo/TiJ6xg/kb4LA4F3bEVDTxhysbAZyct2VXUJILIyB+Xk6/2n97gLfyhb/dD
gTEHY+p2p7NLnGvSv01NDvAg/RqTsavHyrnKDFdHJbMHdYqO95smjdNlzCmZ04nWizwR9IS84otJ
d2gaInuO96mgWE4aSG3S0e+C4rcpViJlQCXIjPd68jHfss+7nVZCqlcSmggCS1gGjCBOqdlPuNkx
YRUuNCLKJ3fHH/arIqQYNw0uOqXLfCzc3/2AUETIp78Vm2Y5xulURIqgNjBWt8ptvOOa6/DbIXsU
fU61oPLoEF8086mwGTTDLWk/5FDdbxJIBg0DG3tsK0pQIcGyY4NWbVgwEOVBU45p3tVdUJAp6Ysn
Jugoj+PckdFOL2Gi1845P7HpkGFWqXiuEuZJWNxspR5pRpsWpiMxgKvIbbsZ5i6m+mE0/xCuDV1H
/9L4BW5W9uQv/U3ud1Z5j0k2lowxGGVnHlgwrSVJgvZjVQKJBqmO1fLKtMCVwktAdi7PfuuBjB6Q
88wc1r7+c6Lb0ukr7r784PUwpKR5FPgFyqJ/8G3CyTTs+wogPkOxAd5Mdhp2+AhbGZi4HfHR2uv5
xK6oQDpYQtI+wQO0zo2zgWY3p5cbExGHpk3sNFtV3RJtpO3JMjIfmRZ0LX3UC0pIJ3uAns7/Wag0
u+uCT16icu53FzSCkd/541MGblB50kvP9TRQ53+kwekRLZBPsvF9OAMT0e+4Ano9CQQG+ahnT+t8
djlXemwSOQRiNgmNCAuMcpks+wYPE6N1+gBASfbCPodOzfB4lviHZN0ywLatXjf5Z3cmGsaN8v/R
PpwbsAaKiPznRNfNpdDf9I3t33OsJyVNlrtf9v4igL+0TKgY76tD3V4ts36jKePo5hCE6X4KlK/F
mXbXlLcAvYr9thMVrxwqjQhN68JEKa1edpnNDIL2F4UnUfL3/btx8cJ6SC4KexfjXVKKhnm5Fi9B
C0a5YilZ5NBu7AyX3BXn56SluN0p5TmTaTd00qpajp4Q6YLhvoeABVc8wgzgImjSeRaABDvCsbqA
rCluWXIJBud2pC9chLJ03564LsVYvotpJXnypOMyIIRolmteu8/TRX5fhTxyQQPYSjN37h7/mY3J
f3iZ4gDLIZ/ibpd21x/913sTX6dKD+lQHKhpvL9oAGkLX2hwv74r8U/CBEMeFD1Utl2bpiaNLzgx
du5mGje0bGspHpETXfgZTQQBWkSg/ogPnETd+Xm8b3OBsJ357mo22W9DcszCKp2gh9PDuKDtReZW
02KuRD9Ki3f3ytXeQuLKUmCFNjdKeh7fMF4Q3h9lPRYXvtyO0qqErmpJJIqW7uObU8xPB07hY9zz
dNquq46l7zsLhujxIpq6indOM1HJdyIKI2TXyQQDBzav4OeZkMjJgqQDn0pw2QhTATC+B8pRE/mb
OufQOPK1hHmjjTGxN/2sQrOqjMidUxybrW2ioTQXS/4Cg/NeVP4KHn1G4YXHcMjEcvEnf3vy+eMi
WJwMIMJBG7sZdYmBL5qFq4tJZL5EFNsbBS7eNAs2GeuUqaRJ0z59felNbPlzFUMwDRFwK5DyXOOT
cKzdJQ52aX6A1MYs96u08bUbINVrXn0bRiPr0Ilmk/N6+CkExLWnpD7MITAdxUs5thEBDby24aDa
rycfUe5IWCCKe0ocgbvBEBwvo7x/27ySFcXZwbdoQi8QKya1F2vZRr9peUNkXWvq+wk5CCFb+O/L
QrsfVlE5D8UE+RgK5q2t2sILdXD/IkMgJvCXGiacGKo9mcP75jxkPm3x9kI7MIGiQsGUFz0/OW6U
/fjkIAb3my6EV9WNQXNfHUfbhuCYBYt+mUmDfPPK2b8JJvQ3MQa1jnl/lOmcZaG/Ds6bcFC2pYHO
lrrSSDCNkX3+BUFJSSWC3YAhci259830htOGmLxrfLRG9bq/F3Jq9GgAFBqoWOgyzfxL2lQMwh2z
Z7jw6CStKCfux4XHejRGL70DDdBeG+47V3lZuQJXUuL1ZenYa14r9vinc8ADs87nRnxHh7YKKTYm
k5nWyzw3oRax5euYUxLYiNkzaph8bbgBpyVfoqVXEMwvThOLRhl8bTS3KPZi53tCW5vuMntkgAYG
QAPxl1EsT81G7YCjyBhdEurHTTPuK67/lbacLk7Upr7w20bveXAHtzOzyi73BZ//KD3jIvzKos4f
qTUQeuPJ02NVIn6aUKQOJvA8AsEJPlPT5v9n3KuEMnd0wWsz/yb95jrHfAx5aBoyd8sdoWGuNICz
63l/TdDhrbS8T8rxw0KfwWiXCUHlv0Cmktw5ef0AeBjJTF2GVzgDMEkzf+483cwwRanRBcA7Caqh
4aCdHRYWX1iFpOo73HnUMeg1EMN/UlLZ5TLTBCfEPieF7cp+MhBluXqWfxyv2h20lpUwoOdD++kg
bZJqFXIgU31Ta7eMwiTpPzmuaPW3dijlV+mqlJRJXZZwBWM54K1kHxfyeLEbw20WMGOawl5VGSRc
HC8TmCFrlUCQrPZKLgc3YFDXkrBf3JnZLeLET/DsIvJPC1w5tn54vgZhdLLQYeM2LxicnMzHpzpA
wAbbD+KZmtTA30Vazw6kzSBYdXYFLTZTNJBMzkdkzir3fBZf5Dfn54hGNH13hOS5KVMWjrIyzA2P
vtP4Py7u7Jy1wmJ2jvr9+GOC9dmnEmAs98A2ecCBSplMhQucIW0eGE4dfil2ZPzwycX9HwOGmcWV
j3TDjg4azN+S7S9o4KQ6D7a2px+AsTP08Ezw28VwapeSykLAF2cUdGFOlJv2QXPc0VwFmzBq/Cmt
CJaotp3Xw4INFcH7hBFyw6iaiTl6k5GVTJTUjIM9BMRj+JJn5xbgf33REixg4HW4QQeZE/niaKo+
LANfL6Op1azuE5aoXAHElaS3PP9b+R0xsCx/heO6F91eVx8wo6vCuF6RrF1GLPx4HLDhW/kvf2v1
YU6AnK0Heb2iCdjCPt+TempscV9HEB20Z47oOTmzdppq1pbFw40MRnWD/GDs+yDKvXsrjFeJJ1Sc
apvOVPHfdvpK6N2eia7PsJK2byJ/EptIK/H/1ljeYv0xWZa1EDHXded7RoE9q4dFrK/PPSbb6/Yc
0wFcqLMt2t4aM032J4/zNGEAS7nuO5jupuf077h89QLIW+YzSS9jWOw+oVdmdzTFG7Ga8ZRgKMAZ
FL/+Jrktu7QCD9KZPYH9W9kiB/86xawCpd07v1+eXMJjKBV41DeD3SNWBm2rpz/YVrfzGaD+6wk/
VXyoUav08iT7eNb97manyVZZxUZp3Ev9trO2vWmyPOhUoU8qU9ABA7AighPwdQYoUZ8dtHrYIdV8
OHaPnC5lZaH8MmVIG4QDMyqXNHi4tkzj6aFDDT0KarzVaHuCdGsPKymv8FesmskxuayQFoV3qnRk
iMSlAlNL4fZv4uTgEBzWtHv9qEV1QFHeRSh5vcUXHVZZLKyd8QB4RMtSY/P/55HeUpPddtnHGxJu
W+E7xsfk67e2pP4w2PpE0JJaIzI4A4MzSgmEwJNHDKTe3UBSfVFUlwqhRi2eQ9bXeOETcbnl4bjQ
u/pA75uKivXHfPO4AYVhjnbK5Pr+SqMqTj+FE/q5MOOXhNxFcZ+SO6f0oAdPvNgyFKBECC7fpKXX
+7UO9Xgu0MCqFLDGyZI7/QPkke+ykOqoqkTNOrj3u2Usp6DHtYCF7XkSQ/jJL/k/P8eUmmhBFjDg
dH8JJbXR3Lam5wGqQKgLPSu1njU6the1z027bRvYXn9ycwOxfGbMV/7b98OM9tGEDOvxUENOLbsj
YaHv+B3ZSG2ttk2dDXNRuiKACpGZ9uH7KJPjQeCMbRB4SfY++hoUfw5NsB3ksXx4b+QzP4WGTozj
v8Wrb0hjsBpzfHfD5YAQ7KMEh9b8VclUzjGvaPI3FFWkvrnZ4XcWSJ8p91B1WPeOxyY+hTVUiQgh
ivikV+HTXBgf5ISTCmz1W9d9s747qmE0nZJ22fVhZRVjDBTl5JlToANLRwVGiFQiOon6TBTqq+vG
iF1CvtpBWx2X0Vp4WYLfJA7jpeNRMv9a5JlAheoD5MuKYx8Im1ULmeBG8pJGmMFfh57a3zA+i6IW
seoMeRSDbxJdoXVNNxxSh1rlhNduJdfjF/2s4ZUb39craRZuc4Ac+sm4oHngG373XUu+IukL94Bx
HP/uZFAhSkNq1vcBptmrpj9jW0NeE8oGntB370Z/D2BApeCyvvLXmj+Y5P40bpLn68rkEbACLOFX
RBMVjJYPRr51WZOAmmXJKuzTa2cOVl6I9XjwB6X7fv642fQgEKG+wwmg9N7/jhIfi0RFTQts3P2g
YX0bjNxheZ9f8cJX2Wwc1wyzMSFnpuOv0JPz5V2yZtPy7c2CZLFhwez+yOGPn67BhilMRIWFmPT9
Zpy67/JtyhfWYD/h2mCT3O8oGRFstaW7+0kmjsa0S0rsNfHxIIGM4YMeD0WGz2PM4VFy00wpriKt
WeVue/1H7j2u8oGOmMytHGQHBgo2laMwISmaUIQ5s/LTmA1ceWPKjWKbtaCr45u1hpu96iJLLJvn
78aUTvLfvGGB7qEpTtWReGgo0WBANk6NNLhOuDdC+RSgF2ZVYTZTeEA38VnKTxv2DRNLcC//SzP0
cOWQw0GJekL7FdVPSmq0E0rL6fAZivjuf4IrUjUc8CMo+/f2y02rVjkoQDleRo6x/13lesLaRJMj
q5GLY5TT7tZEvz9W//06mScaGmi9ge/esKj9UpoOmLDO4tACHYvElyRpqA0oZv5V0kZmG+85GK4X
sXfY9JpujXFqSgmCWRZ64XWuen9RvEu8vOBeRUngSOpm+vmfrhfdERHpEKqSdJVZRvcsAh064Wk0
+ksdrG4Bit+mUGgBtUfXyRt722cVJhmLNWvydjqrAwn9dQQGoaR7FqBwyfX76aZhuRyygECLoLS7
uls0/ScqHsUbvw9Y2rCk8hDFhC3LSjWboH/QRmT878bPgVKZ8eFtIsu5LPMVmUsvOuC+PMtpeALx
9MF1l+J3bBKGJnGav9dVQcLh+nakr67ZU+qO6MfF2+wP6gtr8CdDldCJJB9va7mlNHiCaRqhxtJf
MiJwSpS5JctGYSMNMdhyZr7RPCVuNOdgMunzTx9YfbJgbjR4TOSMcrHJAb5oRpGMXnR1ua0VhPgf
mdQAxrgEln0q/Vh+b41SVjRMgOCxdj0gzW6EY0GQbPpVpiwzuC9D6PgVHmMlq1dIt/3yBiZb3mlk
GiU6vUTR85Ientpm8qkfZ2er3siw5htsM95Jx+Gxyq7Eco880BsZR0Ivq+v9AjHvwBzjFW3I1O4x
9Fq9OTPmfpOzSL0jTsn0ZnwUnj4taMrdIy+79H3wnbcBl4LTRMDN++XqHT5n+0752LHrszUrQIht
jjNArW+BbqjNDaKxacAwPVJkJIb+UdIugGyQiZG5Rtt4F3PlVHWcG76h117ycQZTLyxYnPK9pK39
N4SNFmdkqZkv01XEDNR0cbb0Z8iwgQ5wxINN4welWG5gIgxcPmOqFJmUNbASfb/PZXSmcBzyomAM
Oco38sBrtKc0Ne1n4cjsG3XdYBSaiV18LOU2g6frZDBTao6H5UfVCOLzrJXJafDN7jpvqDgKWGI5
S/XZ/FogFI1gvdUX8ez6y9wOvgNtbZ2Lu8van1T8Pd1cQ3od6XzT3ndWqSMFDPogbVF0wKfqPgKe
+mQZvR0q0Bd90LT74zg7DoOd5fJAU9Wr0ghbABi9oQkMFOeWamB16XvR558zaI2bbWMB56e1WhXG
4he256DkD7PrykgWuvdySD8AKKBehLoM5SgMlDOM5+3TbS1DFchqCGS3nucCruO99X+I57bO+X2E
41fN0C7hAYfaYkBmK7JzO10p65WBbTS1T8ihkhp63ucG7NzFhwq5fEI4hX+PfZnImFaWMVE+dZew
3X13OXEe0bBd0N3MZs83hEOtVt4T/9yPBkDlnDH0yhHsv6bNWrW/DdLD2oM7FEaiHD8E7RTYzc2J
KgKQGWLPRQ8jfjlRHn+Sm3c19dsR8FtxEuYBZCcppdXJ/6sZiSUQkf35ZmCzInoTblBwAtZscY+n
J5543IdTSX/tq/fIZoUZiBU+9B92kRecfjxUyS7O4jZRroxA2sc3pVDDU5QkOnAgATpVg4r7Vczp
xpRXU17svjneA0N2IURtyzhh6VKRgoex/6mCfF76ax1JD6XEGl4kqkNASGDkcg6D85FhoHyKuf4/
wcrO8LFm22NfLR2K/1hdtM1XbM2ZpecKDDOtg7eppG5GmNhVEW7MO6miCkQBe6P/pdBSNJuzrUvN
RIboKw8CAggsENefx6R0dIdigzWoMg/SKAAy7NLQM/oq7vYxFgzg3zDOaZ4mzXRMca/2W+/VU80t
dwwAQoDtROOEGX+MDeOa6f+PJV/oNGU5e1sEmoyf5morAHO0RvlC+aqDA5pa+yEEumIPJgT8YYjg
EqNxh3Elxpo5asaU069MpuLcXsCFHa9+JPASkpJTfkZpHOzt9Cb2dkapY8RTXYd65uRggO7eqcrw
9hdlUQBVFiRYOIqXgqd5ta/WNqo+fSvmtZKWqnof7nCrOahRlrdoVyywbmcSmMJ6PKiIcxe8hw2B
+D7mPCHh0JH0vbeAbNQww8D/S5PoH98t+0zUuD6z11KEqOxdev8YP5p01NHd60hqjns+kH8SsTMa
bqZYFu4YmWkhvi3G+RG4I3TFwheVOVj3CQkJ8MDqXqxEN4PYLUeqTgiGmDk24NZAu0Jnbi+KdP+l
f7etMRVnukA0OcG5qxPcoHFcwEm3lj7PDrdXzH8UioT+KOgCXbjgSRevydH4SEfpIusSW3cPzTyc
EjaIlIZNdnUGIfjC836hMTOWVdiaRDtFdCPUAjUoH690otiItduJgtMe9MoLNyIo5BfTMBGCYzWw
1Tydyho2ecvrhOgws+OmDN/kXeOelIMHeSGN90w5wkHzKuX1brhuqpSdZluQUK6A3jESW+c5Jm56
SnvrVoMSORsNW9rqs+u+JSzkgUtow9dx4G13mQZoFCJmqj00P+26f4l7/tHsG5U085h19RR4ZS2f
WGaScaYucGKyMd/PwCnBp6DjBzLYt0llEuRCNJQWy/vMBaezm49REOT508FL0zhPKD5Lp02hu0h3
wauUsct+d0F5n83JFyQry46i/APQ5uEXNNXkdrt5j8lA9whh+G8Xa9o1sWRwtEsJtFTJCpGq5AOn
h/F7EL08IFe5zws6LPWwJm/F1LmMLC6dNByv0kqxYLmLLpW+R6t8uYDQ4MgWRtek04sISUtOSL2w
3TICHPhzI3Qx+YJpJasi2ifFqxExIJcw5/6DGex7nUclAARWOchG4qj4Fj5qQ1cskoWu4EiTy1a7
6zG3v19QU6yIgCst2U4BfuECk6prWAzeEa/c9FqXV/i8zfKUbCa0ELWYfjkjNP4Fwuz6HBGtgC1B
CYLzm7I56lrYfCUZjgI3gzdj/EKr0ggGsZ8xr4edhkquvn9hoXuqyJzjXd0WlpEwfCKavXPI7fpQ
AR9Ui4ESbBxvX9yh9gZ4rmw78GgHJIE1a9WLiTrowOj/Oav096NkKHKJVyrQ3i60dXFkhyzz0J4J
L63x3UMgCAb8WnXB3rb8nNKpHH/W5+ZznYrXi4X53uYmt5gAf85N6segL3vvaZC8pO1XIX/WRrq/
m7NQLR4fcaCxcRGsGnBa1+KChsdl1hUXqZz50jRXkml7EUFkwCmzd5WdlKfRxXPaL5VS+aBl1wB9
8KXq0nTZoVh3HNvoU31llrvUyON2Ae4gecz7ldCdXdfdV9wMMZp8j9o9tNxN5QOcKk/ukROAliXw
zQO2/W8GbB/gS3NRVqxvBqN2AKGHG+pv3Me/w4ZZF2C2NgUQZPoEnDaysHXbYOKhqF65nkb1o2mI
QwXY4OA5hxRzSj04zCASHV7Os7YW/pLnVqVHA6L/WZGbw9x6ATaYsBux2G+XQ+5zqdeV/N6/fxSa
O8j7E8bSqbnGhszEUU2gNcI4kzlzN1hIhKWSwnv5B7VrMj6jsmJYr3v1ksIXYzsR6OSNOhX4YzgD
c7Qs5babg/BUvdSXfbU+IVzuDuxP/dnJWPLFKoLS9EdcHucLr0ZWqGoPP5wU2+vQh0Ydxws33NjW
73yywWTxfTDftxaNhePNc7Cr56wdVKM/oLVjzVuZ1P4zHvh3a30iMGteTM9IwN1xoZE8TCQDzJwt
S8d7af0cMmIM+2OPwDdBWbTIfH3Tv58673HJ6WVUVsur3HqnbXzTyPErK+mDMkYd8GysZBiE/Hn+
qsS9cb0WjLIljACNzUPlJVw143R82CEEJGLQwgim19lwoUumWT7L2OJCksmXHiAonOH8SbvIv6Ou
fao6meE4SO49XVRGbwCUKI9+kitzUHI6i0qcyBjtB2kB/Fx8CZsnAdhb/zjae1KMbdtHnr1C2SW0
lVRlyfAW0qXb2ctsMiVDmGF9CWtXTRKb3sneNy9oOpQIle7SoLAfiHmTn+XiPjbDgED/aujy/GQu
Q/4Ctib4cqvcsubclV2GIGg03L65blFERiyrKL+JEzkIe36DQPh8DQP2w9BK2/z/QqRLKgQqIkFk
QIIIajCFDnISpFYogfKdHhSYmYLSWffupG4xxWP8etLRreRLQB76dbW9AheVvOebxh6WQzqqiKyY
eViHT9SqhaxsDCPuNiS+gwDa7lN3eP0cIg8/LYaRGkoFDPEqhHq5N6+pCw7MGTi7DbEQMzYvZw/s
Zfzk/pAGG5mcROcFY2Vnu9CtO51IEbjQf28mOYk5QJAZKwbvJkhREzjumYXP00iYgicjlxJWMD9h
jcebWMX+/zB24B40KeFFfn8SjdAySkUyWGklHPevXYsG8y82ha1vhPojRsEbOAJOrQB6pH0ofIE2
0SIqpT+KW28zyQyYV2XO1OVvJwUF2j5h0TFagBXwk3MZZ3NWvvvJRYd8IDorCnYdjgN2Nc/RlCyv
nCzPWYTKhVOeu0iVg7T64eSbIoZJbZgvSJA2Z6MRVWis0HfwTNpwgpthQ4pk5xEX4YxiYyi1f60J
slhmXdoZgN4bZhcdJaJh5t4nLWaeteLRQY1r4sTQ8oEDbkc2j6IpAPr9ftw9ow0hFTwCVggmYYIT
Uq0wnhdtzWE4549cnQPTA+vYJSD+Dhp60fxETLdjCo+d52siFFacagKbguhw/bKa0DpyLpE3krj6
7MaNVEnkKEWIo4TNAQWXpdhU4acmjTHy+tE8q6XX7P8pZ3Uh5Zjt3/I8NuAkCIDNapFy4bRzaOoN
pFJY1+FyDfPaSPj6vTfrFovNhIO0ciJaSqhlQLOzSgjP8Eqf7ScfXFxprOyBNmyZceH3OiSIGx4V
hk2qHbpEYi08IPC6lOtmUOZHfGS/zPhqenKtyIWInprx2eFKyxuh8J5wOwkff4dOTAXx6H/GZig+
FU6tabjBxOQUoy4rb0bf1sqAn+mySKE1i6VaONP9oMApZKKJHg2kr/zfiUgb/vsCDj4Q5C9AQ8DX
OXEDJGyrHKzxsigA6HxAIrvq5QuzSIQ74UAkIbZZL7wQmLsG+EbCZ4+lysp/EJLMuYq07RaJTRzE
ZhoyeUMlKjucoMFNZKlWF8rTp2/8S4pT62YGb3tKDcQAbvrnIwIYcgG9efmBgr10y9JV/F/q8gD4
ClOblwv00fuWElF7N2sF2ou3fTWOl/2Y+PkRt6nuD/a7M84stQFcy9/V6luNHIzBNu0EccmT0tbP
GNygj/O/Pau0ciG9redchM0i8S+juIYs8KbT1KC35xoaJ3cHmMZQi4fCIrBaQUlJAR4wlv6K5dKj
MOZ+v24J7NT6hOfQIFpRlWh8m+1vlaTzh6woANBchZIheMzG9++Kz4Yn1V6LXSKnPGee0zG/1H5E
AtLjWlXh1x+9KubfiEaoT0JEwy/STQc9qpEccdJ+N5ixmGJpnVv/cfl8aDh7s97shPqPBRehbCdj
GC2Gtw832AkfSApGLDaWYGc8+RZkBfaYLslA3gETiNdZi0h0OTexmwr/nqi9VRKyXT0MigPpdBu8
dW5u7DqB+6fXTl7VyhR0sr19CiqOLbbeQTkl0tM3lDX6Jo3KBA0WEK/AAhSTNI7DGnmEAyoHShq0
1+EWGJfAfBbs7/Nv6z/wfawnWcacX6fqZ5orbOz9sZ/DLvUrCulxmkyfOYMdywZVlDdAQX3dliOH
aZixaEHidWKOmbqCrl461UILl1WUKDzNT0wvAEEziFKbKNiTWJ2rXuCVPU0t+XDja/hOI7s50d4V
0L9dgF3FHFdCkqPKjAcjasLr7UmryGxdSYiti3/n2n1jXD5RXPUm7jNFkHmKEuoDWFses67T2yJZ
vtK6k9Q11sKZ5LedbGzz5SEizq7urmaUoPp1NL6vIDgMHedt/6Z2ZjFvpoeyxl+7VL1Fj5qgwMYl
wPgyP0vwFlQIjVQQ3vTN/Rb6y3sOw0Wg/i9BK+RFamkHVfnNqdGrQzRg3PQdpxYwxiiH02myYc1A
pzlF5reUerKYQtcMfqlLixFHJelPg3qeDNgwkucdsesEMEq0Ye43KVBsG1fZvRAG50NVrT9Awljl
j/Svl5N2whqR0YZPItfiuky0NVsuSy6dOelxtDdhbKUZdCuAh33R4hDxleeiVUTgt7PSay/mvGxn
vqTRounTlUY7o1z6byjki1G+/GwJOm9o6j0bMUzCLkU/zJEAZDUBGhzPSwzdnbPDcly/uRDbSmNK
1llTeuzQP/8WBo8bK/kYhy4BdOUPucoo0c7csv0k+7wPQ1pUO1l75jHl9wUOLXMKhodvO3OHWL3p
3HjdgjuPnT6bIpDX1CB4Uc+gG1JXiV7QEvTZS7ogX0so0+yZKSzaWcFCFu4nNRPFtUrJnNV8f8Vm
3pC4r3Wz/IKl6gY3ZajE1U/2cke/v2+AEBpHyTfyKu2lzF+7De3Wp9Y7qw/7sZVAkfN9kH0CK8UL
OSAh/b6XWpF1d16Zu6vxyvlb3yoU+ZnDKGVfPctDTb+BVoMCPEicAgFlP4JzqxaKiP6H3zsKMOU/
jvBMCGvZ9DELnwgODEZ0nJwFzCNR2LlZyzRi75w36nxfukPOER/SYvMblvon6/dqDCWEa1k7g27l
eTvne4g6RfIgXfYrhQdMgLMfMNZ0crWuDXQwkF8xMgFOBLxo0xXXoY7u8pNyAyPqjHSYOJWuTc6b
JgAMxTkqUlHT44o02ubwrAOVvgg0hSO9VZvlmYzbGv/3LH8kSJvxM264pX+ncGjjPosF9dsdonRr
usA6h3h971snfBf9+Zk+usYYozUN75F5HlleVxW+cUdaH0gByZz+IB5VSi/4lXQOPp/oGy4GMHX9
3hZ9Q1Xu/qPWyxbqofCtvFihQ0/2WwFDNajNNtaNrSyEXrwgPgLnmEr9v6vusBAUQMXfqAwnKxqW
vU5l6XQRms/kWBNDOMcEcaVy8cvda7Tirj9QFcGebnlzWfiSkWDYFBdey681sdmeZ7mQIJbrSY7D
gRYFOVATk0+QBC3W2LdEavWluiAJDO5lVRiJ6q3swHJUAoPlzxVT3I9n19tlwBF/PyZnPob6SibG
juws5UPBd8lkZ6VYywtXiTPSHmSGIr+KKnDniZYgl4Nzlo189FhhfS0qD0BHGmfCu2WEFMMDerpu
Dqp+RU2ZKKt/WgppQspURN7eAhQk5vaZRoBcAtroIUozFAe0DM64YvCTw1665tRSnpdOGziE8H+N
wUXpkVYNJ9UmsBThDAjCIIhtmzrK8L68NqFo17H2ChicUVe5y8XzCyvGsYhzcBX2VTjJzyw2Y/GS
al8m2McI79rsp/Dr04JbdACaTP8xq6C6MqbBNYG3TZVsvrHUsROnj/TUGcmZUcm+q8BsXRkyscno
X4HBYmi55rhn7nwCnqOWRj1TMwrPm3l1BVYD0MeMX4e+YLuphSPsn5yiMywNPybMJTPtcfHV1+5D
dTTAuRDnPiaSriC9k9L63Ao8hoaB5EUGSzW8BmKtgPd3bEOr5d5zt3ZjFmSG9I7WpBpiOpV4HvIh
kLJqWVgzGi2LVdTkRvw1gCKo77Cqtd5hm+nWiJjBGoQlYxUeZAQDRKZBfWSD2rEONWxAYX0MupD0
llhvNPgogIUOaJqCNBlSP28q9b/WEASFf6b7Vw6XU6teUkiIIWZM8UIeYqNXQOI+ZMxiwcTVhHof
onGYvTXoogy4JsbJwyB7G8KqecqVFNJ/oAxz1Jvk6jPKbwJp+Tv+UULp3X0i0QNNCqXF4GKRWMsT
tmAWhfv9ZeRL3SjRNmMcDJ7DjETiL/XL9pGT2W08DEpibBtv6fIHlQrrqI+LU/PAAtR9EW8OotYK
3tT2pXjxWCZQpFYpe1pWMqQ6EendSPpeK4QRc5XslEKTKOHB+M76CxJkiKmPidln/aJuIvlEHlgh
ZFt/WETheqyi634gh/HoIlDT+MRMxv+OmNwWOWIOVY5bI1leaVysXTZ/lFvZj3pZgmTvXhwkSJ5Z
Oiz5V7B5UcXbx/o6P/gNnm4snF3SAU3ZMc6pbNofXNUwnP/va+5rqU+N4LUxz6NEJrTQJkeQ6Wsd
toXE5YhGnvoT1J60rxEjCDrDRu2uz0IyZgZqCMEDZNlznl5wsXAbDQIb2262qdI3YB+eIwmAsHyP
ywh0k2spu0075DCq7UA+EsR7TXosfGWrYmGTGN0WzdTIJjvhL1D8ru4zv575HVtn0zE3+AokVTwB
j3AoCqB3z8Voql6x5BzTACByMpL2jMN1j3PLp+uMVoY3uBVIG9/AtPOnNOp3au4EaiUSk+DPV4Iq
gMRnEkZy+bOj8HRSVREtESX3i9h8wV3TrNTbhm/cIHJJkFu3ZUPclFYSuM4Ki5dOFpwF3zWDVJep
h3sly71rHbFOyFP0bAmFKXKywJU58misflYRO6JiLxUf8ZXg2OVcQPSYnnau3gx3omyWxz0ZGoHS
ahs8CrnSodY/cs1JXnDMe8T9yGKOMvlaILHLwcr8j4Eb+pfnYz3+Sa94yIP+hUnzGdK8/kikKlQf
4ehgGvDJgWxhdf0S0Sjcd3p6SdpKj7bvdOPBMdCB7S+idsydlI6qxWEJpRvq2Aepz167Ry2mVce1
06Eh3pUJoCtCIjAOgus/aj8IkOjWqQ+oG8B29U3tr/qPJiJ3pdrz1KiamRGxzrJ16zbY4DzOIeAb
Qg3qz8lcFRa1GQkVDLBNuM0SmL/mMyomLyRUzvIHziXt1UKbiMTkyOlLwG/gdw5p+SzcLfGoF+TQ
d6aaxTfGEB53QhgStYbPm2fJzGGJVxNVguojCOTcF5HXUF/lA1BQG3W5YwLTp/tdItpSJ5UYRKEH
gxRLAD0ax/lbeca1dkbYE1VLeWZ0s/tqygdPRSdOE9vDf4Sc75woErTuk1B3/zkt/3ypSLa4Faoh
kkCa1c0GOcSFdIp6HJx74kHYw6DHamrymM9h4WCVf5eUU3j3MeZgL5+acqr9oatLCaoURBHPqe+J
+LNAqk5kTxxYKJEedmu3r70r9dqPDpb3dnTs6EZTTytOLXICCmJO81fZcFW9ohABjaG/ZzYq+vUP
+xXHztxbRVVmFbm4Dw2LIe3NJ97gdVhTRVA7QWDzIe68QYwsa0zv/2HBEf4+b9tHZy8cigXXVuev
rORjrDuZ5++HaFPVwip6fT+lLiCuKX4HMwYFNtW7cxpKBLNWwmtPw8EMq50qWR837A4RiPZnT7an
dCwNxW81KE5FOP7C13kbbLof4vSfoGI7qHguCpK9YvatLTeH6Lmq7YmAV3Nxwlraooqg1CjfXvdl
QSwVk++cip5G8sp+VEJRtxGtYXI3jVdh9SWFY6uc4+4/CMbieMzDTffa8qJl/21eHo5TSKHXZku2
49dycC/DdKG7Xj6nR/Fw8++Rj3iAV6DTY+W4HT5DeLPILVEqmpt6il31sdbAfvUqSaf7GwoZOH/Z
St2gDvtP4dPkfsQsZxlAHpYQ3/65xLbJN7HS8VGVebIHE6kdgiKp8EgTnvSwypGaYie5PQzGPThy
pneJyaiiHlsBOzu7hy0SmJuzAk32V/xNJ2/s5pmu3xwzzQFPM2VBDYV7FOUQLojEsaPzZWQv0rty
T+HG1/710pa6MjGO/nhJKMpAjTTx+mlvbHGc5bXi+tktXGeF13z1cT/mEAWRaLlsItJ8s5nDDISA
z9bHpcDHsPydISyZsRitMhxWd/Fzri7on6Ipp4Phn+Kdu/ncV7IdBrJxk4pkr6nGv1xJLGHZfq3G
kCTw3j2ogEfpetcH6ggSqwGwGi3hiNQca5f0ALWchqQalp/uEC0+3GWiYzRR8kxodtH+sW1whfJ8
eNXst7y8PbAGzznksRBCMQl2cr2M8V+YAKHqNsiYTs51Yu0N15kThMXKVOqG7v+I9e/k+cQwvh9g
XRZyrURJWOElmvxbQ939NEdW2tQiRuetLVGuVe18JXdQnFAv4uTP8NN0Zr8NiOJYWqYlo0TEYUFB
oZ1zGyxFva6wzqsdtcQy9u0Nft90SR8wmDelA2fTNkvJFsUz2AztNjnWd2CM9/T3qoe9dP5mgUji
fv7UXqcwySkBVKinq7Be2FHi8wmUjOkAuc5OULxsd8wg4s7SFtd/K9Cs3YGxnbCDG/SVntcJcgVA
geZbSGsjFiynuiLuNxNQITZjVMFbcIGh3WcAy3KtPvELtT+qj1NwEzFdWNJYIsd+OIG9ncBojvYG
y5xnlmhagEd6hpQV2fjy6AqFnJ7Mo0CZkdiFzllfFMObRaG8m/t54Pfc78Mwg8peiqERlWl8S9T9
QM81EXT/URUD5XkTy/iQoM4Lyotz1j6rkYVZW3GcFO+dbeCWcAdZNWe5lHKOaxFw/7AoOpVRqqdU
NCbv+3TVQw4D4QDt6ZiBZpFVEwNT6NkyKrP9O+An8duNamRYXbE/Oibde3GxUNppF/ktAU+l7y47
ttp9BusFf85o5zzzG1FjzmBKtgtc/7gOc4FD9iqBuhRfQs/V5XiXVsAqlSJKOWcg8HCL0jEx7dak
zpEjk4O29xRnYja0DuL/QvIqJMz/5/sj0zCkPmLE9JAcKFz/5T5ejbEbWQvMDZK67mAZnHv02zrB
7zjX56uad6ny0cHj1/i+aLYlzqFbkOGRC01jGlwevDeaptMgnk8qLZhZ9Enrjx7xBL+zmFary+0y
9cg7PzTgA8er58Iyna6HIOcrKBqN+bSXlJZgGccYilAw6hgSkDY4s0LstC+RopJ/c+U2Mu6Lt3FT
wF7cu/lqDlDqYfGF40g2+F5/odKsG6la2c1GKZvybkRH7G+HhxRdKmi2eAU3+X6+vESLPrnfeZod
1rhBIg6kP8MnQIZTPOB4jJG9rdFrqx2dgfG8aokgpXPc9mLl22KwvcH5A7oIZ4pNuLOzlEyO800S
qL6ctnZEX5vc5k7J6msElz0v7S6ZKAKPESIPPNt+W9vtmcIASTpdZJo4uWgdG7C22KHAHSHz9l5j
MvUr1fQgGMVMfyVWe/p29bI0pb+Bn1fugTwSxqwkSVVauWawkGbaE6fdbcf8l2GytULNX+4Boq5P
DiO8M5QhsYMa81bsN9LyC1AAt7XxRKFUMwEafezDtslfqfX7wba9y3tb1rGPS3P2NcWom9Lr+ytD
QepBdri7KfCBLBZAgFn/3NlfBIKZcdQChd4GX4cvAK0kDgN70G5MfF0ttIQoBJ9ABGP+jPuCHOBJ
tr7qmwvMbVf95AE55UPAKtV+0hesB5FhW82hmU8r5oOO/3D+Y+tpzi7asCFpuBEETWNN3vzpQcY/
5+OHNOyZnIG4NrZlT/gLVN9ZOKHb5/0dZLIodWDiGA62WKJVW12OhGCQGtj02MmoetqjHg6c15er
5wls3CJUDPEP7qOjQN6A8mr+qgiWjfrQaK7xt/S7EKmh6fPsnOQfUuazG7RbCcDJiIrd1cj0v9uV
X0dQ/luJKI+7lqzId/TbwxeXcZVNGu8kYZ6K3mahKnumtuR54YNAerC2fu+oPucVbStjQZ8xKzxY
7rgdxodaNBoIdPTVr2fCNDdm/83qNXNXIUint0UVUy4KGM6Cxh4n/eyssVGJCVmw3Lyutqyt5A1i
Kcvb3df+rWQdE08qRHfr4BCBKPMj7TK96wf+fNdoordept3j0SRocAXmglqxM2GCD/08TIvUiqZ6
1lipag6uecr0+DJLOEYIGeA9bwA3FmeKNDXzhjxK5YUCxch3lnioyhVXLZMWInzt8pQ1QapJm+cw
DWdSYhnud8GqwlEVd2r8SefYE225JzNuQCxU7vMidsIXDfnME7LyjWarw2X1gW1knlc3GpzqBNVG
6N9Z79qW+0pUPTpDTLN33C4uFXeddJL2N/aHXq5RgZ47wgSOYypubKuIP+/PAVvJRF9/pHAdOYw8
wyFZwDOtT6aX+Y8PzkZVfoS9Vg9wRyB7YHS3i4j5j8hJ9ydzHuxJI95fgWyTjhYtHsQSAEkuCfU9
Ug/FVZ8Sh7T8Ili9KILE7lIMHldm9pu7Pomthp2C2QzodhOpuNDfx9/wBFFOv4MGAJ9yiHQhZW+f
2hu/COIIEskKM4xZXyvK3+peNEJfLLsWDwv2Epb/kZEZB8/aRB48IDzA1R1AFFgOR0Pv+NdkBJXn
CVcZAUgDpX1AdjNO20uSvVZj3W774pPysY4XVpbFOmH6MSRmM3Kc0oGCgY3x9db9lsDvfe3hlu87
fPR+JaSIuJBv6IXgXTUPoGGVViX+iNt9Hl72a/wk1YrC4YAOLMmWhJwOunyvKq6oaqrjdDV661Pq
AQSwI84S3HoZ6e3BtDe7FZjb/M2zf7iikRWZJriXQFxVnbOiT2g9AMsGo2L7/wbjmi+qdDktsBJT
Gz2Jlrsc41b/HaAtJgh2B4Dsd00zv4sYP5XXGFOB1tfXRxPn4g8oHeJy2suKFZNM8Or26IxD3Bs+
j/CWQB2JnGHjkIWVW5skGBnBSEHCCX/J/0FK1rLpq3c4roQeSZAidxpZjRbDxwJ7Zr/S4TbAo7qu
4GKaC2GmyejWtUCXdvr1GdFMu81crbHbpvnBaI9gyQr/f3rY6wZHnCgrDqsFDhYtKjEep6XECeoL
begoGJ6NlNJ/G6atDiBLkEDO4WMVOqIqnSOHic94SiFA56iAEdlvjO5WwVbPk/N0/Z7GITk7iPD0
yNH0ik3D/cCkvsMaxdfVmUtQonAPcC4RZwT/4icBDdjDFFKwsByBDynfTI9Nyom2Yo0YJ7cqPtaN
UO+uo7SQS383VxQeU/cvITdvmvFI4Jt0H5g1mDLWxg98o9qOGUZ47Y5HDYqsyik+mplKp+ycXrqH
uS62/gKHHar1KnfNfyOETmga107W9p9kYo5eROTCDcRP7NMcmSO+AJSzkO/jYb/aZUyuM3855IOi
wiN5g1u6Vxs9ascE38rfiCt5m+FU7bHRnBKh/lxMHnft4XI43G1tqGgKKH+4BElALCCRNmFlv2Po
UbbTUPcBjpQ4hAjBzSiWRy23/im/w0dcO/4n3nnrNYiiUZBNh1goqfJHSgQ24l3uYOvwkmwTF9n8
Zr4vhAxsx3SMePHx1wxYjA8NFPop6Ji6wkmRAoichle2saN2E5PuPwLdYWHXc4LGUlN7rBhN1hv2
FHAg9jJnG5/5JvJjL2FTxU7o3xpxgBB04n4c3Zfeuyo0i5KrunfM1aa6Lc1C92fB+NtxEIEDY8Ih
g7Z5X3eOKv9IL8V535lJ5B7xMXkxaup2bQoSu5T1cJdj/uuiRUNBy/FBKLFndCiWe/zKZ9C0Ud2z
YZxgOQDdfQjJTou0Lqui69g1n3VdlkJZlcF+kArv/m32klTqAqCEbsUyqauYeBWhBUDteraLHus1
w8iU5hx4aITcGS8W5efdMTlLl39FJOxEcALZC+kXhK/Sn0yHia8rhAEt3NOCHwx4QSA175GvrXAN
UFT1ptaAOb/EGwi7FL30bY6hfgN/2k4BzwfO1mADaEqFZNJl0WBKABqmrJfGRCoZeG4I15wEnvGg
0yJ5Z/CCWVG5xmgDT2v4TDv2+PmRFGos0NLc2QY09hI5eXeW6f3nJSRajKgT44RSMXiusa+HikLS
77VckvUx0x3IX+QHtudS0wn+krN8V/PkBpOSF/Zl3CfJZAJqrBnM83FLMWY3ONZeFBMl113rd6r2
DIU/xkfpLg3zK2gA26q+2ZQ2KMst83ySt/ZbLls4CcfCnSVu4BIJ8LxyO+v5HumgQ25pkJ92i6IU
SWT/ndQ9vw7kojcHgZvFrmX+g1rOdLA7Ld0fWDJBdhoCbth2/Ugv9uqHZokuhiLAYdip9w5A7GAl
jQEbiEkKxk6Co9NiSbS0Egbr1pjI9ABqvcbLZlArL035ec0Pbgsn13hY/oBJXTttgRdjXDF8ZqzO
RgRPm9e7+I050pbe8ZJQOBJ3KkyPkpkx27ckXqY7GwssYP0qwFFalzWhRSGe8qz4SRO+tcNgm7NO
EOIanemF2ZZEHzn4pbvZ7LioyHn+0LmLZQcbeeTxqa3ygc2+IzJRockaR4VL7za1ilwv0RPJxLQ9
ua6QHhQCF49r7iHRo0Y5OvhTIHZnWHjv3jkFl2woKKASXnnAeaBS10nfVDUWK13zL7J9y783zRSt
1Eh7tcheG3OmbLo2oe3C34GAQOrgZPzu4A2zdwaNOZaRZklNYt47cTytcJrQzRMQTHKnPQy/V1Ah
fA7BeWuYvdnSNgRVkfKR5qBtIPoalOoTptgL2tWdNouO+1YyZa/UFfcQu4IiAEMvTRSKVJoCOACh
S7RztyHhpbZJFngDwwNvhDQF4gp6ClYHmAyiMlABOMz6jJW0hKOvFUtUgFHw8V692J2VUrn6o0aE
f1dkm6aSfGHETlRysEOMV2P3Bjs8GseMIHsuufZiCXKexqsnQgSbRjyKpnQMJFPQfbalSe34Yjw2
ktDCoElAdMUIIxWZmc0gHoQ5PqbvfwJ9Z+b99BgpLvOkxsq0IFtOJnPTjfc89TClgRE11AWaAivl
1REFiv6YIYdnGEFOh0He0qja3EhnW+QdcRSVpipSdpK/srzeyhXqcuXBse8ibw3SHk5MA1wnL7zf
JuF76264QDMqMj7EF2/ne3QZOg96nY/IdSNg1tD6zzJcgfcYwTB3MXf0t/o927vNLfzmd0CI0rZF
SYLGzyoiTK1exstyLqNBud+ozMjqzbQKBQ/VHSvwpIwgZR+sXkdVX2GaksiXCyL/zHmFZ/YA9ZYn
p2yoGleX3v+ieOngUFax7Er7qbgBZ5rP/rU076yE0mzeCZokZ4JlSy1+soiyRvDZamufCn8untm3
8SNzrZQjXXhL5ZJ7bvShLgOD49S4hgXFJNxtjGQ7JeMOoPT40m54tKyHnxG5yscgcQXZG9hsAJi0
bRJsrJng7etbiSpFjknsmSzEuhL2RyTDLQX01oY580EkQa1jfRU8lXevj8wg+VZ+H/bXwFw275y5
vJVuDtE/ZS0CgeQEdkvm99UkCYsbqHZ1FccrWQ2irmTt2krI5kAnjomb9gl1ei4h2GLyBZRaTVW7
G6mL7yMYyhgILko3aSXlE6OZjwBQI+iLCfHzzb+WidwlokVmkmvLsn4+9m8OseRCiP3/wuhtQ8aF
jt+hlnhnaMAVjWexBIiU7uDNEEleJYjJLTA0T75SHFneBQ+czMJwMiu6kUut1ZK7Dt7LDEf/Z2J/
gjHLGbxJneuZJOXsR6yjfqAS3jVIm5K34szDQCYLN7dDKkYZN8vgh0UIoWgG53FUD4Va7W+T36hD
NmnQ4ozHRx9T8br8Un+W8nnHbar8Q2/Uc2NtQm7ua+TlsGC7Z4bZau7PMH5CpPApC+UqF9f3MlTu
pPizKdvM8Ee4J5Ewh72tFh+ciD9zGwF9cooy/cxPFOCe0DlLa6SM361I38zpK6kua6v4GaLLKOoO
hxvBfmEneXpzZghS04y31cNA7xiC3SjL7tjw5y1u1RBZzqPTVXSOOcjWCcsYIOy58H2JSWl7mB8e
mg5gXO6RmG4V9k4FxLTm+XhqtYGLcGPuHeypcp0224yrRcSkYTQXEHdTrO7qkb9vXRjE0o0yuN7L
yo4EmdCCHBue37Xc5xOA5Axb4oU2x4/Cbd9VSzgc4jjCy3KhHoWFAZHeQ12wx3UEYxOosaHlWanK
mPevTP2wjji7bknNKBT5LZ4f56DIaSuVxwQJWBM8QdPutz+G4WfTU4B365ziNRX86vFihPKjdviA
/JHhQjp/GaGr6bfT4IMX5HxTTNYqaoZxRec3uUu4tmKK1PLgmT2wHDjXU70awnUvKoo2/buGtOsX
lZeB5UzHlJTl+jdtxza8Wf9Fb1kbGUYc/uLmyp5354QLONmx/DLBela0nuc2eP/KZHWLDlP2zc1E
qbt7dnfm5OpZPhmyhFgN0f5KESC1Tiwocd80ydMFUvW3NV/SpUGzwkf2j3qnHkBE9wDo/B9AD0Sd
6W0q9IB+DNh9IqNd4kwRbFfEJABerPseLSs/dax2pD56CTeerjnAO5JuKPSzfofZj6Boo3xcTzLF
ZCbadpmmA+so/l2Ai8fv34n17W03w4MWAdbtJgEarYYHB4P1fPQNGOE/wfIZkU7gdhClFnII6oBR
26Lx7y+fqdsUxgF3llExXO7cF60Z75IBFvO3okPIug4lWaK3kHY4w3fypwvu3Fa242Em6KXKolUK
luOhxtNhwYQ3NwEK5mAwnMAomU0hPY1nR0UIiDiwu9mjEpxlI7Gt+wFoI+oc5MTSOsOWRcRGy4s3
EqF2tq+GX8M55gwSWFtID1d9MC6gLg8fBDRs/v8zlIzFrAqwA2VEE055RW4atzSbJrUVpKNkfRzT
9ju02XMUgTxzp49ECmcGoHUSuSnhePewcOIRit9sOLG3Qs5v1W/mgAmFzniBQ9A4+ZLhq5AdMj+D
wrfSOM4hM6nhNL8VDrWRFseBVSI03O4iJ0KNRmpt2XQXk45FSlwR+mLqLQXYJN40MbwLMWiXdw/2
PO/jDtQZfbCr75+fbvTNn5hr9ThOaEC8oMJVXtD3rENW3p2mRAy8yiZO1Ky3kE5LrMCU7e4OJrI2
CeCxBEaR9XU3gCVxSEHxxCmikbHIKHh7zFR+XcADztvmKY04ztVm4waoVUvNI5aIXE1Kl0H+5nO6
1ydSCSxfd0zEsbB8+9bkRHTqRAYEEaWafHkOSqtXNG4JjR0vMv+7CXcw7Lft+u/f9HhWuo4Qz22m
7+nUofgYsahiNBKcNmXwkGzz3VfHfZldIsjTQrkbknzC7xGOYLCWohufH4nrU3Idn80+qAgkaVIL
et/GIeqX0K1Pzmf+s30ns+8CwSd8+WdCKn2/4EDexMRuZmrAJ2DU4a1MEbmXp6gg6MenNZFG7LDN
PzaZ4RkoU6TDn17Ex9J5z+HCfrOs9fVa9CE1sjo+yj5kxStnTNpSHUKf5I6vq+6/bRRrwPaBwoJU
/7kpj4N94Kec3vUiT6TURLZab3v0g54uRf2AipjxHNJU2Zanp0eqKvs+hvc7Jf6hgrisTz6MW4x6
+WNrYyDbvk9oJOI5LjTws3OHOHI8Fi08xxj4KZEjXU3bHN7Smy5NUqoZadpq/M3H4UCMKZZ4y9oY
sTNHrkvvjuSnwWqPEyrD6hQXNz9nvHbv9wF79Pj4e8oiHqIpWC6QN/SdgJ0fhsz83LYlXhG/Hdnc
pj7oH09UjLaZgM5PbumjL226oOpeuDS6uqxDVhthZUcKxBnZqSw2PqK5gijH2pLrX7IvQE/0Yk42
5v+lWS2Xv8IrVetAXftGyVhapSGNEiMDKOpEEV7WttdSysXIGJhmCDYp3JmpN9YMsWnbKoy4GEHP
n3G+WoDW+KwwFaxcZO9uONSV4Ai3WrtXosZXH0W9Ydk8xK9lV8f69LpuEQRU6cvbrN1V+ugbYLJF
5vQ1FSKjP+ofmD4GY6INVJHNtLXjegP/Cow8Egnys+OwqUF0LeLTfCZt+syoYvnMURsrMngS2YRb
EivfodIkQnc9qY8kEO+l6jOBfski6GeCx9XUZ5H3uLkHY0wCEWVUfK3nfTEdcL4G9Gl4S/Tmoirf
Rl7iY9J6A7jK0J+lB1ZPksc8sbN91xGC8KMzs8C20aUJovGHjXFOTmEjKCMNcAjsFW1AbuoPapzU
A5FPBqY6hrb1qt7VB+hJxNKoFHT4/VcV38MnMOgyjtVdgmy9mvB1lfv+G9S9fTbdz7Y2igLIy0iC
lKe2uIl6ZquKjLOFuE7OiKfGMxJsm6tuWJxqT05Gd+wNpXw0LO4kox/hmih0c6TYYEPk2tM5P6dE
ZBMbZs82s9r67pfJRyTsSkLUA9FZ+BwNfoBZuoeqcsJB0Hkz315UuYaG/RnPXAla7DNbQHTTUNtI
A84XBoY/TxPwQ3UX8wAH1DxzykcBeFniqkKo48UNc7nHhTsx3InhF0D/PzGC5wj7G8V9qLw5QfS3
8bWE7zZ8p/4lpHtNXSpx5AiqdcRwu4w+R9SeXl/AoZJGPLLWOFLOCY79AUlDNmjlqdfsRgEbFxBx
XJZdd256msGa5f4WIB1SjZvZtkDzWDGFWT3fkm+WZ1ekpDR6XFygWA1LfIIuf8SdORGk3JVZI+q9
M3ZD36o/x4i7FQEKgtCwqrzIkiXt8XLh8gSxFVf776xwMYyt8Yd5H+48VZKW4a/vy8vucmjdf8+F
fbQH7ezsW96eggkEQ+wc+aN+0SxPOAsJuBKR6m+ztkipCI9G2rfGFHHeoGdwhTtgu76RxmyM0uVx
noIqLy3Z2CthKNtert20vY5GSGX2/36ZygXs/mQTQ4nPJ9jaxqoMK7tOucWaQ3EqcrUSDMtABXtm
EW2jyeckKZZ3Ts2JH46Glc4PaOWzX8qJg0aWPLuId7Et2WN8OF0v8TYNMfGVI5GWG/9kprgtJ1je
jAdjWd1RdX3kzpQTq3DNIUHBUjbHR3QT0aBrIMzkrOHh4GhKdA/MsWByg8pA22knIEE+Kwh698v1
wiGgBJ7spAyoWhF2UJY338qbhDG+2UmSBwioW0Ybz4BDS/Gb2uj7fgj6L4R00jAEy/osbOOSoggz
KMWg+y6ftlZNIbdI032CueH9v8ZAKW1QdxbTEo+DgxP+JD5DoEGqTL4VpjkH/cYcu5WzpUG3kp4g
xoR83sOzqCGwRRiWUJIuw6sX4RXdQUaHV/AF0RCKMU0uZnjZ+xZkkJYIoEQ56beQMUFnKoEAbXCa
iMLQs5nJI0FqXsJQZ9YgllnvlT7y6mx/FUM7N4QgAdhp3f7iC09YZVJwzwwwQJ+9PzUlUKGkIX8p
aKB0WNgDFC0YzHCyMLsqY2gzghEpX53JRcIXrAt+rAkQwXESa39EYUM2XMvj4UBB4cSUgIdibCxJ
59JolcnXziuNmBPKlio6ae5tb4zAG1SHyFZxVk2lZpgwgFjovJKcYYOHFuAX4mjH7iipthmuHZRO
Pgi0RRe89yWGdhoWadhE+/ZoIMo/OeaeDSpstQd6xBmb99b1T9qKUwYM95WY7I+Awbz+LmXvj1b+
vD3fVacxZxQ9P/bO+aoN5E43d+RvpYjFt5N2oiv/k01QT3GsYv+ZLIt2zry2y8Lww+quYMzyaFC5
qQlwHsNZMMXhjI8DJY5lHEGQnXjol/cRQnwp/TKDJFzVcD1YoN6qOtcg+SMjm5EHYeQPx3TYEF6G
t6uUjj8fzzbdfMNoC8nsIOK+b+NMI/IBGWWgiy17YiAkQgClynqEWU/Wq0WpxXacuKkHngS5IPna
347V8UlI9mfG/xzYtxft8FXVRjoEt1qLv0/Fad9+8jNHJlns0dQ7FxVUYugO4K2+ahUpGWZKpp/A
4aIN7T85Rs/uBdT6YGLWitXaGl2j6q740mdAMeBhpP/jxO/cI3V1KLp6Kwsfs85Djlb9Do7k/ecC
qb2zpxkG/Vjn8dn/A3O7VK6RCMNYsqnvTI9gzXVy/qE2soGDQzfUK2ju3pzB4WgggI03YfAKo6fA
PmEJn78r38cn+6OalKHY9imYhcokVeu7gaZt3HQwA5hpOycZsI3KYki3RHXBLsgwVmBCUhqNvmb8
XXhXU3pMrqwiew5i0QTL65lj2fQK+F/JQ13pRTLbUj+Pqp5aQ3JO1im38X6XrF14uBeFU0Oq1hIY
mtXLG7i5DMlLsZ4nbvTswkVdwJYhi+Cn14bAyvTkn5O846J75CJMil9rjrrV3LYOBs3aEdNIqr9i
O41EAihLtE2J7Y7qbzYdFP+fOdf+qd/dWN57Eb9+ot+m/n/in8v0dD3BXoUP4CO6PF+chA5W5Xwf
Zlblco0kyCzuCEZ/s5crN5rYkhw6WK2np16yslYQtI/DSQpkY3EYGXvN01IOSE4IyLRJ3Wib3yZl
y65j5/Mq8v7DjlXByBlLv1BulD1/jHIemmHaSs4WEbICwXiE3Mkt8PcVg2l5GCGUe8IbShHirjig
oWCe1tTiLuscxcF0AZFrh/4Lgainpj3460y8+ZT4NvrQKhuG1zZpvXRdUvSjbfFUnBp1m71fxTNl
j9r5PfMzuqAFzhjXxOEE4dBv2/NQNzyfw/BfYqEVTD9ooMHYOVy21wBnJXn9uWIQiKslLKkWs+B0
EuNUSqfIat2YaBFDdCmbgyBmFK91rD0uPdbw+B4R1rLDemyIY1FWiuiI0hXvElfTrEiMChKbZg+h
nNeLTCJ8kLtjjpD2QnV9f0EfL8b3pNMTwNjaNuv7vy3a5/fnpTGMGhROKFKQWPWUw3bvgRB7JVc6
AB5CPifBzqwjn61sBxQYEsTxpAgAcvUD3SHHKqP2SlFYeV36u4JNDvaYnvuWbAOnzKd1Myle0fqO
FTB1f6suUeHF0pyRUfbSmKmuVik+ln8H3l3lllFbtFhwx/VrOxSelpTkCk8J/iaF0bp0eafAn6CZ
tvzGJck4/5gi0E3qas8E8ID+F27T4zthb80+7jTyK1jCnMC71zX3NyX8qGhlfaoV3kn+dXV3bItM
koAMulnXLXUBib8PPpO0bwZlwZbuoGVTTQ9ZkoPU18QCsxKbM+1X9Zy1AyAIKAuzYcAk8q8TOjYt
Xa/pd2fbH1hQVJem387pNzqE//BOMJxtSPTryVpamRpq/dSwvxSVVbA2zIMKV/7enJPD1o5OFyAT
we1ME2alkP6fzLK8wS8pPw95uWuZaZkEnxc0JEcAFgp8MJLffeHls3OBhff4621zYG7wkfq0GDhn
CNAgABXMbxdi+ACe9/ykcqnyNZ5Mf/UrONbYfQO3sNYpPrdzzIZJUYM80nwW8di+Hy97uS5LhMLA
53UocriSJznt1Z/Laddnd84wzWmtKa4Z8jZmjP3WY76q6VshB6p31F8ISwndBI7OLHwcpsDR5ynU
0yEmoTJX/lyzuCP2RqkElS3AJFWR0dxrEj0q5u58XLYS3rKATPbFwIJnbGt33liHxOuauCbBWwoo
/VRKs5Hjg7s7Wm3Fh2RGu8tEtDiBn7ukUnL3EVeSUZkiG1gAHIZvgqnqX2CgTk3z7AXk4q6Fayzj
3v5lf6TlSCaGIjTVrteIpWocefHkHKoLk3WXUVwaDw5c1EIv6U3fi9tQ8FHF3AtIYriww4NVbl0N
kjMya6M1QbI2ocJ91DXJpg3/lma9Z0IJJzkFR1n6WzrEAfX/IArXyC2IQxzq2yQE7aPDkR01o9T8
2TKzZOHbo3Nf6zgLjoxwSjXsp+9Mo9u9eommSftkRNpSlPbATfV5dIVQ4IKIS1q0QOoi9C35IGMV
oCdJaepJixEtgGmx7SraKBWuXsmuhwrnzP5Ttw/OMnW7Uko4r/qZ0waJMHuJ0YIEqx+2aapt7HgW
TgoUvHq0V/U98mcA95X6SLxUh+m/FGVaWKKTxNB9F98YLqT3Vgs9dOc4AglnVjAM2pktLQtmgkxf
D1PX88CIFs15cbmsFUxJsDJZuSpAVsFxPR46Z0J6X7zANMrmhDg8//vAlvRJDWJOsWRJab4uzi/z
opc8oQcLMevoQjV4kvzZTi2WeSIMPgirIokagH43suzp0h8F3zY8ctfWm47K/JcnUcO6OXKtoBZo
eI9bzCHq/pUHpvz3Tp5CN8v/ZJaOrL1lAN3ywgPK7z2V/T5QiV7zla8mpS/O8NeqxPZ6zLGDKk0K
Mpb5mDmq/khT8c1+AEC++7ymZZ1MFHBG46/JJe5TF/pDEsFIkhC7mHHM17LxDTWc+pKg/pcPZUvR
1CaPShZuF4S9A+LyJneNKKr0c0g4nZvdY3aVK0r6LOzxUECb25tsLfBfcdPjkolW0svEh30/V6sQ
2xalTlledEk11mdJt8V7hSSVcJbqyhlvrbhXXA57UrWHAYExWgKRK2qK1bnp5YW0gIfbDZJJ8W9O
R2/kcqPjVlcaVBSJHMT3AO1/uRiDFJWDQ8uBrgkxfatWMahefh6uhwA1rx4B5q6mpl61uILEsck7
y6yST61Oh+l9MwoI6JU8LFytjSOn3OCP1n1tManpvIb6gX7JQL4cvbea1jKTKDtrG2kZZ77FLBIN
Ed1z55CPh2ikHsj4tXz2GdxC1Aww2EXU3KWj7M5nWYrA3ZqADOEyOZXBAZm/k3mNy1ghOidFEbJv
fuLP9OufcuKvO5eW2N9p0u+WWWnQbLa65TDzRJwvxHqmP4okX4stDBHh414ob738jSWhTeVAB4wC
vxVUTdQDsKVHCPGSUbQqYf50ZqGKSDETAmLKx+PBpv0Gh5DFG0OzZ1xUEBLnaJk8hoEmPlenaNRQ
Lp/G7t416cbP1Lb0+EO40tfWNVVtSvLFZOMlHT6rX06jc3AfLondn2e/xVT302my8w9Rzv84TS8q
DR5Aqoar4IMLCk2adsv6Dq3OGG2wQbOq11xUkAHVeQB49gkNDEU4TXGa3JSNzXLhirNSKZFnISD+
Ek3lclHeghe9AcxAmg5znXEKe8yi81DXawClLnMcYxGL0FqYUqH+iWnrejU105vN/iqwzVwz7PgE
dCseZtWEQ9VON8Bjr/5W7O97lXcaXJ6JI8+KeeEJD91X7a/GmDqEahKjl7CO83FV+P7j9IOiaZSZ
xqKTQ5e2KO6H2MWEit5d8WAlS+C70yApwbKiJhjRN1dID55NyhGQHGi/hArhjRa/TM1UKF58ctLk
Qr94PVsbrFwcfMycntgtcVl/pBbufQ4LR0r2BsVySDec9iYz78q5ofBQWL+rgb2n3u/S3GkJ6i0f
Qm5e7tlMmt61OHOfPYedMhIXrp7+694RuADsi+OTTrGGyJw6ujjngnmt7c6RKVqPXObdkO/zp9vw
FGQNXKTQ/SIt6nuN20uGxYSlRMVYObM0JuWchSLWLtQuMkCaZeIi5WYPewvOCLmFDnTSFfEAb4VO
xxtE5ozloZQKa7At5seZDSn+ZEnAmUz4bvZZGVvK2RHSscK18IrgB88BxML/ovM7UIqlFh/zVH9u
zTdZrmHLrA/JQkueyY/d5m8FeUwzWWYI4m7xvi+XfZYxO7wIGIHJbhAsfkhiXtspFjbX31sbZ1aN
Yoa5jN1fiQoGzgiW94IzOhyfR2+IPvNb0x286YjS1oT/IZ7Caala83KjfyzXz3OCZSaVZXQZj4ve
wJHE9t0ROtw0XwKPmqpqvtt7uwcsBqNj1yaL+1rBhuGBHLnhjCagL/DM3rjHmUy61LfKyBgYKiFX
nvS7/K5kkwh/TtbB0in4U4o7Ti7kkrkmKgPRHKyf+eTFSbdhW6cs0hxMRC8a4e6D0vj1gD8ZMjPi
xEy8v3rdBxPL4EGPL/0Bq8VQ6RyrhTJXaPNVUoeJtuXXBGnqWJvG+1vE7VhkPNKKUA65Mcj4Ock5
6u1uGeuOKhpey37tTTPQ5EVgjgfNnXs22EUqRpORynMvGQPleCDiQpHV4pXfTrLlNIhs/Wp1xn7F
EN4J3g/oO22yi7wOMbm2kx62lqLA1hslG+vp7iHGx/93WS6U8FpCth3Z3TjiTRAFTcV+IfRq1rPi
9/EK5GlSCbNzGw3hIvbo3/2ECagSlEmMOlNk51OI3EYW2wE4KgIn70N1c8iFPQjq6TgUnlRvob4u
/23lVTUQW4HozvJW936IbRPWuUTYc7VKYCa+jkP0k+lEy4Xn6+p0pLfyISEKXNLdr5ClezoWxO04
0C2/Oheg+8abs1qgh5zZlpLY/CjbJ8Yb/Pv967dZN6hCQSMBzrKbt8EmPthGinLmbsY/0faYqO9k
YkPrgqHdKDlJ3bhUrKrU4E3htYQASg9+Ope8zVSt2Ts0NZbh4F7SEa3SIkW32+SPHOKqgr6cprH7
6bShWVqXZPAobyimYEV80vha2LI8yXGjyhVCcBLaRodjqUq6RH72Ig59RrhcVMbJ//WkFdFbSxRs
PXhyn7PjwCshMrOwtkhiLY3bCAgFSvSBdvY3uxTzOODxdIeSL/B6xRX1hMB8fdB6DpZf/GaA8eds
lxHlFH/0RyyrZIpgIq4LZEMMIcmceioBG2cNGpC5PXNZVPw7Pvp6GKw9iBCZHLV44le19j+rVBzZ
Xiyxet6kIIZd1waPRGzD2S+rWqrktyxRSoFUKLrAHSHIAWZo8HG2w9RluwLx7JhNaAWdYOIzaer3
KXAk9cBOq2YjH8HSYsG6arbr5/PCaU+EOIC2uhLeTx9o43I+JA1aLE+p46kLzClZD9K8yjaxj2ea
TEQkmy95P2QaR19DKo1DTKzaZA6Z0J+3Zm6n8jL9k0yjia2RfIT2dIRGGDGiWZAblUOXny0G+dL/
EpZc65zCTL7hc0LZHJH8LparQDrwdChhWe8O1b/hyHQqZYa4afCeALRu2/ksgI8vytoR0nB5XYds
HuVA9128qb7KrgrmYejJ74TRXEgXGrsRChdyO9PGUgKDfFemsd3uIi2gJEAX7reOG+4KBb5SQb2m
Lj/7auaRA51Q1eZMCau6iPdOC2AtgmNn2RGfUBxgAy4qUVPyKS5psxe2Fonnq43DSG9bEjE1M2oc
MKh28H71gZunwe+c7+DcwKl/SEDYPiRFGmsAeBju9uB1/13nJEmLOIxBdMvfo76NRJaxjZ2thtAU
URFapmJ/II+xdjxFsShJJLm/yB2IkU0+UXcNK8g6ToOIgklSo6DKl6e598orGQjzCcRR1GiPAkZk
YHzvCTxhBbC0aPaL6d5vEUmJIAiwOzjPJQ29/d3oqY+KsCX/jveKUyvk8W1/8EYM+DeM0c+8Uong
sNVV6MFmO9QVrAJuurnnscgpaCKRYlFi8t6VP1P+KUyAnO6h+R6jH7RgEUeHQQgMPcc7817xIjCz
ERcBRwaRiFamnt1qGQLtoxZnaoCU9utEPhsyBBlQQwYVzmman00dDW34K0S/Tx2JL/N6z47jp7Yg
mfooCBfaO2vyPwAzl7zKGxebAvaGOFzpb9Xy0ODKDjqkfskHIyLNU50TKFZvUmZyu+x+2Mh93c1y
+NjCS5QI71jZ90fyMjJz6zih1yAfEto/Y8CKBiRXtpW5Wud9Q59zww+akaQ8fH7azl5/aeiN2Ntu
3lQa/DZWwJJgR5xvV4u/ahx3looewEhO0LCWUs1ve1Hhsp5qbWFOfQJXunlWV3BEVvFI7noaixn0
MM1aHtdWG3ptJ5KDElto1HgxoBI50876RCVuhkMngDXW9IrjeZDOkr7+abpTy8SvR/BRo+0iktDr
mXv8A4+1a9QaRxzdBmmkiX0pgF2ssvTX34mPNCuU71GOl049cCqYGFKxL1zubHUlPuI8erM9+m1y
0NecEU312yL2J+wFTOlw169JddVcZGylAlaiUTHsUPPS7x9NMqURfYIlpt4pzQ/c5rZH8mdVsxB+
L/6gQ20NBNojNTC+2RSWZZbShK9oHNjddpWjHnv+pQModT1JdEBBwaZnenhfwNjUoDJnK0WvnUqw
B14UtC3mLHlxs34a6XspsJ6/SsMcFI2pphY07CsYCBcnqKaVEFwVOrJqs1PQESqv765i/Yw26hGU
1gBiOqFqOZtPEE5zZS0YnuuM3YDPN4yAHRRhsRUPm0rNcCOQZDR+x7fXc1RC+urz15bOycyK4u4G
QuZal0EgJarb29uzqSb23Xj5FaM5MHagBES3ziC+EKZfbd4KsBL3tYFi+kRyKHwhsCJ1wS+Ds8H9
Ci940BJ0FUjnrfh1eao5Ns8JL5TfqrSF0SKUdYxlQVRu8sDMNzHNT/KZKcuYZy0sZY3S+wJjBuCe
YWDENjatE/t09yygJk88wV53L+e7FgTiq3pJzjeQX2fPKEIq2+t9adqsaJFeZswJsLrVM2w+ATDi
OmU9C1ekjlB94EyO962u3m0h93cBuGHPCO4apGaq2XPTMfzzhzvM9g2BL+DxBgZN+ZFq6H7YP+5T
03WvCGgxkcK9S+L2T3JtGs0Ya8kTXBcVzS6Ip5T3wyw4E+PPF6uaKEWVDxiUxGLq3aBT3PxBDUh4
aUs3evC4XujbPJquK8WSPW8lhVsLMmYS1/MUjtiB3t+Aqf8z0lElpFlnv7KWhJkJI7w2c5K+iwG5
8DpHvL+j0+UT21/osaAsFJt1rdi9tsU+sF2fVzo4NtcU3wNR0rOlOhxgzNufMGMqQsAZQQQnf8w6
6xwyJ92n0rk0LActiAmy3Hg5g6/vhNbvuQd55Y5Z5Ija1NJdxA86zH3o8I4GuDCQfhBy9aeOOWsJ
9+8C6kqMdaPGN4QMzkdRuT0GBH2Rpoc6ByDx7imVPJusOoIsIzTEml40je2kf05/mkeB5Bz5B97g
Ap2GNKLbPoJVPBRNo8Hr2FuquZvkja78iWl6CoXhWFyW3isQUSSAYeB0cEKWmm033cr2MMW/+0wU
klPufdSa1i/MmntyRHu9Fsat/CLkG5eY6Iq/y5d/gUfkWwnD5Qit36sS2tiZS7KM1Pg1MEf2jBMY
+15Y7GQuSXvVwP/FNGRp5DxRHLnTcxasVMMcoE5rl7WIjTHLbcNKox7bQWVLZoxGSnfsCLkW9+ZL
HxPXBIySA46MMBZ0f02QK68ZZvd0daTXvBYW24hG6kq2ygh9zDrHRFM3PZJTEOcsmqPPJYQa9EIf
5cAMxvHdzTKAUP65nZZoabFgQ9HKzJ5XRuXXj9MzCpsNvYHNV9bXHz2HJpQzeN3mQOTTpnauo8wn
eMCIpzkkN4p9bOazAw5B61fYEBM1jqV5WFM6XrhAcUFvi1b8wZm7PXZjuVp4LSZTh0+ZYupzVVtx
kl6flEXQqXosGvDPFJyIiJILjyRfqIHqoB61zhfMmUgkLtFZp6e3NgZvAcIIexxZpWkO1mZxJ8qJ
cuCXWsH/DckAyIZVo0KnBEZ6u8XDT3VZHadk4FzuB8X0U8GI51Kl8VaIYt0RmqZNHebv6ZacE59U
I12sF5qYQKQHySaON26epFv5/A4Hldkg9eqFBWpRXyUtorR5aSZ0DiYGzB4LzkhBtrOUkBFIJcss
wI1H5r/itSSR/LyM54n6zNcO9lspqwWeuGG14QO/BXhEWaT/rKv/OWB8/l6APSYPpvKfDrldOQgK
dOwQgbwXv1Jo7S2JbxsRCX4wG1Vqdd2NY1nl7p8D2cif4Bm9Jr7ImHfUN2Rg8Ep71HodcRGxKPZZ
x3o06BzpQJXpGn2pQwlsghRlTYhJWM902fneJj/LpTvYuLhH0iepdE9OJvb0d0Iz6qTodNqzJa4A
3r6Ebq6En4SgmdffB/uD77zS107z1BEBQ80HJ4HY/uimPCUI2jo1vVzcGLKl4tCMiLeTBQZemm1Y
FzOQM8qU5Z2Y3c4KCucyRR3+ocQdhf45Bd+FhPqITODZ1kzYpMkZHqKR/1wMIcGYfyDpJJ0aJahN
37q+0P5tM3Zv1pdd9O2mAZZnwESR4/KehuT8USxpDo96WauZlQmJZ6/NI+mTs/hDLJYAQBO2HCUC
8V1zMx4tMrBNaZPpYT2+XKkm7ZznB0wH6oYlE4yQLe6KcJa7Wdc2AcgBxeg7GgvezZ5akhnTy0fq
aYug/4P5aQgx6NjQ0gRwCG1R3OAXnofRMYV/il9Wfs/iaFxQNqYqiPiXah+4CSQFtpCHCowfEXOp
2mFR1+K5yfbkzLES/83TaVs8AV2a2KWS+N+kojPweijQA8XTvoV2E94JDHejOCJdqbzAMjkTLeY3
X0Vu92E5GXumv0gDYP1wPL+CnTA0f8cWqN/YqbMtcLpGcqQDhblMbRTGR4pZLPUenPs29Quw2HtD
pnRs24I6anHTphfmb+wjL1OYwgT4nGUjGkr26aW6/xeg3wM8otC9wsyx1Tdont2QfjiN/KzP6VFw
T0Vjtmh/Dia4QB8eErjeM3ELlZfLMjyyTPEvdGMZ4vQxMjARIUK43c2tRuWXuFa/CWDnFdOdZgEB
ZjAjZ5IDLv4Tp8j7Y2KNefCbKk+mhW1HNby1Oe2y1MfQTx5+eQclZMpjDwBSAaxvuZAAvcTS33Ir
D/PnQjN9V19c4gkSBQZgw9CfcRr5eKPoi5J7CQ2lBnLuZ5ARDUaM5jf+gM5548lJ5i2rZcBe8ZIO
Ci7F4/6mRwnlYTQjEwBs47O3/MVwN/LHBq1EGrblMKxVZHaHYkMm5wyqLnDeim8ao9TFTmPzPAHe
1D3p0uc3R7BbuHl063WQwFMaYv8BVVYcrG9CIo5Cct1jmKshAd9d+gf2ry8QIrvD9Yd/0WCrW1DZ
nfVrHO3sV/vavhM4BFRUwLTyCzMFbBj58bTxWX4vS2lLsP8W/c/pDUq14ubsCRNBLCMF9jQtkIph
qEVgL0s9hG0auHpqXU6qj9Eh14NKg372AyTUFUv+ff4flSeHmg/ZCA9ucl0ZRFERaqbTtztUy8DS
hKBnq0UCFijWH73cVn9VmFO6/AHlkBqJyFOrYB+d/eKvYK/ofXgIytdqa65JoB0aWwG7n701dCnR
NOHBp8HzT1qPjq0kiXAr35EoKNV9yN4aPWbC2FeIoEtDJ1F34tiJHJuz5CjWuijvAz7/Ygl9lNNn
tJT6w/GxsUCvW15RVKfVUoUiIV+F+36+gkGDNY0efWpDwh2edSmp5SE+ACd+ybXKt/we3kJoCGH2
ZTsps57Ccf+pIgBHQfL1qSUdleogK5EqQOUQOLWJF9di1ClCNcK5Ln8kv8Ve4S0tb7yRKLP+LzxU
ZyX+K6dT7kZUuUgepyqjwrmh8bLeEiP7rdD8pwWnVviceqvyLS56mUQuT1ltHGcSH1Q+Grazk9OO
PXFMxKi3iW1ogDXffwmO0t0L4vha81Bi8NBAG40DFniRdXhM/waEYAu2Aj3XdDS91Lt4k7Mu9AEi
AJnypq1+8YTukkok+5nRa8nKsmDmeG01FtxsnlQ4RpkZLDw7qFxGgEuK06V+Tj+E85noZYgCbTAY
YJABlMEoc/Qd/NEGc/dtSvsfMzLRHl4/eHwV79N8zHZhwbw7RV6aXGP9wPKwywu24pRTdSlHSSdZ
LWWg//m8yjFyNji/LjWLv0bJQo8PMpqsjx8bPLJBAVoT3hdC7xNj27pXYs3MpnoMujvzjRVHLjkG
GXGbR+/EjZpG+tmwBvo1Ry6reCjTX+38a6CMFZwyBJZ7BdHvuWA4Im5lxWyRzHYM1dhbEDB+1nE4
x+HQ3n99yzGDnqjifMquUjYoPd07j2ozXyf4B3G4cFpKBFtW8vHMzUd16aR6uYV4qHJd2GhDwQR8
uX5Gxou+mvRFVP9jmbHl7IosgZgaNQtarieFWQC2BwydljUBJyZBMbnHQgUxJZDV/UYkmr5JyaUr
q2lyRLXEKXJiE9CZaTi5O5lpPZ4z1ZCDm6F9AcgPLpWjCWk7bU2RpfIk/EaErQsHBp+fTkOLXva+
zgSES0IzVtqdcpcCUc2VyT5XG1cYBEVqfRztjrI3NFTwv/YO3WHSsZYe710dxVjv1SHWIolhiX5X
h/OERECbV5xC2FCVOoVMvN52HWB7Hfqr18hSdhYW3/eq+f3Z4sxLCJVbPM37hl+FEuIeV314U3Ur
wt3/XvAfbaCYnVzS0zNyeQ3pQEG8200UXxbIZ8h3Zh04M0bYRzEXaz7RwYGlJfo/z6apJUzPBsOe
j/VrpbpKROs32S2X1GeFJacwfLmPtE2tgixYHeLtlJZk+K12qzSY41W6WBkhnuLtiSvpU7QI5cM8
VozioPhgmmiTbFuZNFvLqfwpOnvgbl5NUvj+ExmOPBqwl5Vpai1EJO+btiJ1rz2guUYlLUmQekbp
ryLLRgoHJQwxamNq5YosUoELifRmYXIfbbW8MvxAfaigQVunwNfDMeBjJyDmfn0wHSlmjdy9n8tP
BTPasBD2l5xrwXs1lJywc00oeuM8/5B99Oi7uONAN60zTjTRk0Gn0Bs36w3VCzRTMiHBbnxWL3UL
tXAMthcvUJbUz+7Ze1XLaYg3Ff2V+ewdY+mkDUpYCF9Mp9Wvqfb0ls4LaujHfwRHEESbg2iNuvsO
dilW+XxdwyqvBKV/9P28kjJsLs8di63TcElSpqndIwuNO2Rz1AsbZ5uCFJqgsGNXzWFKety2W5tD
iK8NpO/1FNRFlm4zr5MLTR/2fvuT0c9/jhEYfiiAyfFrTZBLNLr65qBSYTqSaLuXX+tmFAGEVEQN
c7pvEyOZvGpAi6jiw7IFch9llMElU9PiAxxJ70wSfByZNngFlbg20+YQXTWy8W29NpIGVBkWX71y
ERNgT+BII8PHepBZL7cEuOvhSSFXYiDYqoEn430tPwiE1A07UaKcVdD5zmjBFlj2jrPHhFwC3Z/M
BmF24poX/F7plgHehhoTvkUYKfiLvO09cQRbtldMyrR+Vq4fc4F7fhSizPlzkVVMP6UItHg2AnKD
rEP2JaFAjg1rlbbeB28rOtm0Tdd9s/Tl8DhnYroPWjfG9g/tKi9SnlYEUCxiY6RXLccNKYQ2SoWX
PkxnpAxJzg2T7utx9VdvVy3KFYiVrvFGSJMujs5CWAi/s2Rto1E7fNYXwfFN95neawP5BIfe3gxH
D7fZE531g6diOf0e8teD5mo0sbqlOc5N/6gL1cxqKFz6+g7f9l2iGBoXJH4fjqnb6BZr2K/5IioQ
qQdjf2jJrKoUgWqpYf5QvVCh7OxEnM9VjCcaShKmrZJ9skrsHBElb2cLo4MweSVYjupz20wmtD2Q
1lbB9FhSxPTY3NW7yVdWY65AwLnmkTKXKKE86vO0uGYCzgioB8Q7MGkxtkRxItU+6LkhqRbl5nzV
MYMN+6Xui1NsfMZGrzXTLRu0ChI8Ww84IcPENJT2ILPzNpBmOdarIz7tqjLEpw+gXfKr+43L2q2L
hMyzgZWsZZV58hCTUzLaD1UAReubfHu+WOfcI2rbLsOka61nWxk6BTxmQKTczJLg8jEavmJBHryB
64/mmzVuO69L+a8ZopEnV4GuIA+SlMMx/F5tkrxnJ//Iqg2D4pncqH6LqFAHjv8sRvGFY//7IzJA
T6GKx9qbN+rNO3/1KgvPmBDsJ+Rl8P/B5Z3UfA/ZPDR2pAmyaeibV76OgGjE4dKj6mTvEpykkTKe
6L8iQCB7KtB+mdGuvpFw7EQllBFtFS3CLH9n7N/tGnpXgUlF3PZafdKn77zxZWFc6IvLLvpRm/D0
MdzexzKp0/6OTYlVFN92sVF/OXa2krEnKdDHXAdsL4PR+lZVvWlLcyX8furdq80N9wX/x3szpS1K
KccrKN5mWOoqDeMhmDkOxSm2IzY2c4DkPiujKhH/MJoMP+Tb4vNrml9ou9BrEQ5dsSOzx32GR5rq
2FoSjLYZXdoIyS2y2vnWRgW++OAh0QwR2FgbAZRY9CcRjJ8PVCAyyZTJ+uo8Rt7ObPKiZj+ILULc
TOleUj49sthNv7Fx1dp1qPsp3qr7q+s5qsMEMdsjRQaoN1Wyn5Y+33TES3tZIkR1RWE6ZV0b2gKx
jzAIqVmbWtekzJAAHJxz1RhGRHGKg+uWPP3xVb4N9vUVwb74fotIZ175MUEpzH1kHNMuMwE2e/t7
60PWuCl8OUX1tr4FV0jMisE0srFOTZJGFBklm8AUf/o0yTxgCIWhMkuzasmOI/itw9na+x5C0Bl3
O4Jnjln0WLI9x+/pudjUeXg9H+wbs7+E4YrZqkeBlOjOwASB1HZk9oHIGJfbqH4ddQ0prs5//GLP
Jo6R1/IWv5EgahytmwIhjyKiAHquuHx076dPavyDWJPoADQqC6cn5rEz+Q/tqGGEZMEhCG4KOVSj
62zBwh5CoR9vMzweY/j/Yz36Z885Qdjnpv41PXOXdxvVuILHouNt7xv5C4DxAkF63d0lNZmCKzKx
WNj/qgqb2aJDxlHasQXORsoVgT18iFWRzOi8EtoEZ3XhFG1I9hTcrkS8J/KMSC7tZ+3QsiObAMzh
8Nv/y4jVHcS66ScEBSXxcpRhy26D+IEzMJ2rDOlIed6ZV3i5R5o47hiohXJtfABAb/hW2q98CGqv
2/K+VkZ8WZHKDihXNgFqCuaA6A3fMN4shhPa3rddGyFAAJKIVeK18YW2z5EkKb3mOQ/mdL1MLpsy
EBlfQC3hRc+W61bSyUUWyzbwduP3cFOJLn2JKj5Kr2kiSV3gsasDu06DMbvHlFw0LR6ie7Ee1gbQ
64TxeAnQ6qoC3/386wEGAUsxP2RXw8xdSWvK6euiQAvG790WnsXgkiy5U3RFnNrkYZrw3YIVPNGN
EkjixVifbM6BT8EqO42zmtKwWRiEtNwROMC+u3d3Myt5kip+GTB8VPZXby/n5feTssP0GCK0WcTY
htofJrKRCR10X3L1L5Hnz2EbnmXkwv9atLfaOPejf42F58OQyltp1NlYPApVY6WSyFnnTojNma/k
Hu1TXr5k4EMss+UoTGp2HYErNZFhaUb+m0jzTXr23jUDpsIudqKnn+k3XSFMhjl2uQHgwwrLvdQE
HDrQ8U2MkDXGxMH5UKpYYlgeMv+NK2BSeizYoaHuaPZnbnJDjkNotLsChtD+JZqJ7l2y9SBc9gzM
SnRyANPCyqfXDWfSXqe56eYJPCYZR0hsS1L0kqP0wSFRek8N+HnSFqFQWtyjbdH+5bv2jVGoojh3
+1h+OgLeK7mjzF3Y9++8a8saQ5TQs43042UWrmUcsP8WThFu0jYA9QIDV7DXLpV6F80zWRSsI1il
uMf+Ca+gcA/RvHVu8PhbMUlcb40wM6G9hksmaTv4viS6TocL2hffNjytAt05rLs3oyA7EL6/9huQ
wKF/BwDl2rdsR33+yABVqZeBCjHegHhY6gcl3rG5HiNQaxKUm16cIWpGi+VwCKg/sqqz/lQIPyAe
b/F4oKUn7gQ6WTta+ABRiW5xeCsOlvmwRYUVGdjT8U4jSzWaey0eYF7ywpHun9gJFhjvUDcyPw9l
TQq1PTXc9j32I+jeQP4urkLeyOyi2PJJzfv2EVHxbOY1/ez9/ilyQMjjGhBOIZgU343lDptR2ujk
BBGl6gktor0LVFODyP38pOrUbyiq/Lx7hKq9Huy3mc5IVpWYL2svSSMhvtKds8L5vyFHtI5eyO/Z
KNuWus+1a+ByEAy1f9x0GexbNnCYelTjU5CIipcp/1o+KPvF6t4PHRXWOqMaYnGRmoCr6i/Dqmyh
B1IVBQ9HsOoh+DoZIzpIfnfInMNkznmDGvmwzF9PylQPDWGVzgFxHnZtQoHE/6kIpq8/U0C/iW2I
2o7RnwQXfakP8Bh+/+dU83GmIBX07hFoxVaNkboMhC7XQ5W+I1RTuJMlcx1G5svhOW4lQq16Fmz2
6ZWKMQQsOLERn7LP3CFf/47WhY4OiHwxnWgsHg2ZSB8Mmxn+jqL0aWaExK8tms1Qfg6doOqKdkDt
TqRKO81pGrDR6PNqeitIoAJ6iNQe1u/9uiBdeLqEr9OK6SY5zZmbSWm7L4AZ2LcF2PJ4lns+oaL7
ltTLR6/qZ1B91zKGzCXUk+vY0ifxkPGFo9V51q5DSyX8oEjpR7kwF8AlLQOcQg5FICNDzXrwSmp4
uhAy8nXMD+BOLUA20hGyFRqJWHd/0CBFyNu8mXmBW7Yu+q7ZRI4aBE8vm+QXFLJXYmumAfhB0RP2
JKk7y1YX262yRP4+u8rdlP7KMCWp+kjSv7LSFXBjlHh93XtEhaX4NARfGmbSMxworKtOCwNYIRtq
BoqIJd/orBkyGmaQpNkUjHMqop+CW8rN7QU8Pyw4UxnaH5UeNGvqBqsWOpDCjxVXJV4BzwWzgCpi
fNnYRY/ISZ9vYNlBhgkoMLUfqyujJ5CtaQyPyE6T8+YPu5fxVsnxKZkxkRn+h+wu4o0Epjuiz96F
J4F614YFTUJNoUEyUEtSAEdmvLwSj9Rt03P7dzIyOCocbqDi3tQXz6Jx/ujL+BO1ibbE6KSMFmcU
uRkZbXRSoMyXt3UHhOGG/OpmeP3FdOYbakPHwsjUB6H7phjUF8yfuX5b/jIBxCg8HBVzIBhzH5WG
4Qxt4CFTdGS6Fw5F/sIAV1sdhC38mG11ayIrsz8+R/Axw7BkV66F30w5wJGFvVBEJ6XNv3iAv5cj
qh39xl92Bl4MWKZDa0CbcJ/Nbs414GcM10eQr7UihRyv1DDrTJdoMMdtZfyFNSIynOQTA/Ao8uEL
r9F6TScGFlnml/2JHcoCLFjYPfX7vVQxqv/2JlutE7CwvI9HdBKy9SNOVlkgrOZq+0FlJ2OVZGFw
DtffIXH4VbSWdoSDBCfFBNZk0PhlGLEIapd25/sIhkwsTZjbFuGshhg312QjRKM0LXmWp3qmnp7p
Syw4olRRJ64+mCv89iLz8r7Zb7eokucocMCO9yVrxgBQj+Nt9Di+b9XKqS1gEm12Z59r1xUCevhb
jOkUzZ7lMopX3yszgORvZHz3GoqB/cumewKAcW4/g58pMF/MQRu43EX58B0PBXt8hLtpyOgKs7sn
/7JPMDLf/FJ+OXfLq4GyDIsCBEujXNtPsWMSx0i3Nej4atlpE8LQSdxsTwbU0gSQbVlftNxH93p/
WKmuJQjmJm+9KBsOgX3iIFf1hixBrYMZd27Y+h0cL4OhBXthW0go8fscl3EuARyTQe+VFySdwsM0
4Z7K9xeU76krsVqcXhFcnPiuK60PHjEiUrPWS6Wh3ddOVgsy6vewHnF0d1BCE5sUEx6micp+LG9a
PYJpwNxKCpD/lnj/6XPADQnuS2bETY5COKfWXCttpSvE0itzh2tcScpsBzHhs/u7z9/ghT0na11Q
DyUjsekq1K6I7ZOs33MzpCZHRsng3aPO5FS8CDTJ5vGR1cPaaUdL6bexf9bvuftEtUObVbJb4hAa
B7RJXdZ1Kox1otvG13c5aZPWvw04rN8xH5KwIlGpn2BMhi0/mdOxXw3P+LRi/jzvU9m6fPilJ/Xf
wA5Ns4c4CVDSLO9Cxs68wJprGrcjLMN409z6xB08F65P/FbDavQVKadkRNfDzjnsRdNO8U8t9Vux
59P13/tBF6FcrfpuAqaRT2m1/VL5WHOyVrTsNboP7d/iyHR5Eh66k4csxaiN47ZNUaMiYJELWuwp
cxcIvelcXi82jls9OBMUkaTzk3A08tbnedPwUqkAicKhXYtNTPbpT8dFyQksBEpyuBJDEKg6n3AH
uHntifi8Fpcerf4kZBodl7DfKSS0YY21BzZyYGvzYQ45N2fuVk9ztWV7LxXw18mxo0FfZEdeApzb
w12sOGBBodANTkWCqCR6DPmZ+LwPkSBVLo8Om2DdQuLvRDf5YcFc+IAbBmF/TJqCELM2mkullMi1
hWinfvfw8sDetFO6fdLPfN/5UqbcR5cVYMGmTWrnRnnb94yTfWJy5CekWofSmizCusTZLWSvwN/z
8Iajrd1jVYJ4aAnc7/tMp8+jWzGvCTtw2tWJ487cIK83NoLOf+OM2eMKS+oH0VI8wSlmw7NNSwm9
18eB3ZATk2VgT55kLJMr5bF/wb0DKkVtNotsgA2IgcMDAgeDaEoZ0mlhXoY8Jvo5AfA91xF0zZoV
qm4VG659YQXcNwt4eCHc5VQcvcpHo9B4MRefQpoBrOdhKIN0g+smSbnbn4aYe37jsDUJPdBElHhx
8Lz9/C8eSoONUJVeb7atzAem/4O/yJnlRa0/M/sDN2fV9g0QoBCM/ojMYMpkT8YAJsrh6/8Wah0Z
1G57gh97lLR9vSaisZm5LWJxImAIeoboJTOGPLU/v+6cS3FVUgF48E9p5Fz8J84Bc+u4sqsAmljY
fW56W9n9+8sWpfti6I6FwxxWJIxKKmXGWJlRHFQtbd5/Ywc2Th37Yv0MHMmCiOUjvn25AHBFmUon
fzD7wUSuqUiqMaCQKiFvltO+XqbX8X/tHoTbbE/2YCNpkUO9cckmgkmkEQybUOUwGAjE6g94RJgp
XYthnwWClQD0HegrwrnzgZP3xCDT8krfu5xBQAcxzU0nqhNnGNbjhErYUusK9w+NTRgdVqvhC2bl
a8jNG3XNLUoSg6JwSczs9rJ8NWyKiSS5EWbEiNJYnDZZmO++ilORwQHs1yfvXXzDQ3JFCWEFO6/2
pj5SY/Xe7aH+XT4hJUAOnm8uGjcrMwVYMEw5d6s654xRRvyBeGrGwnti0PUnOiiFby3vxwgN0lSo
QrYbT0wlg+E1rX2lVXj+kn3/pVQ7OI1bfLhGvovsOr2r8XVPaiTQ+hwaqzwUE0np7zbBa62Y+To0
wlqboNNZbYTum2rO89iEtx9UA6W2CpoNd8gJMvIeG7DGI/xguUjWtSindhLt7iWa6i0QdgMyMybe
wxvchFhcbkOwkcmAYLr65pc0yy2u7r5gcco7dfzbsQTdgtwmXhEsSaIWkRzOMEB9vgtv3ISK0mRP
S5AWCJA/21wyeXlQtbvc71NlQpMKOsJYZhS3bxLf+OSR5fFflRWEnr6xlYjodQBPL7GOLUVoO2X/
8W+YQgBYbrElov9EhfjiK/KtfQLNkoSNeZYmvixeGekgc85wNN696qgLOJSdB9692K/JQp5xvDE5
3KoFe/EJidPflzRxZqpJz3g8Vi0JdnOzD68JRaGtTdp56VJK8d/CKcg2dzbC7TA4NtfEG1OlEnjg
wfZER033DdfYglQllo1LrKSha3bmF4jDDqYP/krD4NUvBGNRlnqTCg//XeOiLUOg1rwexiqXL8Z2
NuKarxoE3tJfKvh60rArDB7F/5ozMw3MG/bSteNOvLMr6647FRCuswcCi3ziTFOhd/7WmqtqWsQ5
7h9/uZUD5PpDOaQ4z0giNeMvuwqTP2kZ2mkH/Xn7qPDdeGezZvGZr0NFV0doAhyKtTzlvkP2eVpL
DlZPoBrXCgxumsWLGLzybOd6QolOFJ9RoDDFM92oelA1sKsn32CwieiG5WXywTzxkvt25x7CHL1/
CSW3/0jpmm7BsT3I7OEVBn/vZUBBJLdOvWSHRqzxg40ib68IbRhrYpF2B5lsWfSBEN6mQ9zefDeD
y9k2wIUJ3CJ8NDyB1NJ8SjUqkTopLqMEZ7bz9IWdlkbFsnCKLPFYCTcXJO6/hXTwPxJJc4K1kvFn
8i0/qdLvcvGwpT66XxqfoJW0W/PMqr6nkNrvgQvEqITATU53tedbXOWwo5qsJLbaBxNb/IlIaAmc
QS5B75DxVpt9HLsPA19ap9wBG8r9l0ZKonzv8LbCglF3Zwb+2t2oBobXwJl4wjcETnP92iZi43o+
znGwXo6392D8ufQGlbMSeSzo8YdAefnRepCLxc19kTP1zATWtnfkdFkMSaQS9i4viCx4z2+RGscA
ghwlsrqYNtBs5x+3jQ+eOJMCllKeYGwipDQlX3GlFACdshtgYxe+4oeIEsqf65qhufyukDztxxlm
CuwiqGrX6QtMwDVFxUD4tuXLV2c3QMG7Fo8GMIuUl2GoeBYo20yIfzulXqCpoenXyehFbBGVbDSR
AD1e7irqizoCeNnVbTfYVkTJD3krEW5dQiZy5AhyZF1MHa3usXEVzKNkyG8nKsQHTynVvNHtOM/N
P94TUdCUSUUGXZqjuRqNe4C7o6IARptDUTMporbDUZrNZxj8KtGkgQtAsG9763WjgoMCIohnGzSN
MeOG2cYP6fQuCPqnDzDPM/w4RnF9NQ3Zzt8LGFvCAwZIlMk34/c118SRbC9NXGFKU09ne2yQDBIc
kH6ZpT00DKm+s35aHIschAiOWepUmBt9fDAFB+3xGqZgViEtKu+lPG3Uj/4S57B1VigqRw21HpVB
1Cm3PQcGmDL1lk+GMjdNmPABZBNVf730qwPqhIDIV80DOFKne/Ui1N5j0cKkBFSc7CFas1YRiAei
TMxyBNJVzhwgYRHXqri+hWnpjg1tUAPoJl0KuN4yZJfujyXd1K2SF2CMl27DlPP+nw6EaqEGS1hg
XSOU5FSJgoknEztsd0QCZ5T2/hG0HL9WWTenYqN46H9kFTV6zMc4/EeTMQ+9z1x3+4zaYC7UQqA9
28aDyOiNkTVFGGl7C2vAthfqoDsmQ76wNrQ5M5W2RNrLoxwomC/JR3ltwNTM363Kd4mpX9PnLJFj
HEEAoADedJWfbulZtLXx+jnY3qgyhOJqRFjYCdSiDdkUzT0zkW+JlEGeorIkHZtb5oQuTNOm2Puz
YlM6apq8KkYWp4AXK2sqh96sV1n7tA2LSmv9HJF8noayI9wsT9bd7Fs1+c0t45feFaZWaOeDWK5G
7xMIxiWInUNPtSMGVrcTW6e1pS+kgGW9gkle3jGwqksVPXylBce6dOQTcNNWvKeFoNcjnMVGJ8TC
ElWW3OMlX+E1zEzVdnZDyyl+qmUtGc+bLbT9FGk5Wwc8d/uDU4nZjOhXABwDxvlzlq5vUsvqYdv7
twIkaVjOAL0KccrxG2nC5PIxHjujyxk3pvUmlc1xKJEFVWd7lEX1OMJOFwx8XPezBRhV0iYCIVS0
xyCXfEhGCY9CPoAt+C0KjihbjxuMVSNnPvtCXHVBPXamVQTyXT84mwR/vc1ExJx7aXhjwuAERl0f
rlTsH4x2liSv5C2uFRrXzuFyCC6IZlHS3JP4JxhvMXCFsCQaZzsWh43duvfHHq36k0atHhbcNtiL
ujr/ZB5Z1ZGFeWe1HxMxC06ET6IrGGtthoHlJALvU6o01A0JmYpHC4rPpj0dz6XUMzyWHOmM7YK/
4uLHohdQhAX78xg9XPGv+eZiAfTHod4zmAemeC3G7HZZjxAGhUyKM1L26AMLhZvnLldCYOatl+Sr
GqaAin1UCE2ttCdwMS1VJmXcwfcVO/Ma/Ouo+5bKUwuxZp2AiYHv3dSoMA1Hxo4z0YnnCpjKmUSV
mgdnzqAnvinUdYNnluc7Cm1dYEl5oj4RbyBlzkvlSsZKfIUhjABTGN4zMfZXRdm1WRrgvOoA+vvk
1AQNXrzMOK7Gms2cw4Jw+USLDrvfIFO2eOfqh1hWjiqdrai4W2hiqo+HYGBsUlLD0b7WIZHOu760
c7Oo96NuZmhUYF31kWK7wfHXWGvrY7zI8+jLxWOYBf6gGVXMDaVbOukcXyFmM/AzfERCApDvoMB6
47kWQICrUr42pJyzvtixJSTmbyIFPTs8m7k8dXvNhvi5PwfxvsiYq30LU4/mYwLUfBMNoeCYnT/3
KTCO+QIkG8B4XZhrubqRs+Yz1xe8ki6zV8yQcAQW6P6uY8MSLhb2lvjlxYjzIY470zvRIqmBDNpB
iW5P1WIQS7iA/rVzSDJDWUBp2VX9mH6LuHNXY9StK0kgiW2cq5eAvb8gvkUDxwvVLOxqULCoC3wB
yHkEpArnCMKB/hg5cALyNXhzWvAUW0T/DkjJcGuPrKUrIqA/IZFS7Q4bR6eBtc9qaRg4OT52t3dr
iZipffRzfQLMJjxiyMeYuOy3iMsC87BYky6J+T5n37k0ZFTQ2P2MOIYkBbDhORG5NBNw/Gg8abX1
ryT4CkuX1ZkzQEp57W3AbEbeEwbD1BcyxqYkvIbZ0zRZ3CAkbHLoc5wKeB8mR5xTO28JKi2Tf3ui
9QqX95Yj6Gc24mgeljBm+uCrx5DPGCI9h6a/S7O12QTaDa5VEe1Ne4KoxEwVUOWD7O7h7ln3EEot
UiUKXzAHF5Bh09F8m0sDn05Qzf7w0jarUTUFKb3FJHBaXVKeBt8bUJjDo91V1MdNKqFBsTv9WEHQ
rtn+vTcOAtw9udqJHpAiiqX1E6hqAtxkVM3P/NsBet+iHDYoDeVBeK6CxQsEwsFsmkwo7STWg5JM
dkmJb1SGXLigyTn69dSbLm3BTP7CMY9A1Wi9c3WMWZo/SGihllpcVXyZ1USjGbsUpeQyoJ2hVyCG
5svcuNHI5SJ/ugDRjA574ySBY6M17N8CbM9JA9Os0hn7xAtEHx1g9UBuVgfB9PgWJ107wJbT2BpI
IiK+SFcJ3RagtcUBezSOtGvcQVTB3lPU5ZAaEPsTsKQ1fENShr7OYQprpAq3XBc8JXOY0ytAWtdk
z1GpWY6r3m8SCzef+hkeJcBgretJ2lyGbwzKmvAyJyCWfHeDqX/IaebcdBi3KkDpfGz9YgrVIgSv
UHY/mDChwrmn7rmUJHK19Pm1HMKqVlKoYso9kxpWd4oTYcXytWX1YO+We5Egm07TvDegJm0JkOP7
UIKGxr+waUWHkwl4fYRfHO5v3YiDsRFYRYHb0SeGXwF+FJEuWJ/Flx6+foQUDgGn3RMj7aGVek+2
JmDoMI+z6IgAch5RWsP4sFK3Cm0XFqTR7g7/ZCpn9a/eW1dqkdTMBgXJUem/se60aZ4SKNw+m8Ym
KnLGwZMzqVDRZ28RhCe9Pgc2/ajtMBmWhorgB4MoYejPBdnAOAzY5E/gc4l6e9E6qJMPIGA76Nx+
CEkSo+7Wintm5tRn5OlL/7+62m/LQnOiWnqb3Vw/PqonHkg41NYfW27+38fV7AG1h3NTn4rX22qa
ipYg5odCR4MIAcZyo3qWFUj7nnYW+TY1wh8z8BnEaTak/k/9Fod2FHWF6M83PWnyF1NS29yCHp69
hlx58dWpsSQSuKXHm70xhPFmr7lkfeYDmruOGVPBg7jV+BILX2wL1MUALEE6mtHLFBUlgnb76i6f
ORacUiLmzYfPA9/Qw2zxPDLHPqc75C6hHlNDenVJxJoyWADzwVX7uO0yXWqK1+El3VoyE//732LP
Hb5KOmHgyPMPTA3u2Rf4abs/q3eAca111/y3kOQdfnNw5c5YR8cBjFAVZ9Zd6eyrb+ZumDjuvrwh
o+oQSpXOAxb0chvvn2MfH0soeqa3Fmpj0RZmgSknMBGC7zIjBC3J8EXfnpJWjVkreLMktZr6OREc
Jk0xpHi5x546Mnl8U0m8bKn6gYpsyI+xPUejsNUDSrBgPPR/8E5R67JHTii1NatFSbJPKV1SvLmQ
xzH7CSbWkQY6S4bPLVAlTgAudE3JhOwivpbs60I8M0cuqbdPPoj0W5stRbC1NvtTdwfsSbLNvsIQ
5xnD0wwtr5s3FwVbWqSUJBRzbH1Etw05rWpUTzaA0r30pF64okb9lOYU/iTj24hIJEMzQ4EEbltA
B/pWFhoaE71PYQ0WZ1EUl7xTDwWhmXCaN24nQHuAKJrpbeuI1y4ifuJaXeeOCaaEr/A6635ZHC6S
eCL9ZgZkzshE+6EoRf6gTHoEMuLVKZBAV7qv+T6LjrF6hGmLrfYKdcCqBolbzY/v4HUnqc64ZhrM
M+CllMI8KgfPa1Wlne1B/gpWIpwLZFAyRQNXqFO7lUSD8Z8OTNuPaMQY0ySMAJEeBZ1ram/Ezt8f
cUGRDwo990JizQb9oVUbodHkMuUXAZUdGMt6yF3no9FW3h/Qkr7cjGjtgn0gSmm2TL9KFZN+CDLS
6UWWHQUoWKYOS12n3Z+Lu2w5icv08LsRY2zCblD9UiHiHXaxnSbZObXIQuIFAXGNpsducRYzSDRk
v8mDuHadjHTxT3UEIhSeiQTSxhneB1Sf4qVjTrQM2t9vLKu2RF6SvV1nS+BMgovGWE8PJUK/TyOT
3+IN+l631pSMfHe6Lu4NcOQcpUcLxCxYIY86EP1HrU6zcgqS4DYdiUSbvX9HdiMPfK/09Aa5nps4
AZ3dFiAAY5aFLGWcZeB0LHaN8ifoi0ZFr14lV0IfBpbcjsj0xvZp3+TCRA1OukFKKM7uFzZ4WIBH
zLV1t7Mr75SQQWxPHlZYzIl7nvfpeQIs5oUPf2RvybPgshcJ2lLmBqnDUh8dr/TA1IP8X7vjXjqY
kjp7la+AFEUOW/mYMxifkPj1W0HaG8UgKLnbri9JJpALG3WMNeFZXxK1okTYSgLChoHdkSGoMnHr
oc/A9jQmrn5RjccUgTNPvz2cqZUM3YUh/OXgSVibsU+HBNFbdEUrdHuKe+5+sfTSnRnsEFFuV+8x
yuVBejN55NKhQXP7iM4AoQkEm3N9b5Zdm03nLrohzvrqrAm6+lS01LxSRnsuXK8MALwQwwYLJuwX
7ItLELtFNEMnJI4EZsB01mhXwrMeM5tnzkEalrH4oJWr+p5Ohyqy6zzsY2d4UmxhndxIVordGwZc
O27cXyviO9xK2D26OwFd1DGNqSuUr+p955O4a2kbtj1u+P9/NVzr8lKTgggA7ulVHC6Yd01Yz5je
ysvA1/ZcezL2sCs2Xl1v1XQq5l5RbzuVdEvN6PgihMDowgmuHLXm8ABufuLxwF6AUOJXtdIFKBtD
GOEj/eXxn25be8z1NgicMW1e5BdzF6mET5/i28XIhbPZ2A0fVQp1/uh1CpW0RS8otzpRMdwMAM5r
iA2/iL2VI5u5EDQdSEb1XNfT93JEJ4xEajUelvv03Nd0EnoPW26qJ4yWtqSS0E8X5D/msNqLz15W
4xzf+wiTTuZe22/1O6j0I0UW+r/VKxN/WPO+7qaORu5Egnnk5RqKGHZJK7hayrv/t+mjHWBQrsBj
ccKJ3CV8BznYj6OQTcmvYvDqCGv6V5E0t4bJQVwujVM+Zr70+tCB3ythWDmCkyNOTM7cHDcRAA3y
t6uOXQAe79QYjs8TYfZ+PLui5yQaeLG0bHQphM0wd1kmj36SlA92SG2nNdJLqq5SMu7rx/28Wvwl
lTW7kCD/hgwHtciswdFT+wL0MZJ9BCLWYmVZlvvxedVjjT9Ct+a2rMtSMBsdYFPZr0VeYWJIxtqe
SyD682RaV27M7JPzr9R2nIS090dl0ifoGvn7ldfHgYO8quSaKRqFRc+K0kEvm5o5zORBblrAj215
2l5GHRWlfWhSdZv6N+8LLc38VKYBhKwSbg2AGQOIfhnZDfFcN8JvJdMN6eJKfaopj3/0I2M+hW9J
bT5B5aNHCFOiBoiyesiLV67ws3T8+Lvbg8v4SEqKd7hv2TYYO8sj/dIwNmSzdMQtyNayNDb7xZH8
xlTlYJNzTUl0Y8CtJUWrj4D7zokbiwMbUdzTAt6SIOI2Wz+eblNEl+s14n+EJ2QraNyfmPyhxxIH
OCFjko+AVNuoxEuL5wKHF3h6KOEY6LXu8NWX3XaX7WE2a3x7Q/LTnBZ+E/a5eEfCO/wx0woOdXcR
cjhU+co2bOJQ9xoLffKnbS6fIlO6eTkUvlQrlEqsECPCTicCA4jKrax1JCkKU/wXxo+u69VrHaXZ
EggdtuwLXbUnvVDk7RVbmbX/I6gdg/C5eMDl8AY3UDDlA810FrxK45K033PI8O6aNYXxhhbWBQj9
x8lA93OeYRHQyEs/OHuXXGQhIz154My43NDnclCum7WsGIZiZuDDlmo2ceSFoEbn4esnt0IokqRy
vxl7Zivkbyway4aGFWwicQit6UK2NJEQF+x4KpPJibWw4s/eRumE95JBjkx4XU4gfvGO8m2o48fq
www/ss1XvhWRHG5uyJPok5nAc37R/MhL6vVRoAo5ZXS4e4G6kOj4S8vWD90Yy4pXQdtONX4M787n
CYZYJd4ey19Wk60K7WGkbBJXJ7A6KQb3ns/pdbuu/R9jUZYR+4rrgbWV8dM6hArRoCaJPb4wY35W
kJcpHvVGhS3Er7pLTM/yoiuEWMzJXX5rnzGhHkdWG0QZimwCJscgKerzRfy6cFL6eFZ2aWAfqhp2
yObwldjnyeOZT+v3OMEc4/4JR03ZKAzVaagiGOL1Pa6SRgADHH416D3Sfhb9N8alZwpUWmiO7wlH
5+PKYDpczSbRZoY6eY6LQGaehagVBAdsVwI6nzlyKTfcxGY8rMWa2iRGQxytzicBEbp+7OqR5kp4
H6nemq9nVMWFwBNIkio5Z+R+pjkcdUj8I5LWqW67E3oPBebtbq1UiB4Ud9xhbCfJcJuYzahnx5PF
S1pcRv40SE4kkJO1kefHip+cRoVuk1E4ctSlLP7DRfjeX2r2hbelsT8ZM7cCyaOiBcodrBIBf38i
uv+DeGVpI568IXPJW1j5Bsntgr1grtk6IJJU1mEPJJhvCexI3HcPY7L/1QhkqHOQYeHJb5gqBAr5
dYaAjOXVaeG/mvwxCZ4uvu5m0984K+cijbflsSYAzPuDysb9HX1FQgF7LB8TcilL41RxB4pBakDd
tv0EDy5dq/+ToEBJsW+/mJIm+4vvGhE7QOMhT4+8gPjAVncVfxgqYbVkHKp5AH6dmCi/bDqLor2X
8TyU2Rcg0oczWethBtXK3jCAZjzF3h5HG19oy1d9aFfhJMy5RG0dNhyeieBX/HA3wYEMhW8jRSga
zmvz+YiSeiv3vCpUn1Y0fzfLQD/C7Ge5BaP0Qfr7kxAcktDT5KJWfxbM9RVJY6PjY5pg2+WhUrgK
G2pvtM5HhwdEDpPEcciqcwnB8ZPsIhBCN8rjs063CSoBqWbcJewHBD9QEm5gEbuCEL3xbKRqhnJy
vBTBQy7q8qjFdF9xS6eoYVET5ugSEEDvVz2YXZ1uWxbQTmCGI+ptU9x3JgbfQxJhd6ZkKy/k2hUW
ubeMzG2VvlS69cT2XCEWv+ux0GbOvLaf+j49tqNnnjJ68l+kD0wWJoH/gP7fAZztfpE+9Cc0Est4
ADMTqfdTvb++fyBDxercUlBkYRafk5aINDWsPzAILpRo5N6pVlzcQDbkr/aK5A+QIJqmD+O+RIa1
gmroOFmXnDmRqmdFAQ8iImIeY2PpxTxABVcumGiH9kfyctBudHMJNN6BGC2OshIX5nuuEeihXBz8
on49DdpW68mm9eqOhHTrUgeMjL211W5PLLcBnrq9zcujLiEkSdO8eg4J4e5EWfwZL6+0Zck9Q1bE
1WK4+BU5o/pSF4rcA+jeA6InPs2GIJpe0VB6C59EJVtNzhL9hkgen4gjtpc87EBlGaxK4pOeKDun
7v5K4OMQJihVh98eNt2pol7vO1nPKBS2nPhNpNpXHmrqaX8eg1bA0FKDJMvR/Vd0RfhHXReWfXCh
jx21zv6brpD5lZEi33uDjYJolecvL7dtoG6VGTyxuwMo93Bgf4JkRbTeKORaxeHLFJZmMNoJGgjB
VSEmOdyAWZFZ39rEF8ZXKgNC38qHuUMcm/s+bxAsupAnBJST/I8mBTb+4ns23NepdF9OThbk64Ia
icBbTM2rI5XlQjzcpvm8ijQN6kjnflSDyz7PuxpTqpY2oXGt7it4o/Ptzl8VE0hy/Pw4oVgiSvTW
srAmdTCri08x6OCrVAww0wccK6fdAAwP3rJT3LSmCJzkY0BNaZd0HDUJ5ScB7iX0FIhT8If1cths
YFv9KO2Iyxvgqkd2MXYD/zbYox4y3oZT0W/cqN1o+5PA43eOUJZR8y7MAkYZJj9FbpJEjtu/9c/y
ut2I6ctpNMYIJO4A2abvMFgjantX6DFvk4IWUiXp32duLQG5IocQLeAu+N6AU2XGpP5qzG4czwPT
oZBncdhBdEOxywDD04lKkM9l5GP22QBuCvZgQnk26DM2gkmIuhMGeGOnqwCJW2qBJK9qtV11CN+8
wOoMX9lSEHlJd1eHTQeAIDnOfOKXPJdj/RbUoslkz6AZoDXF5gi/FDDXTz4GMP++VxIWodAhHXBh
PXWb0iIqwUhVVldnSAHB9Qz456dm7GJJhAy/vbwjrkoKoNVGFfvqsqzy72b5CB36BRXwd7D2AoWT
UJVi5UodCxwv68jm+g2vSGGVPRl3WRIay1g32eyj4PjN1nll3mpO6IJuKH4PDlwplwmskPWlXHlk
F2vDvKD5MRHe9g2uR0eVuHPRXjvpnj5WBrvbSS63v3f8PB//oELLTY0j4lfD7GpM/BFBQGz2sw62
pkXUXrEKIYu/O6l7H8QuMQ+9SwhbV4TC/eGneq1WY/YvbhrL5acs4ZIz0xDDhC1CipoYdKSW0JD4
CLQAbaAQfMoyRCLc4r8WQBErf+YQuYnjJfBC1w6EwnZdwaOYhfUze8qJtMq91PrK5PtzWxx6Vw2v
AIFmYBH/HCgf+MWhK45MgOoahm/71ngUDiGxvqlk/69Wly6WwGbS6QbvTs7J981BCiKHim+8q089
hMOGv/o4Gg6DTxxXvv8ugPKZiAB/s6mYP7Y7Mbcwszv/KK/XBHZ3UTgGNdIZB6XSEospHmAlODWk
71keRaT6ZFfqhlnCwaNiKlbCm7PLnPcJozHwjGad8lH2qWcDGVhrjeNd6hSt/pwexrNS3yL3B6NF
efSXpyc3W3I56TLOovMtIkcWzaPjBfZNGwia04QJdOtX/KusxBAnhAMTlifIO6IzslR72RmwxUpk
6y/gC7gptFKQkqRmE+e3wtz4cEwvdn6Yq+1jk21KnyoTAyI8RHllogxftxDTuY5bZbx+Inm5NEol
kKqho4AxSd+XKjpT0b2MJYsugObIqyzgZUCGM5DdPeUOss0nMP6zp5iAmDzAGaCpYQ56ZuqDJW/P
n/+y58bTw/oNIksVEs7wOmAYfoWLhWuwR1kqGmzCoTVGNnrSaJrODFTUSGDJ8H5hVmJhr7Vq1VTh
JjbQ8qnI3UcGYmFVpolZe9fssgxcclCgC+HgLMcxBYoURKTtALQTkxQXpCwi65MD8B+/jqDRRwQf
zv98Z7HoyPNA8sd7Yh7ckae06P0riBpxDqlw+YF1kGPjmyZ/oJ+zW/r7IEWs7kdI7mVSGDcIQTTM
5Toyp3uzRj55Rb1Q8EN0rq3puW6kkqLsxl4H1zolJVAOeekj999OAUt9l5fXOjqkvLMKCvhwlmKB
TJRRWu5ygsEIXnpuD1mlFnwtF0WudgtdvZmFBz1XkW7EdlMjwsdBQSLUVzyT0q5YKYZ/D4UNJ0Cq
rG2IFgl8TDVwdB4/2o92FhU0ZlMKdESCcpZXvzE2s4rnMvRU3RXB3muOxGcrD3IeIG5iHTzLoUKu
mYWKxKn7+a1X6/pSlcg42PKHbrWrNuPbQWwl0EBjVnRQqrRvZ2kGSyrS1D7n3Bpr6tLatwEQRfXP
eZzuFY/Hr51Ul7wfgh44dFkxui+36gpqIpqq6lhcKOkcQtDgIBgPheGSa8M3L/1Vcsj2iFULq/cM
geliVpif/Zh/fmh3XB0+rLlD/0W2rnvr/9DrCOff2ZwVsLVhGZ4f+z9kQS1/31fOxkp7N09PREhW
jN2xETeSGJtiDwYV+0LLvizFzU5Aw9sLtjSONRXalZW9/SMLDH99ZCEP0mvM0Etf6NTOirR2r0h7
WnjnoqWLES8SIci/F9YgLe977oBR5aliWQM98SlXuywltaYpe3hXky3H5vsecNXxfELyO7bKCJuB
ljY8L0LSQJW8gsnuHC5Mfnn8F4IHEy7tCXIKtq/eR2o7hdI9+oIwKE3DP1iRuIbywYJZQiXnSX99
Frtz5ZKAQIxAzwzsiEoCL9K7XNvq7xL2E8kY6EULMrNS+Ij9aBV61JbyzBIztp0mI8EFY1EJLcoS
ojGCPkPfrL880vK1rReC0lW5PGKH2dpIILHghWluzUsFFFb10hhr2VipAiPA4S3Rue0htmD/kzg1
w54upfbRS+jBEnPxY+VtC+RbtyZ7/dzfd3oHb/RpvXb/pgN3Yfbgog8EX8RMQHCRysQZ9BiYGCdv
l+kO/9qJhSe9k+Z52XIdvEwpkaGemzquOmKRb0UDD0RyyKOsqcrm2nDkEsSrFxyu9sdrOpXMMXQ3
d1kMe9+6Z5wiNlbpsdDeinSAvAF61KTxPrytUT8vJxuKZKjK+i79ypd19TOWJOMUjunUELFdU674
M3DliF2ruxFxRa2JCUZuEiDZ2yAXnatt/zUXTVcx6iT0+ySGkg8seHf6/cEreK+X9hfZmhSYrsjU
RMUeDO9xii3dgIxrt9KPuJRXpG1orD23m/kU/8eCmdCqUTCckQlTYdsahCp5oFOgPN28/Y/adTU4
wcV8CZUo3+FH/rwIYHWTqlr8wEoAGA3C0h0MBZEHtc+QSL4gmJcoerY01wyki0FJkJBwnWBAB1b0
MhngK7rCJwkr7SU7vfBu1u3nshdVEpwkH1j3khqZqRF8+Ll7/CjcboRLthoGNksXJyu+iCwuTqra
qXSpHE/Yyg/Ux6tGetb4ufQoI6qHY/wd0t13RKpbf7HjDWh1cXSGZQdF9/UHBkPKao+SDXTuILjx
IuDPKj+bMfKPvQkCTaCtZbEyhAOwXroPgYV8mm2/UErbLZ1NUZM3RPSNvgyykvmrb57Hent3Xp/l
BBuuFE3/ou9Ypn6awg79uWzL1xF6qXKpY3C1ZnuycA4mOx39jO2CfiFdKiTxCePJmITFjNC7iym5
RvY9VhSOM+YXPFdJQSn48xfK9GSv8KsiVabQkJTesUET3pDzHVDMezL3nSpxfUT3Fu14voQ1Iqey
1Zz+cJ6Av24bj8We/RR4Q1iRIR9xwCWAg2dN+SW2xSZfI5pxH4agPxTzb17XCyHtZH/LHGssrhyY
464qAs+6uizQoDwVI7kGk1LtYDw6O8IQMjIZRAxHkpV3LJl5H40SEcQorm1OVvbfDzyHHY40emM7
5G1TNSfI9sDaqsfupkfgP59kK0jEKi2z3chLdQaSoiFff6JQi9wUcLp/RpHVV9A9gex640QyyVPH
iSLaa2jrnQIqdwe4MedojgbHLStu4z+ZsSDOZf45ySCuKKIz97ua+IDPmMrz8N2q+ko6q/QaOCwh
BFnwazAu889pMDa3F8VWeTmBNDJWKT1Rh+kTXhd20KtJeJm0Qq6lObJM/Ze6PM/6FGV0qSBGrpRr
XYcyoL+wEOpxbWstxwTP7mIDFbOSrK3xxL05LWi4A+fS99d87lijEnbXcRzUwQTO9X7+fToljoRR
fbS9omjgpsRvPz2aDXH/kXKQen+pD6I3fStvLDs1MsPoWFsxQ+uEjVb6zZzhBlC1b3bmAtU+rBKO
ViS9xBJB+rXEjzhX0jtGMrVud0AeytxE8ddWYG9SDic8Obng1nwrDREFeK3M4oWlgVJDfT9c/gNl
PRGRJ40cMiv7JTQ/vitOhlesQwrVqcGC5Z+bkh0VMBE/bHYyUa+Za1PHF+IMvDoKkdyMVfwJ7nJE
5D+PKQwEezIiNMMi3k1g0BwKmKPa2Cxz35HLqFg02P8D8irDUXv39Sk3Lye8ECOYFyMQkmSOxwc1
s1w70FaoFNBeArCeGnHnmspBQH2r7FnrTOVRbgmDbhDLhVGOqCCXTeIC2Q/FE2kF+Xbxbw69IbAp
Ir7pKuRi+uwGf7ymwHB2iJbmllhTVMSkNTi2q1DgcxtrKSU5tFjvu3e8AkwOq2Gy4lj1AsY2O6yk
1wPIs7XtFeu03mwc7CR9I1Ip7B2LLXUt+IFlIWF7TMb2zEejitW8+Nkya6UE9j77rqEHoCECS94W
ef3Vyx+aUX2qQDT0a0KIjvD6kbcaW1Tiv2xaKhvXcsIJFLydL6j959mvXcrU0Xm0huNlyefzndpi
SbGuQVsCV8qqcxP10nylK/xWo/BEKCc0s0Y7LC71hByI7UCCuF6as953M2Rle4HpeLiPm5nxjEjK
ET5qJt9J9KSMTRyNE3ue6NsgwtHxVmmhG/H1TMgLXTBBMEtbDkXwELwODTwYPD4NjvZbFXDsfrss
bWYpfRn22bxlYXBVePTPPOHVBSirZRc33sjYOOk2eZu3so/OEuyiCivVh/i4/BK0oVggv8LtMcxl
8/yTmpHLIG2Mkti5fF5hV1SCxLnGHtnKQqULr62V9zpkgOFCuBPf0FCO0HSbvCKD3YxPCwI56xUz
7gdsEyxiH1NuarKHavyXfJhO6Womu9t4pe2rUKEK759ctfPGCMfofhJgzNJKSP97sGh9F52BVBxj
xAyTH5kI0PsLi+m1ty7Hi1Tz0hO9UVjlIYA+0zRZIhsfyVehZiAxz0tRvdxHczmHoBAoEH6shntA
QUZju1k32BEffkLtqL/fZFQQ3jEs7HcnVJSt/JyqCWPuJaqKI9BIhiG6QDDiwkNPoQ/dKzqEbYk5
4W7AlCpQC5qTwXFsMLl9MWUxpfHA1ceeLJDdr7ft/3Wde4gxjGVqM5QEfRS7t7f7dspPCPT909W9
ChTIoxN7JywZTh/sQ5qb/md3ub29+kDBBOoj/cHouG2XSu2u7V57k4ESXS03FTlADDQcWROh365S
iBKe+2mpk4O406MzwY2Vc6+qoiUSWnpBcgk3iYIaUL4f2pdk+f9mDJkfUXuzwNKYIN0tZLSOeEh1
n8RM8FTtk1+XgCTXVqT80GVEgey2ZxHf70jOfSkGIdLvRGaIFx2f+bbRzU77pCa3yYpEUaJ2AXJI
Nte9WHWAA8DhgjNV0Cg94esbbeCu3rrzDlXo7rY7Rys2aKF+XCEHhfuCdbiPtPft/J0tPR/Snl6b
56iJ3qhNybOZ2qSTR4/ZWvgD75SJCYJgHRV3dRWpE8wE4SMztY3YoXIqm+lt9wBY8RIEF6wFxG1u
JvsNk5TFNdwPKGeqlrXHOsyyijfHcYNdm30A33L7B7K9RDRfrYrh4ZF+6W1Dpci3ddLFdWNwt/MZ
+yv2LZc1cJg6yoUWGnuNL4gjP+k9iO5+kY3fffRxa30jd+dagOn0DgBWW8R5dXeFRYI6jzrWZfRg
uKAiZyt2FrtdUBHqMoEis4RQ3oN97A0xaI/924ztb+Bjy17AuL3DtdGcPaLSZaeVfyVfSp5a1bg+
DwcGAsFdFlmmDpPI/DKRQFdd0N4cCMibwzdNbja+Au/ELB9p+K3/lnLIBKw0jlZ/OymqlxdFQeD0
RDUG9eMS3r/Xv2Nqk7sxta3NxlDCIwf64+MbYpGtJvSwynBjhMoOInAx7/5WiSDr0CMi0V84zoZ/
8hiwfWzZhVIJbTOav/PWfVIuSfb8U+xGIzTBpup8TPzFfbW9eAMHPFSsRSzpzjvWjtIgNy3UwX/R
wCP0nk6GpeJmdYwUN81VT6tVNod87+1squhkPhjM1+aiw5WPcG/8uL1ps13MsQmbKipaFBm/R4Kx
A2X0NuBCGQ/Yo+YzSIondrKwscG8fB+PINtbg5bi8j/1t9xGbPjdO4e2k5gwfnlgux7uwUbA6ev1
HZpRal1w8irkT3lEg0x+6CYNyM3IasSPioeNFJdqWDHck6XuLNC5x33gpaNSnNjGSJZd2fn4jE90
Js4Bgw0hUumx7sDSoh3oAmw+sP+YhUmFg4x3CH1GEflRf7OrsNuTXISXFLgUB8FKE9Ijt+iVEAOz
secfSAtzZ8Who+HWEmRFsJNgwBK7MxkSO+oWamRUmwJ+M5NAYsQyyRLCrzWNC14DEdlyk3/FT8od
/MdIoaAPz+2SpsjqZLxtO3HoHTW0W/pWHXxs40Q8sHs7FrhByT5V3oIHCdxyF70QyvOTdiWiHgpI
D9cHLDvRTYNDSzDa0awC1hfabKMRJuA37SmFPrDlwcc+ktZ4LvSsi0Sk1ABpmCvXCh2iPktS/U/I
yarEH031ZfoPi8SgHf6/nx6+s+3dsC0YbXTwD7fPAFpQGLkpaqvspaoHR25VKsW5MvKMu3NB1yU5
shUt5LYmEV4tysPQOw+a0M6q48mOuI0XQDY1WdWSPUMOf7/FhqFI5oKWWEKlDhaXybcIqE/2jYBC
d/1/ht7h7DBTOMhLOfPjCiQFygsCfvztw01lvsx6sQmLpT7mZl75GH2IBtDFVDBHiBFOkOuMMFPv
I5MoCDyFO95fNodc3sEmzOHgt4seiaHpfWZ8IcEE4qoHqXhWNESkgMQdnXU4Ou86RlHLUC1M3N7b
SsyZhvGKL54GRC6zORx+l7WRFXfHCxKUAHx6BHViqcFhHaRqr+7TdlTbCnOwbrmmnhVutdbJnAxw
D6i0w37qUN0YD2Dm14fAU/yJ78yD/SMzfiae1WOtnfabdZZ6MTB22nlV5lGxJ5vOmnLu4cPVJEBS
JhuDJJBL4lj4YBHAZjzM3QiqKIRiK9vx32q7/hvhznwQJgAMCj02wWUugS8CJnycwVXlQJXR2w7w
yS2qijvXBVADp+J43soYfV2j+PkxLNsPmp011F0CJoG6OP/hfUKHH4ac8bZRJ34+5z1XiVms/hhn
LKxRRiLUsSxqZi6WfCnjMprhibe4jHaY8Cjvbg4pBQpS3qll/U9Of2QNcqfU732aAcJyg3eTMv57
Lk9KN6MGX0ihSzqUUDjmD5ANsjlIJNqNVt3BsJ+m0YUI/WssHpBZqyAJcDdlK9369WWXV9wdGVJu
rCg/scJlgxOcfti96vraA9cGRo7MFzsXuz8VK581KMFka82x/IW8k80Xq7/j3rZOjdXsBjHzdjgE
rc/7GJhyzaGiy8KPbS7R9QGo6n8z2a9KkSkSxZyOoFaB1CVHb7jTH77r0coneB1po4idXZ/S+wJb
rFGFVKrCOVGWJ3m2lqV1eowJf50lje5GRLq+Gqx+0/MMGIrkS4pQOBqOxz9e2WzEYST38PcLAT+J
taOSmudfDPDh3lb99Eyk8kXyWVq/K2bYVFc7zql+hpPMogUfER6ULrlvuaOZZhQEgd6DniwpgQHS
SI0LUkdjra/smetoybhQl2KW/gfaHd79MzugWUWrVWPJMOyrJdHDHM5xQdpdiRDQkBEAkynpK68/
zjVwMRtXuAztZ0MMx5DYt3gXGdkm/utzGb2AhltrOGN/82gvCcD/co120suoQepMJpy4fa5PlXQe
OYO392+OaE6+8DJaxFaioA8GTuyKgCNG4fhHOHL9Q8bgW79XHlLKz6Nd3rmjeC9YLcdMAp/w07g4
y3vaPE/uUK3KsY5f0Ye6NWJbwpCQ98rY9/PsynXdUriNASKVCwb7AhACahumOaEcX/ZzfVtrwZTm
ntBUb7RR3frG/P+khoBffABgOO+A5loazonfDBnBe7s5XlKUMgEGzEYEZ8HlKxGzeP0yFGRDihF1
UKR82GuSSzmUjLWimVc90WF/XFLdoeM0NTTSguUK9uDZPwDmzzyFAHTm0Y7ih4dSXcVv1N09GdNG
L/M1jxEKAb6tjieYjy6cMQGzwCZsvQ5iHZxPf2Q3N/8Fa+K5oLf3ZjWZkFroB5WfoGFJH9jYuzf6
3BHkJtKfcVC0ru/eYSxXDgv5Xer8S93eqPm7zXOn0FoCWnPn5wYPX/DKAT3WL6Tl4wdZU7hWjvdr
YLYnC9XvTeVOSwkldvCpB96fnkO5/Iuud510lBT7a3l9sqbrUGSSOnmNO//aUKi4jsrym/VLrAOS
0czR43PE1J82sUEsIvUWU06nn0cArnySx4LU/i2EV9YAp/UPBRhUiU5++hON4E0DxaV3QQijvx1S
GrF4H4l47p3V7/4bmjg/kcWMDIPbOUMl6Uz9n/9TAur0qBVRRz1RusyrM6mMvuyfcF8RWZn1Rst0
KCXZYH9rgJ5lTgunzQ+9UYNOhRGLvxKy1iUEHmlTN2cFMkOGe5JiuAh4EeuQyFV78UBHJTn1JVWI
+mNRSOletPHiL2R6LSYNPtYQ0bOQSJZ6woeZAtgyP/XH/IEJ4rasH/9JPhYeTiWiQXInKlh7Z4kD
gE96keSnSsbkIf64AncY4z9GdzdS7saPJZ8azqRw7uMdE2MPnCiCpZJEI1RSzHZZkCqSfqGR/1YC
A+tUhhVC/NfR3AYnDNhxj7Yqw1kPpAobtRZXSVD6wEC+e0Cxtd71FNaBFLoAmgUC+t+B9WgDvJpr
QMeNH9LGpxTG8lt8A2gNDa1dU1THVSEy5qBo23fuhZkDhmdAkfHQUDTfix75ODyEXiut0ifGdaG5
5w0N7tqRoafSdMrA+ZD+xtqm6NZf3FyV07r3TEoJp3VddjzwRnZDb1gsH5I33Zbw920sy7N0PjKV
d6SQcac+sA3eM54rGezDKsF8fbaqqd73ZD1yytqSpC5ZJtLJW17uOsHlD2/B8WJd6DgC9nIu2ntc
IgLEjRzNb0djjcolk9F5ECr7rgetCYsjoukgSle+uPX/KlTcCuOo3HL2Kgx1jMPtNTL6lJoZk4pS
+VAr0Y8bawJyoV9t3QR2yRKAcfYPs/t1Xp3Z/Q6ht05IySSvPlmMc3nPEnS+cGd+Zk2eztSuR77G
X66wajYmGd7AN5uQyRSndRC5gnDtopQWORZIFxgtNwzE8G+VnyWcVsiw417oSvgaoVmzSwH2kQxc
ty/XjRqGdBM8bdTC0CFGRyTuKnirbtAfsrQ8xVzbKhoOaeQmsekEJzD7ui3CxnEAjoLU9oQJNKtf
9ioJo8YT7CU7QaUpp4W+fcLd5wxrZ9r7YLjP2z1LdSKqzoLgFjSyRnlB9cd0cD3FWggC60BJF7oA
8YnD8z8mPjns4bCT6MrVAWm8h13ZHGlks2lSB0lV3Y4joR4c9hWi0AHluU/sPoDAB6MVdM6ldCBv
ZeXibNgn4uLzFTQRXL46RBgmdTfW7lcTGEyzmGdJit7EPoneR6tRk5OogV2HmXA20Og6z6cUQr3o
W5JlJV66Hobn5vIk0mpV45902zoZrF50eFe2bkq8xG4qclGrIo0GbiOvM5oQUVPMAxiATU7oEdf/
neqJeZ8x3Lxzog0oFGgdQLuU2v9b52e2YwZneoYNmenMZvB9tlhsmuychrnXXjVvR4YKrAYy5MwT
9Va5eiIrLSebA6HtKn4+QD3Zuj2L1PcR5XG0oyi3KPIj4DgGU6OVDtIG5+lpYK6wOgFls4/PhtR9
YwHg0n84uIZllEuFJ9OIY1ooTUhy40VMCia/Sz+cpTbvHKhOcncBrpBFQTSVRW+huRt+DHdUBak6
m5DDr1SE2hi3iB2yZq+qmzDTtB2CG7eFutet1X313tWddKLPhSe0HCD8pbhRpaY13fci8dMUvzvP
Z0W2LmZufh6wZPtedYvKNR+0GrpzcaX1m0a/bAQC/+t0zfUnyhbqDfG3SIki5GvdqI4rMDiKFma6
yVcy3xBwafMhYXsQprcXActZ37EFeBtDQut8dl58mjyhRq+ht4NawrYV0rLtQWGFhdlzTjvrHyiK
V2XR2O/TEMJhw7x+afqh2gUdxpbaJyvCiqHnZSuh9YZoZR+FJhLJquDCyY+AdsrQd+E+if1yDq1d
OgzrdM6xzkREP0ItqsbFp7/Gjb1YPAWTqt1NO3NYkowDfkV/5oxcuXJXGMyI4oY/Z1XqjJ3oTaWy
eeQotLrlBm7csZfblzYs4m+jp/GAYxw8bzUpUauagPSFgtXRJGVlY1EKqXOfEOBCXDkB2pOKIkqO
VmH1j0DgtXp6EPkKY+sI+SB99mFGDFCtS0LXLkT57SznmbbDvqnGog4A1KVuhoiCtZ35QSX+yXGg
3T2Zlfr21ZZ2tSmomEMpU+Z0gxnDFn9Gt1P69Qn/eo7iTvXPpE8G0GjEuC27SQqvTPze3eH+GHqv
hGo8MbxmUgqDWcT5GYWEWwiaCWaBn7ZL5+pHZPzeeuOlSDuXgT4uoVZfMePr4RgU9K1uwbByGuei
eyFpZx3ch+ToknycuO2bLXED9vVbrWCJVG0XOtYonwkClfrzybKqJZWiGfcMR2Sw7ySzS6yjOT9u
RRyQoG68e3RsLY+SQpb8noLURSSplyC34GZmuSfc1Hfcmxu/gAjiaeJHSAzFeLxqLNcNH2nIuaC3
Pje1kKOia8UZkkGP9Y67YaKQVGCEfU845HohdAsWo/W8yyh4vTK9RedRrjLRWUSWY1WzscG6P2zi
p0YJI0/rs+PhPm9nYPN2IcSHtTdbdTBYli6uZLxK+epfjptqv+V6eHR6ScUlR1ujd5ttuCuNkHnw
pZMsbWwputl3/Wm5IiNddiWGW2Av98ZHCGG9Be1EwngvHmyk5Enkgv20PY+B+aBCSlLkm4Qj0iqQ
1S0PuJfnoPBFvOKJx8nfYcXbcbUVB/88oEOceooveR9A6/yhI53vi0sjb635oDpwA1URt3rmqIze
UWmTf9q9lPD7Mz/PZ5PdNz7xoCHNiQjRrDfpE5tfidGCg6Vpi1keBClUPro+y9Nd5gfZDXogNy87
OYhUp+Xj0WCeK6Gu+srA9yedmSXprQCi5yIa+67ZVxWUYxU3xjUaIv9vUWhW2Za/c7gucIY5zB68
r9eE63XejhvN/0ZMtbhIKJCeUmn9cgZn1r1XXsl2RD3ZNWExkai834PNn5X4J9u9KvSTIewqjBXB
j87nHN6GpKQmltmfLad+Va3QgaW8XZd69TAwffMOyyrcmNEmPuo71lD9tuBENwdZlY+yem+x2V3L
XlbdC1ScMUSA7AH7blzKbFEllY7GQXnReW2L0my8biNLZ7/C6GwVRH424F6cd9JHWZfrFoKZohgz
kP0x0jP8TFhztPWuWHtK74miXbs5/CEv1usZnhV7qPTT56hWiO58tWBOlecFYj5jD21RY9omdaUo
dHs212mEIondCS8WnrD18RAZlOwCxHJWuSlblPKpevkv9FK73wAVUjD/8kTwco+lff+MJtPvxsEt
x0nSewjuUHtuoA2h9yKEKRGrK94FjwgpXfIMO1TIwfhYIVAh0N88WAgfKvbiD73ERswRGkpL9Z9x
qOU0+3PvNp5H9E9Rez+KPjOyCv/2VzUTf6UlO+k07c+PDknNEad66s24vyayQ5HqIBABk8oRl16t
8j4yGOxvy3fye17pfq+Lz1ozol4/Eo7dYRwHPAKHRpfI5aUEI85aRCYGJ5v1dYiGiLJUyICr0330
sSubGBagW8he88FcMLOkMzYAtFto1NErI7KZ+NwBKZr0wC1ruInzX6qmHFsYnkvrDvNR13Vvhgxo
Qd3w3Ec/i//c6ISF4+g/lqmCu0plNSSjgsiTk+EHRGyG4sSy0VV4nvYwo9AD+0JkDnTeqwzXiuJC
zYVQkjFX30qxOMaI9BjEjg/N7o6mCxfs60GQlY0j9ZdQQ7wb0DrjP/TvzB8GXQkETxZbzrixggdz
M4xqRxLTjQkRNgTCYtAI12A3QKd+Wa3kreHC8wMNXneQJRFB0w5mHOGezgrJtSxGtEgcfFEu88R1
LP2P4BW27wzcvjpRPzHXCVxoUyxLp3NM0+2I7OG3JHg2pjulYMaz/k6e46kAw9A3SNJwn3X7kraH
9TfObbvKZ80qeZNFEUjbpM7WMQd/oDryh2WBiBPkeHUupDNaZbfGd1d1t7pMi4V0e3ZA9XumGYTM
5kg+OAn0MmwAXK7oSpB5IME8AhKLAqEDRHZyxWalrvJ3MabcUXj+5cOTu/LyoKXfdJdQAFbV0A9E
+0IYpSXYPliz9rlfeVBonTdC0a4p1r1hXW2AIWu+fvH8TvtKvP8GixpuJiCh2DxmIGUdCdlFg0Ha
4p5fjwO3IHrwnEXV7emDUXojQ0LmhbNG9XSsnhRzSodmIrUAgav9f0611KfVQ+coBHBQhrBHS6Im
dJe2eTqIxoMvjsuqTisgdKnN6UM3A4wqEg9PN1wXHjJit9jF68Sj1zURAsRLgCwH4jovEGSH8vCi
EEkHWzGfAfIEVQQqbA4MBmHjAlbi3ARl/WMzlC1cBX3dtP2xqOqA4jBhSRIv1c2WZx2yQvT6uCnh
3yoZ7XIeAjQgku7/x20MEOpVq1BndU2yDknN9AYJyWd9+T5YoSP1e/IeoxoM7oo6QVBoTd6aKOBq
PFNvHMatmICs6Ab4bSBmvT7zW+01qV2g+y3r6uMxBak+9JSiW62swuSpJ7TEWfbtiPV6vdSlNchx
uA4e2aqffQczBaQziBrgrJ5pWBH9xe5lwZ2nwjDdyKCw0rzKKUPbrga2FU14+y8stY7ht8E+eEWl
cZRNmuzP29tid9rYor6As/v4cbdTMezR2idYKzYDl/cCtvB3o0xaa7IAH9AlLBLPKUULBNAw+CE3
BkXu2OXx0/Z+ASeaK1un3nPnD3+ds3F+eEZ6Os7hbhkiSNCy9JsuQz5SUi5O3kiCRRzNR4ps5Zl/
H/iqf+IztKZ8q3J+qClvhOYpAUG73L5KkO1eJefln9KhKOBuftbfeurihqxV+xceAzYV2tsTc5lX
NRAx51G2+YkD4hFxit5zOhgwRg3VGy/EEdCHFUPI3CmedL+nA0oJuOrLyfdG34Su4/z514GgxN+E
Y+cU+T+xCD3yV9bzOqnnQyY2xZvkIQm1jIMzDaAqRy/epaJtRkg7SnJd0tFsfi7Tt7okPKmZcqMU
E2cbDOv8QuPRBS04jIRTFYE2e+/18NN9Ks8FFec/hM9Yq65pVQEuFaKCOrlKojlGHYfgQDc88sLs
zsJ4eI/P3ggo/Txkm/LWtv3mTEO19t1KEXbiBEP2I08tltdp4mFTPtq5+08Ly2l0qhbUaWmofBH8
YshKLdbIIUvOt0O+ZfTTqJt5sYTI7zNqjTwsNmZlAwEjDYfJ4Bed88eclgtCx9+pGIVcL1ahM3hX
GnKfbK9amliynhjHty+6fhxizy4sIVw+5VJen1Lay8/55G5jkZPc+B2GVzidgsxOsE4AOyl+8EXZ
SG4TxcbWgKcCwjBZX9MgBZU5gdNCYXSZ5iV/d42SHJpTjvDPOMgMRx2sB+nkL05+PCMGYm88JnKW
kZTRV7h54xAIGZOHVeYmW5yLJY0pCU7+KG+S/6uu1mwAEinwB7VZ6Pb9Ho4vC+6waMoiZHC/fbLp
lQPAqQPMEq+8s6xHhBmURPgNoOJIdLT4Hh0BUDosCXS6mS2KThlt3Brv959CS9Sec7m3BhXAQiR0
LsLnHWlnSnxOezFtESghtekDNYTNOHB8VJMbiWAzP/lD2m7T/XeafjTZ5zjDH0QoQPShV4+hJuue
bpFOWwxVC+dGBf8DRHcykUcHCtEJms4qpTF4ElDWKkMDGPlw9DbZp4a3A55pKDzt07iS4ZPaOHx9
Gq21Armtrr9mVz/l0i9ZPfyPoh6iBUFPaxXxAarCZGcvOxb9KFobHWorsJvpHL3KMJSSLdZ/vvq3
noGg2nX1w3zMtfzixUfT34m+B6uvJbinrAMhBSGYe7UpWm0xzT9zY/RZZvWUBy476WNYRC+IfUfB
rgBWKfTk/htAMubAWKR2Gs2CWR6uRdZFFd0uUdztTW9CYe6PRlVAdB5+q1Zevk1qcwXjOEQm+Sum
s6ul6WkQJzVl+tn428FiAOeeZlzpbSQn4vncHtyIr8O9uVATfTBU16G4X8dFN8rYchge1UZ+ANAY
DfWLDgKq+hBcXtq1NiQ3Q0zO1iCBhM/mef2kHk+3qPYoUStmx6o0hL3C5HEcC76mGtudf1YuVzHC
6MXn3Dbu0hRCNAho6DTHtL32s7v6AHMs/NNj3adSVREtGMViUI8znlElPQKHfyxU7qKQ0j84s/2b
6Fqipb7Hrs6Js4BfuqCFDIxCmknSgOcrHcsjCGGIAT4HCk2WIWthFLrwu+PlOswVM3hQZeSG4mXb
YPJ8Rlf2wmxh8YBh/39hVNe9RRJS2njcoEwc09ONsMXMIY0SKAqWmRGW3R85rZ2Zi3X+2CxKNkdJ
iFTxPw71fHXsx8/PUxsBWLEN+KW6xsktaHSmZyqaMKAsQF2ihSdCBcqlQ1WIDzSZkSFpLgSMwajq
tUgqqHzoJOvSkinMdNsgAdA8TkIYG8QkegYS6RGlmwG9cwnTe9nCd3T8IIaSJsmr7lGwQkKLsuOF
ToRs2r9O9NA/ZKjh1+NUlGn+DQhIHWBRvU5O57UhpHjjPNIcwNFD4GdJxL25/ot01U9nD9lY+lUY
WXzz0ML1r13PDV0r32k+7HbIuAjJVpTDZU/AXxzBvEN21xomZDBwVWUIDUxzugXYDVDURkVl7Afq
szVOnq72O4NVtwmCZnFrf4+H8cAF0HK36cpB4yvLsi/SL8huVg2AECHInTms0wfd+DTZRr6kQpq2
ZuXDP7Y55rTONlTJ2tHFYNfbmR7qo92oUDOsyuNDIfWnMWeRimpLI3k2r3eX/11c2QnQSra6kRud
uojd+YwU4AU0ZB6VmLFCAa/S9pM8R6dJ715U02iRnkbnYGqFCNcko6WKfEHte24t17TGHLca0+jY
s4u44ICp1BuDfGW4l69KlhP0BVAyyfGbeDmb0LJ2PoKI5ZK7BOD4qYnOpxVVSg7g0xaYXBcGFVY+
gRDPYnNs5YMqnTAtZOJw/ZRIjcsiPAzIteowS+irQKxMvHyltlG3N+n8XEN7bip6KW3YvOPcWnIg
mx4+mg/QbOL1GqqPiBY3KqBDwWdnxaXw6BtRphKXosFC6k9Y/lR7emBJJbshR+D2v7GB65ZeI1TO
QtoivKxtaAQIgEKil2jelak8PvNFnX6vFGeqIXRsoGlykxypuaLeRru1RWugtZw+3uggM4BbfdVS
pXreWR053NbAYkmo2nSuDTesbJbRgUSu8wTjIidSkA6SixX5toS9GQdV4A6mb9NhI8cnhdKlE12c
zFmexzqayfNGCUyyzu99+md0i0IF9qKV8JfOwIOcvhwlMEPioVwqhm39GOlUU6/bhm0cO9XmPPJc
909zlT4Oxd9q+/EQIbkHo4wVFEXfavCX03gZtCq2qk/TYsD6T7X+kQ7XsNzcG8TqqdsLgK01Ck8A
lHyTCVNlCgDQeaPzqrsFtaOMXnrRPHUV/9Wo6d0MyatiM2xFPVKh4EHb+dqs07gNevq33m5jO3p0
yEk6LLraoE+SWixZPgPP3zQkSD3+XUDA3A0AqvnGWjKtLOPsgIHBfGq9KjmAhml+BWAOeemfhAu2
8zBLS5R5jrf0B2dQPPUqqmISOtlF88DntJvT7zkZYgcAdiMIGIhqNBVDIzgpcBApO3s/W5sTiJq0
GnW98biPcaP4sGZPLPF4EfcKxAaSzOabxCMd00dRYMdNd16vAG7C3mS/cTcJniq/WB0H+wnF5GnL
0wweBJYdyWNu6F7vFx6caAzpNGyZ/zkPa46oMe3htqHoXqwfl570e6cDOVeN0fenBf9pkK35rls2
o47fKXwINYFI3q/b65IF7u4I1GBEibotRjuaj1JbSrtQigX5ShMVI7OQuv0rjgpTZmbF+EsG8J1Y
6Ne4ZnFskcfUCC9QqLOdJDO+Uw8M7QDombRxEK0B22TwTqym8w3O6WnWExOLYoKFT1R3i06a5NDF
GfvTwQhvR5WqwhpwIWr5uHPi0ckW5PJiG6G8iAIhN1J9P282FOd6JlIZfoqtM6k8oGRNlRc7dPSD
WfblrNBqwU9S33YivI//Lj98L5n5mPWScLxbsTx98l4QLE3T9hiAo+ZrEAp946rVOQiVLFKpUt5p
pHE3egnTpugAKSlodTQ+ugYDEBATeUcvhpOeACFSq1uIXRFRa/v2fnnxkgldU/pU8BybHx+qySaJ
EGfD9uuVkBbtBfBH1X772wwd47OHgDEQY8nWAACPRzAQKvZM3vVBsgEX1rDQnX/AT0hxBAPDeU0o
27EGCf1UcN4Rs98WbEYAokSIzftrTrvttzDTRsD1ruSwnVZXjkRluBXJyfbtZWI+5bqEOR4SY+Wg
TcBU/2UHYxHT3c/inCNZLsfR8rheL9fYgiSErsem0XV9PUP6sDg+lm5pgOMH4nwj6YARPJAQmsEF
Ic4pNw4sv+ofyBByyh6rJxCxGxGx4Nh2evwGQiyZIz0r/cgSBFjrnO8DGE6Clgusme+feeqGIlNN
L4vE9lOUXfI3U7YIBxhD3WRfTRT0OgvYZ6A/R50BNtNiKY+LJdLx3PvI4OgLkG2xp9+zo/9AeMjF
PgnE9v1Lmp6jVD6o8dgqDSZd16igzM3urt3ybjvDvfAx6Eaucd9XN5ABc5swAByD/fvXBV2HIj4O
gO8MPGTB++2xHlade8JHD8z+cja8nJv7YYZhstehyp3Syqx312nfxbZ24gejbi95GaG+6P2GIMnt
yjn0Hn9Fb3xvZF8lh+jQ3Mm+/1TtcZsywXe0xYW+ndanqUcjSebGxNOneCuA3YNBmgnLJaRjciZB
ak20JeFvFmmwhEU8MfCukeMSTFWN6gPEnN48DgGPmT6y2pf3Xl8bhEROtbPrt/FiAk5AQHUEajfZ
ObzmBMhuVexann1yCAAlCGk58vua25s5RNDHHa+cWPPk1LryLPLpcZ6uADSAMhNRLIBwvfjJe0SK
R7zFFIfLFCflpXtcmMVI00/EVHariB0SS97ksgTylyuWN01xlSfZA7x+QMKZM68DG7rGudnwq9q/
ZB0jIs30orZBiOMZmLS12KXPGIM/Fw8J21hNcXfzTwWn+PYHSd1PeGG0OCUMTTC32N1ca9ZoeQwq
hSdJQHYm0Rp710zoyJkplnMYjAxpuxrmoQcr4Y9431un6JTWmCkwhGNWxD0bwf3T2pf73WJmXLTo
ajrb1rGGw7qewaUNplyQk2o97Q4nGlkFro16uYU3Wlh2nunpT0w8qX2zEzcOp/Fk/0DerW7Q2F2a
bq05NPkos+wWOC3aIfnl6E3FiVBanicOgHoCKIgGRKzvFy7XBFRoOT3sPbl7oZdZUvKsXvX4cmZG
Z2Iitnp1st/+Hi5aZGuXmMQwOebBjNjEPBMwXOfMsjlQBDEppadeeXmxQvB0YuEx4p9iqXoGLaJa
bsdlmA3HBj35x/2ej9JYMYoJ4/L4AtPVNYnZ/3gtvF8JGdQC9xzJ0OiufrzttSP/RK5+M3H2H/5J
Znq4XXVvDd4/eOPaRoSL3l3FPF5vM7naAk+Ngy7WbX/SKEXWi2QNAozCEXecGhkT5zTWQpdmDGFn
PnvaHTDDkw3PBjagDJkhyo0A6dNuVU2bb16VBt+YTGptiTNBSgBRuB0y9Ozg0SQRjv/2MXA+NZj7
GmM03YYx9aCmADfyHfmfLVD4yHtpab+1Dc6mnlh2nXwSSQoXw/lVupmz6AMEC9QyCGeva7bXgnOv
OXiVx3Fr1mpmkMtUpo8IjEuoJPy08BTt4LVvHxUnsVJlTI9V6W4DF2gzrWWBbTy480aN7SuNo/AP
PBgU1VHkqPxgBaItFUR6OIZH//pK9w8TbnzCu4/43j47nyQT+fdFOKdUcTStUjK21y02FZaaqFB7
CSRS7+DCCj8n5XWawjVO90lUPv3jmKB2+rEjQR9TmXV+m6LuopY/gdzL5YvnFIuJ2iQiN+XC/fN1
nLOa+doBz0jwyJ9FVjWYnSl3HEgK0060pLJ661djNf4AhPR208FRkZ+KNauH6+6ZPg3KkRHaNnj3
opEDVkvI5K+2mpq0/H1RT8ZMHBOs+RiMSuDDg8jT7E7YPWnA0a7Q+pLTZTBj8yuOMfgMCn4HQbiy
amfkr5nYFrKPs9y7izjuYG1pGTJgkrZEBAWvRBmpncgza8SZugqlsSoDqbDBoz/l8wQ3Xi+Y0elR
jYaSJRDeLd9tXLUMLITidePT5tj/eD+Bv+U+PPDY3z1Pf+lemTQEIv+5bkb8JCkto/6hU3d4J/5P
adotz2bqSKl5QpAQpSpKB5gNvEG2e/gcW8ueZ/k4R1uv2/jlwY0UhseuUJ+z9mMW8nOftJUsK4CH
FXJcKYbrdl7Tq75UVsFbi4J8bkypKm8FOxlPBusNGlkrds5cOPEfWJ6ulHIfzYO441ivIkx9JbUw
UhNfKYzHSPEinfdqQ1wZ8MwLyDG6cYWt5cN08n21nTRq1yCJrTBfvf1rqXpf2CpxBMoOjIviIb1Q
wb5DFa9+pXeAG0i/ahhSxiLswrZjcMfike0H3TY9C1zYaRso07aRxe3T0s4Ip56Jq1JtH0MxVuGG
YUHVJBF6hU4a5CPvu3Ci4iw2tOxGO7qpGNpA9t7b5yBWanBIAuJTYaUVd2Hf+AO3IQLFgp+ZxceJ
nULOWCpCD6k84gmSwVfMZnbKFQBK5zT7LTM2XnozK2EtwUH/e3ar9bUDuaZl4XG+/TZEt91Zb4Ox
FQui6g19uw1IH0KvorrFQcYrV+eMqiH+8G75a300kc1yTkU1mRDKGPlKy4+EG8A8KxTgUbuqpg34
UcOodaFpOhiz4wAxZj86M3HJ2C9xHmareKNCS4MpAFBS62WqItqe2GRVsgqCQmRaqQNr2zfhQS4j
JzXz3yKdaw2rkBXMZQDp825qUkLsp2oiZy5UwXvkw+aJrB1+uhBxLyx3GVB+YRi5USfIFRm4ZFTX
ppFQlI0LqwiGeRQz1zbok0hTqDK2jCDE2BR0hwwPh57t+o9HU2SB9g2EdhNrMZne9OeMWiP6Zd9Y
xV12FTcMPwh+RoKIbVa5JJI2LpOXadVNB4mcfm8AAZ1eZlo/8qFAnHPyHtj58xw+MzX9S55Qnlly
LxPgKRHfITDEuRY1Dyh/l4EcVx+S6VLZXNbdcZS9M7llEZxDmnKQO2aXOS5tXTbq5Ixek5cW78ne
ctc7+7+y1CRm5wyKmDC9eOjpemlPmWI0O97GRvCapidFDq2wFl1wVQD5AnBtJqGHm98tVAjhmBYc
H6UUSzdhuZ6or/HV9gSkKVrT6MzT+zRK7FPrGZFqL1pzIah0CgT/WzWNWFc+QxBG61zO+mkYVC2Q
rbq5Jw4Mwu9dlif2DNQbDT9lSBn7PK9YJBvitSE+tBVvKFfJLKtrpcyEyZhTNLQ1zoHZJf9/dXwL
c5nP4FP5u5YYRBS/bXlCuKFSItgVOehX0RTeh6VNlJL1SKwBzXGUYPuGCMC/7hmQViMbUAtWRbfH
dlx8xl3jaMfvGD/aqwdumW+c6r+nssyQWU4YoJYdGXzoyRZD7fr17/E8/aN/0Yz653HnG2klca7p
cZ9rBV08ovreahdRzDuFzCL0swYNsHltPmI+7u1i8IYYLsWdSVQuQIN2UK4GMLSqT8hahSuABg2k
U3FWRQ6con/Hhh4YnIpH6IAKlb3kSWFiAlVOtRzHHWNs5fZDjd5ibMVoIS5YWPoA1lhCeo2AFgxq
lwRmyRPLQdtXju0WO9MNDV+5k5SVUVMaWm5RGm+vjWPdHqZNHPiCCbwjqnNTrytqI98OG62/mAuM
HKGCrLCVHduPUiPVt5PQTkzFyHsWPPIDKi3PJ/+mkilNJlwtD1V7mswNBfIO4JVua0S79FhLKF1L
J4qs22ex6nWxHmmjXuSC6LLKddTXdpBkp8AtCdP989L73GGFPA0/7icUDuOFXIgsSmtAf5eaJyeO
if0PwCkDmjixcKKm201e/S11odmwvl2BTTVE7a0T5ivx16ybWOGipEq2mVcWoOtT0LyL5apRGFlI
L+qS7Jh/ddKRud7Q2PMWa/G7Matd6FFQNmfYhlMB/1PfM+Fjkqtt+CHqQzGOkkx5co+ULa9gdQba
hALSy6j9EMiwhHh+jju/85CqYJcFz88UHpWcuEh6tyQuJQaclcMcU6GYHJba9Ej7YD5NiFbMIpPA
P9vpYLhu1v9tFwhD9q3/+XiZrJHzt1CUcp07ltLqL6trp+dn/qSovpDkd/yA7mmTpYPbPxVRpotT
qVpiviX/mkEdaiTSUY9UmrgDFHx1GEDVemlsuJkkCX+P/QRxaF/QCWmJ31Heir6l2Jd+iidn7gif
lISDrhq1EXot1skLWkPw7krmBdJjmZM9SbPslUwUkw/IqVjc7mmIfhypKN2tUQCEV01enPRgcaNu
oxid2mJNFTfmJVvyfBT+I45xKn7P6CS9ctOxmr6PZf9Wd7KR/PxlUVUYiRuqhH0w6akPEhIZLw0J
tKHrZamD5QAtyfNjfjhKQ+W+FWwps1AVurfTCe/syEULn8EYDOC+ebICCFqEYxide8nWmjvnysEU
AllNG1//V6dlF4vvOO/Z9aq87Yv2rUchmqw6u1vpJfb67PbT6ZQLWh8QW6IGUGxYFKyEmZE65FHN
Vwd7xDDOVkA9Bv/JqEW+dE2J4ngJ/o43Uappt/mggUhhehk3wKCqBY1LZlnyTEPpyP+exE+StBUW
7tDQg+CNz4kRY/OlEYNyjyPhmpf2VzZwg05ie59GuJcBrebQDF38b6pQnYHhfCYKLBGCSR9vyU5R
27E4ANPjtCx19tSg/wgZcnH/L/+fCYNIagIN+Eed3oxRcrMRDmrUEuGxOBHQ1ZDVD3BNUp6gwFWx
kK/0mgM18G4Qn4Hzy3uSTHluYJ1AQc5VujRWQ1yr42wWSf2xtdH8qmAlww4A7mEWAM8Fwuu4AbYP
JSxrEoUaphVjiCl68HZe0mxRWCCXVcpcySxqDb5i7YyMy2gJqF40HVsmd4Y/voAwOG4JSPk7PfD0
F3t0FElop4PlArB6Prs7sJ9c6l1BT2L7ZgN1v4qEpvjohMkUqQdQ426JG3n5QbWBAAkf5T/mpCcL
w3xGzEwoG6VXcWKTMNq2gyFfu8PVU8VMckl9tJhmyQhYHc5fjpX8E/bj4VYpXVyrkQQ/Ql8Gum3f
naS8/WzCr8ZcT4kpQjPT48oY88n7IhUP85QQmWo3GGqyL8Otc4sbvx/qSwJQVFLx81qY1+eTlgWh
/Pz8erhp4VYRPtKwyKe/cXaqMX5yy3ifzYh/o8VDDOlBoJzaLIQRg0keAuzdrRgBj0++3B6ShHSd
qRqav+kAr6CYx4/T6ziAiNNISWdS+x6AYO9LVL0YAlTJ8sRLojS+I4NDuVQeJH0oCkOhFU4hy7WV
a9EuHUKQec3w6v7VIILOr6z9ZcxLDXll9Wbh+rhooxmyZuBrl+Xrz/GsQU+p8yIBylR2wCZbyEmi
QqmuZBTA7plkZoQGfZ7jrvZ2zjniDpI0KcXbpw2ZbqQ0rMnQJ3o9DDa9/B5qTdHODKAnz9JjuNjo
pADf70jIJUoUrJFOQUDWDSoilzIe3o8VsuVTSBLy0Aeku0RGm/o04gBmFiaoyRNTUrjnrozfXrJK
9K+WxuuFU9aSb05rFZWAJbtv3X/bNO3nIAxNEa9o1zuW/IGn6WlpdR+5PN/tckJnkSOdLyGoK6F8
Nw7x/acBXTXe04WjhBkzloaYpynr0vr8arDz1shK87/oZPzH5AedJGfE25itz83vTN1bdUPHvfaP
Y6JRghm64hB3cghVvb8jOToF3inwlx9ZSzrj3+4UpH+JWbKkSnvP/nHP8Qh9rAZBQ0/FpfXQ2du3
joqDjof7+9d5Std/wyOmKnsjVBJcgmtQxFRnoK3/cCI7kfsFAvRWhotC7MPxQQpVGoojIcWbRBpz
rErFlzYM2vksSAov6Oa2o4CSqSe1HqSzvRhsM+9cIbkkOkN7pUxAqxcXdJRzPoez1/Et41FSW372
CCxMFYR8yRKT/7RcbZxIeUpF+hADOeBRabJsOjSjPy+9JpIlGV3iJaVkwTv2gMscufaE19GvpTSH
8Ya4353waetZNHNyDGoQWN2VbWfhGTXMFbQDlgprKcuDglgLlvpFcexhHGu/orzB9C28QU2gc4on
4QrD6lWG+C6I+CDQOvfUTLcLEzcgnLXlnwA+HhMUVM557h5+FCy8hIFrzGv/215+kw9BzYzS0gwR
gFmkhqCpEi1lRtoopv7h7zPHTIrWQKDLgLZG5Abl4PBL1/+2c9UqsphIrhTmaCMEjHOst2bFCekJ
mhMZZzbrrDkmNlhJhVFYpLIsSrx7+0FU8S0Qe7vDy+CuJhuCGdy7W+9FZgyD7vds6hGemdWm3znZ
YZAYTs45cxJSLjwnlIx8onxAjJe3ZVwPQCC84dcrvMewfOTXJ4WTG03EX1LeKeLDqEBfNDhEcSgB
dTeMCX3ZhRp4a21BHBL4ww52UQwJ4WhcJsniMaGvyC4rhg6LJAXODKgypVGlUa+r9rGVyiaY7ctH
NBR6Ep8crM7Qbxo+EeMA9w5+hOGcEdmjewcHsK/kS302r7ycouOzkTamm636ywvHaQrYhCW/IrnM
ontHpTXWd91JFaznnBRxfxAreq0SQZryqjcEqxHEk9dEKjefc0PaJL7GHogyiSCNSONBrFA8hxmi
4MgherYvdNC6wmebXJmwB1gmawgIbHQy3Kgx5MGcRQcFcuT1WOyKlKlKJqNW2woArJzfQ0zp3O3z
LQzNSad2p8kASdigjvqHLkWA4zuuwn8zrfAQ0VHMnXdkGuWFQxNW5jysXQYqiPuNjuNLGp5JYsg3
PLRMV8pv8hg1vyiZ35SqjGnnwz13j2EeceaQvHmXkIXBxsbo1261dH25n5841e441UWhI41dOApf
AoFWDQ5wZgxlY7eLYI21EKI6m0Pbwx6dTGaec47/D7Lmd9LVktHfOr0Gev9F9WtbWDlpf4vCH+SP
uwo5qaR19UadDeRT7tNdl/cnn97cmqfMA5lyv2/BmWthhGMgHRFsqxirHCILMt3ojF8uSDDWJK1d
yGDkOKdSx0fbdsVWGPXesctXDocCMfZLwkiShUFZ4ngGMl5litYRUDcc6qW3Ai32/yxObYBiw18A
S10c25It+4Yu8PPfglGkm+CYKCTC+N3Sh49CvGVV04ABxrV5MqsHhmEh4/XH1xGbn8M5wnzZCQBB
z8ZGXAM+tgQL42oawN4kfvGJWxdtpePBJPVuk8+DiYKOiNDDgRKHHvHLdDk7JKNPgrc7YqsNd8Md
J4vkavISkBBWCwMStEEGrZXuGipTEKDDGAAHsDyBcZaYT9BZOyJVDp8UmaScuNQ0aWA58FhpZXW8
J50ao31cMoVSvRX5vJnjXSym7CuOLDVoQi8tSPsF4fmJ8ryF12JaJZWVTz13ZkfHrIv+wMXx8g9m
mDdgXqSkYyZaV+5B2MJZD5vivqVwKnCwTPIuIVoPnDS46bunQ4ThEchASSS49mpinhsfT7aqIo5J
DvZLQUGwk1LpS/z1O4psVWAV2t247uPTQ70sxLq/GutmQcijl2j01YJQXTBIv3eMa4imV+v2Vpx/
2+P2nTjUGjq3cNJDoK3aMWTn/npsFQkPz1frfuF+/YBpNhb1LXg3J99KK2JHcG1jjtbDMLhach6a
2+xZIGQzq0p8/o6UXJ+HWHWMZwu1gN5xbgACynrWoC1XjATOLoRPJEel96aKxaFFOqRm8SWdYvWk
zDm2iglfH46l4kjNnNc+9nqJ1P6HOFPNNr4EkTsdQiQGS5JRV8yXxVIdA8yTNLIA+Y+dthJoai5K
hshojqnTCEshMePr1upbdfifHxFbGmrX6Gk3+vw3dEzdZikOTSAjWoPAghRZo4EYCl5NYpWucXOc
52c5QtSToNZMH0TwrBIBH+RdQqUoS55jlciv1jTFvitVKAkny6/FV44F7W9MRYClePbSdtoPcLl5
tKPzrt5+9YqCiWY5T7dHdxER8EuZZ4ogo3zGjzWC6q+Ao2KlrY1E3T6PB6ymXV++cLdrdaVOWTOW
z51mOuWOBne/SkfebCv4fvxAkusUpJ7UL66h/VzpDD7RklZP6SWkM0yQc0b3w9KYyrwi+3BbI8Hw
Pmn1OQJx6aqNUQLt89IKK0wSwDu498IetrJJl73k6jN1cvk8UrKNbOz5jlph9fudCXj+q1bMTktS
h1POJqviC0ou2GILIzH1Ooxdcl4e+aAsPS4rxGZMMwuxGdh6T0UjbcVmHETSj7sS33f6XsuSc+bT
JYQhdB6kEaGgGktHOIeRyKw7T45FPGUdBpq63DIYh/nKTestn/HHIUQ8Fg5X21MlsypA4/AfZwJs
TkpWF2DZBVq03+YEpM0olKKpTJEb60KyePqM8OkLRGQl7MT+eOXaKx6oVTmbg4WL7NcfHXObzKEK
D6vQmuN/+O/6WF05g7G1IqIMOvv4Lal2xz5hp14tctvmwvYXQTeVFdZNCyoWbOc3Ns+YE2nAHhfc
CegWwfDyXeZokwtHbRGNFq4KpD4D7gh6MA0yRpj4TGSs40z1+ogi0+HKjViXEmWF+eO+hef1hc04
rbsJCBlx2EQRFYGRHHl0nhKsmV2EIAlZYT/DJox/HvsrbwRjwkl2BtTfoImaBZkxSNYa8GggSjPy
i0TnKbHB/tJLmkYOsLIKTr0oQ5RD4HJPF05Jeu10D4lRMQlN75M7oNOha26HzD6Ot1MwQP/7Ksxp
mn1DvYz6nzE7zXKBONJVSIX6LOv961WPr914MyuSkPeeEjQuMsUIf2FrUZW3sL97BT4IuIHoP4Co
oZL738nR6YAx+OHIBu3cdkKCRu4ndqqd0sZyW1h9vWExOsPw7r4YN/mKNrwHZ4PWRjoeKLwE7eHT
EA0Tl7hQfpUpR2x/KKgRSh1sfrOzpCk8WpxcIR/zbjAfcyHaCFZ8naWeSnmV4jznPNR9TUfot3eV
hnQQ0AoGatC7Bds8GQ2dwVfDgyXxlUDCUQV+iTjRS3brCTyCNyZk7dwBdihTRMVaF8zJcMIPpy6V
05xaB2KK9OYTzxP8kGbKa/dtalHvXF8hf2iMxXcrBoKOawKwnvyx1LIsTSDKHciyQzqJvmROUUpc
FLhPhh+5uYPOwG7oWjXbhcaPfxpvrn1PQr0t4mpAg+5SKlMSI0RpudBKAXtS83Yyh7Y/Q7csqwee
g/Ai+vKZEwzxjzBm3ndi0NAHVDPlsANw7ZfSGTq6Hyy3V6XjzY+qW4IzRFtJ0nM1jBIyskiTvOiq
zvsLOXvIDxqChLaPknvSUz0kIVzsn9U/gpPt4N59YnW4HbcwWPR3vFmqF4OLg07hW5/xW4XSyREk
1qoBE575owxLJ504ZfhbzG9R4nFhRuCWNmGKAxZxJKGa8gnPQ1TOw6zaFL+k7ExLfehvIFyS7PVV
QdNDx7UhsUFkaW98hRj0olgVbta/pnlG1CpncQtT7S2JiXRfmwUWYXBvXASkP5SsmSqsu8YO/AeY
R1kK20vlHEDLqKFkX8PLzCJ9SelqoT+oh5OxdBrhUCVxkecd/H5fuOornyOBLlgMpUf5skmpnWJ7
cOnWOX3+9M4v+Br+PKuHRl3F2fWoiTUf+nfzRgX/U8MtUF+kJ9D1XD2bmrENY+/g6fgOb+Od1A+M
1KAWb8T1ikARgTip/bjUZ6RxfdX+BzIF/4UypDxBPU4vKh9P+6Siv/JSTi8tvUA9NH0lzd+SzyoW
7tL6C/FOL1HkMtW2I5IwQPd+rQPX8Q3hRQwx9KKNxiKocKx/Gsc+n1YEOKUgPRXCVHfHCWR1iXYL
rodS8nii2GVs3k1O9w8S21cDd2mWNzeXCwTbceEjGf/1GdGXCjgyROiyoWMnApqy8b6Kg6q5Lvr+
aUyyoP3DmAJG7+XABH8NRsCJAFZ0QPzVoJtVI6ruUXhHidmr8XLtVgWezweDbdZhu6UODlK4kcQL
l1YHSEutQDCf2RnBiEclEu7eqDCRvu3J/+NrJ/JgQohmQPIVa3ujMIqrltfMWjt0IM0xmD6Y8KKh
gcKERZy68cLoZNizKZg4LVXn+eeyMp3gkINQol4YNeBrVeYkxo/TZsJncaA270TRIHUuAvikBztA
gZnMM4cp8ne/l+ZjfkCj56wEi8CrZqMeGWi0sN/1CG3WHfU77q+VGEmu8TflcN/RRF02EubBeN2U
YDBhvQQSEXzN9vYorQv9nTuPZcA0YTqm7YbW24sLKRg6CiT2XtoPZSAWmZl/QHcXFDQfaP3p8LkK
iPW9/H2wyMSMDgk7XKAJ5yMOSeFipoGzaDvdYQ+O/rCzGeoew6C6vIXWkftXoqicPnTgHq46wEAy
m+Fxz894OP2NUBJMNokf2hmnuna0iSjVheRn4miUeehff7j/EdAj7OQCfBSe1OgGnTNCz6Sb3/+z
RjXAi0la8t5cKumc8rPg7zd9wUM14imh9JJHXpnOl51NedFOOXopSX0XR1d+zlJPSEZp9YrXu2Jw
GwpL+6nY1ZTP1iWq5WUvO8huSnFWgMD4+La7IicV8p2uWd1mmVHBdF9IReQzMGS8MtaHT2u6PJtJ
GndPar/FHT0Fa6RFnjs+U/FoymVSTPiE3qrN9O+9yfHy8S1uEmrwjEzbLJ/6yZdp9lLt8grc7WIy
jkTKAThCr/RMyt19rn7g0CRwkuoM4LFZfroffyno9plzELaND7vWMH1bSJbhFP6ZYmORHoW1x+gz
5DjfiDLK6VHUq4rSYd03xWVCv0PtnoHa0ZlwZiOmGeSxwSLA5FIBznOCo9arnL0YhfM5Mb1Ts7a9
OswSYhtTCIpgUCsrzJJYYf0md8oHGXeaDL+1Jyg/dhzy4JO2CxKRmjLUx7zWPYRa4We3gf42Uq8n
OZtxSe7TRKDFVRbGyxuFB4D9nqR6a2WW3ZtK5u1TML92I58srWzioP/I35Mr9f1ni5vIze0sQCOc
wSjqa912Hn4Hwmqc8eN7cJTjd8kkY8kPGhCwpXAflGVm+GKoCFAe4wuL+Kwxk7qz5cLJW0tBhxG1
k+SjaUE+HgMyuvYWE+h8IK1glXaKBY+6UcNxvHfPio/FYVDrnHJcG0Sj8pYAb2mVefLr3IkGKlOb
bwEXZNfpUNbtfBvXb2uvO7OQo5+7eNAEuDKTLStZ5GRmrP7+0zomB40rx/ht2HrunZgaHimb+O/V
t0lnrkaAeYa4WSSlzbQF3YESokCUDzXxcGA2g/csHX1A/rieK539yaOzH8xRmPyhNV7P2sgZdh/w
S9NGDRy7xNZqUfveBSbhW3Y1/yb+6bs0t5Ir8CGQn9R18P3wZqxKjGxDQ4aYC44NDZV1TKq0Q2jg
Zf2XdyB4JeDy0sWfHB4e+m2El1EJhTZjQ5SZIDOsZDYTjtXo3yMerJCwBZsg7GKvxm7OR7pfJKp9
VhH7VLsvKT50aAWq5NyIU6406g/ZyekXWMhjgeoGHwYTQ0FPzs15yxd2wvFiRYhg2nBzRLBNc3Xc
fcn7W7nl3O51RaMRFFBBi5iLD7EFwOvYQsCUM3k7iIFvm0OD7jq3FuRWbUu6MZZi4kG+HNDhkQwG
UxeAkswm7nqwpXDcSaLU4yY8361mWmSjxR/uRBt1+iRXTQuWQHBA/NVLQCy6Q24GkbMjZgns+8fN
WkVeWGuApQJLeAglWmc6iZGsp8+JGhSrabx5i82xQpiZmAgvGJ89KXGhS4LwxIi2PZ74ftuGhkss
YbrvI5Ce2ywARqZk4EaEo4MBrMQUnm++QQR0VdkeUuiZkmoXtNhCugvosw+nwwYlqRptp9aU4EP+
sif9M5TFw9DXbwS4jgaUWd3rSHj+l57gVsovtoaOoB+Ez2a/7MtWL0hbKplOBK8GmhtONIp1eFwE
qARJPgG/CnCyi368PiDo3f9OfrQKZ1j375AzQ3kOxC8LZLVG5GaL8L+YqBfalWgip/MvwWQ8uom/
76DHbSmP/IUQuON2z6I8r1VeWA6N4fUXeY4Ey8+tnGrP6Wg1StYCIY27JYBy0/npy/8horyanPOS
RwIQA3iP6UB843b7CGk2GqSlFcHYFzill3C731mQp89k2Tg8MOFuiCmKdYgfsML29rld7D82y9hv
ByBsLJFHmKAarNdLgsKLNHp9xRATHR/EdEgJQr3L3uoWoOs+MKlU+D3PdikxRqJOF3nTxwNx3XO2
q3V9MSn1/xNa6NanwXsRyG1dOqbxOA904va5B3TGFUJS+EYZYfEYdrl4wGvabWmmBcGiQBVYbPLS
eFzHUyfVithlWX5chkqXbndAIpZ+qgL9UgETCef0uDbVbqmYxKUBMQXjKa4CQLn87OSlf0tXOHcC
1G5pMSCV4KfjAN/aPIWXLKkJstt1IdassW0vW/6J+x3Zg7anG2YHd0bZNadbpxN987KkjtSx5YCt
mqGqrnivFeE2zFMf2FB+QtPeuY4//EoBMUWHGuYlxbuUsz8WLZE4SQOrJHT0j3ZOrJa0AhNRJ5JQ
86hcwxKWv2RXBVTo5mWcp44+rp5TcyoPhwoVNhlL8CxiNrSwZvCn2000ez+qeZhKOgQkO9Mhuuvi
Yv5baIJIHKeiy2/EXELdeaDD5lQPw8TEaaXbtai5Yq0cQDZU+5jlmpOjasRHgw13RmBo5eH0/IyL
HkNk6FBykaeOlHQMQ+aGiKoAMyjocIpXbJPfM0jWePhYM1ZslM5LDE471rhI9fDb9ShuyDDV7iPa
2jD8zl4QD3JBcP82ZsQNKeBXM47UsSKNC60jOk1TVAkkzE4uCB3nxVCJ7x6UQcJP6Dg/qQndfxRZ
J7oObvdyjv7Sx0HndEeeDX1/1bRmnQBW7bkmUj6H9FrITI3De9vpDCto6EuTYGKILecwPx2fO3g0
jiaQDjvYm+PleS7IShOF2qT9Yusp/8cQ2xTJplijQMQPG8E8WZVvoLGRAMtmr16LjSW6xWU+gGj+
YiBt44kebzfufOQTVsXIzr6HO911sW2ksOxNW8FzQC1TcZq7KKpDaM6gS4qfqjNxzIKSDc3y/eRC
BVnq5qD9X2UQsUoQUNAHQn4PVIqcLghA5gj3MIZAnfe3sKUPKFRMgDz5gOwoUdu7cdrVB/AeGeFx
DrfNJ2fglZkMlHBKPfIcEA2Lqm9lVcwrGEu5k1fPbq/Rab9pQOhzGpZTu0IkRi+CcyAsQIc0JdIX
21pH3eiAOG5F/pxlgMVSsmrkZrhpUkEmU6k4I/tpGHCX40GfoTpYJKB3dYUzbE803YfbgwTadWNG
GUCa8lF2Wo0XY11dU96ZNKSf8K08/qYpYq3miORJhT621WKKE/DsGdmLzdETuXyL6nR2XNLQOgwe
diNA4N9uk4IOiteny5yn7PmdtETG7JXk4/l2z3vdsVAlat8etDNSoCroFhykiynx85dB6LdIDLHi
Q5+WdsZhaIeZxDkvHl5sJ5GyYVS/QlCPnHWTLv/gEjlh8wS8J2xFrAFvKef0BJqDc7EFN8BY5WEp
o03K7XQOYkgMLVvPDULv93N+H1bnXWdPyVukiBanytGAsF0MqHNx2hvqVWZk5CRfw3wkmL9tu6rg
sBptD2acSN+Uodgftx6BLFZsV9TY9Z53axYG5DDzYtqlSIlvOB+wIVDh3mtleWhAtwlvtAfI/ih2
Ur4vzN7ozgK878IlimF41faj3Uom3e98IqJYL9MpyjHZLxcPJpno1EQdyeo9StxIifaEBk4z+VSm
GAkV5hCyJVywAvxJOFwUplANLsG7F2UeD5n+qq0fmDWKEwBwl5Rc9IaydtKPVQgbPPlwwcz5Hw2/
IEdj7leQNdMMWkdc5fkKMdm8Y0Y11pN6Fvl0WT4WTvDDJL/9dR7PuIC554akpntLeqamds9rxP2L
DLmXz25uWkM4coAkl8m13WKejwZ/GlNjUNGFfUZswlQqTFK/cflHE5GskWq2fqyBRvDMkrQHA2Qk
zsDbJfiZuuSwXR+CFwjPI8Ro7XpScekBzJGZ6bt+SSuExdsTm1inODj9k2xXyTQZLlHAJ98rqc47
bDF83LMp/mkRjCmiZpjMgEHIyhXxShi/fw1BP7AqpLFYRa1mtelMj6+jjnaqbfntEBGNMnO0TR77
gDxtoEv9SCCsGidKl9tgkLG7Plaxqv908qRNMD9dY/dM3ktqCOYAFC6zsDdMQ/AYqyfAfD+6Mity
nez6RRHr+ka+5hB3EVj38nyHKp+GzRnZJ/GbX8TLrWyBSFU7ehgHom/esNO/PrrkbFMRMg3TbrJF
xpAe4gKT2jbeMjIDOhH6IcMF9cl80gD/xuHEgx+Iy/WU3pITGWvzB+2iv0sqx0iokFG7WCg7caxM
tf/q7MC0RQQ9Y6R/mrxWexJAD1In21/xRF8XUzu6s3Ck90S5ZYyhUujGRwJ3RelE3bqzajWYxHJN
1qEdvZpyifAN8g6U9Ac1Jh4X/Xbs8sOwnSdY8Qj9Rup6eUeT9Tw9fHg8LbWir7b8PD2QOsUQ/6/j
drPChexNKEGeDqFHqM/7cqSj6WobGVarOoQsKFa/Ifjv2CMv0qoW5n4e7gTGIqfGDZHlgkCXHxa0
rG+1rdrROLDgsYHUJ8zCvqrWH2VZPdWLzPK59iV3NKNrjCjpTV75gNBjMb8z7zutD6tLKHPSDLj2
0VgvkoZ0E/nFEAVLi/ccvGvJsjJkmcaG2hSr8w2YJTfeuDverOrZGPD2B2JAU8ZSMrrPkDVWzQoL
2Sc9KphlzVqB2o6G4dg3Pc5xJJU9XPVis1+HcBb6Lk1V2ELROBNL+x5tfnQTdSNbwDqt3wHgPI3B
s0GY3tBJ+LcnR+3yQ7isKAEE9LA1ul4B5zUt2Z3MPD4eUM17YIsg3gIfUaEQFnRad3hhGFSl4Dy9
rIRq340D4HdkicB259Vq/EGlVc4gITURqA2IlI6/Oqn7/XQIzq/rmuf6QtTBjodQWANPg1gh9jbt
dyHEvARgZy9y0VcJuEoMx0u2TJwUbD1l0Pe+hFpa5kNO4LBpwvHmVTJFQPwcTwCY7ASpnWktXpcq
LmrkeOgEBhNVBmJGuZck/tusOTzBq0ER+PFWo1lOR8yZvEKGo4YpLRN7CPo2rP01ehqhYx5UR8JY
yr1RWmONAXwA7hnfnejsZRExEepBxZUKcIBZaQ05Wmpct5ykS0Pc0MYmE0JWdjZSaA/JBEEcZ+5V
G7+7gkaOCdwajQrr6vDhGc1ABVvnTAB61X+8+Z81lLqk9uhespkQ/zFEVM1phHFU+OnDpeNP5ieE
WAVkKj31CyiGGBG8if4sCLxp8HAQB8a68briJUHmSWghSniTRW8w8v+4PaWp9XYf59mOGb3rt/1A
pIpPtdDH+p++9O9yfOa8G/iy7ZEGVoPHNOZ+aV2ccPRJ5RDvS9kUFat97nmR/U65Yx7IbvbQ2uyu
n3LKF0X3s//z7RmtWOR4bT1NwYsYqkXvP98u63/2hCuVE3Bi1/NMdUJi9wCbHeAfjcKJdYn2RUTd
1DRdcETdc44SaGaLfYIWLw711PjvP61UlEvrhXyJOnwO45bSLs4m0CTOFWMZaVWrpsaH3gOzqY+s
QWAeCswZLm7S32Rci5WuQVaDKw0AQw48INrtTqbTbYTd2HEW7JkqKtLlov785p0D9pvFv5PKn8nG
oLzVIX13u2WKWULtCujXoDlOU6NbUBR/HP7a9d+bB+okdaQQhaB1iPl02N53egOzCakZV4uQ+8+W
WwBdHqSdmBmKXW1Wp76+4HD5qMcw5x4/zOFs3MtUVQgFdjQo75GkIIzNyKBQAI26TI0qbAfBWwME
AkSKcf4xHrgs2YCGumUkPYSQPDAR01n74xSW75QdtdpnIlyDp9+VOoRvKrB+Iv5hYOUEncwkXF9C
XArwIjsuuvqyVPd1Od5LjexTzinZdw18ZCOo4wIS1tXgp0afHznex4uV3NsC7laN4OGvLki5w5Vo
1OG1INnUrpajFgewE5k9TfC8GkFMPxEg3wkGqpBFH9IUogQKgEl93/6wwFHSziWR6OWK9WwOphRf
Z1ul1ztAYFHzrFY18Rp2Z7ODQV0Gvws3rkhrhVvsVczjQ+GgrHQl6+T4TXa7zxrvzWrZMK9dRIqJ
771wG/FkzQKDdOf07mdiAukrs2PMalpWNmmrYzZaaIcPfuOntKOXiEhlCDJhwZoofzuFzw5WfmCq
AlYkQQv3OowJO1nHOqA1gCH6zddgA3lmWkNkAUSBv2wTkt57ZyqM01PYYOrrhKW0Y5N7zh39pBWj
kqzhOcu5+6MSm+i66DH5zPxp5qrKzvLqSVq+75c3ppXCvt+c/yBnQAwZGHcRpWla9x+TZGUY3nmS
pzxdkPfi9N6AF58MWzp+VE8MxSapu3x+Nqlq3wklYFGOljXRWl2HHgB5PQhE8+ornLNZQRBqFQBE
p1vW5PxGr5cpI+6DUxyrGFCxG943+0quZx6nwiaM376W/aNGmmiEuiKU22SwANzlOVUkNAm7SaIh
KGE8eUS63ccNjcih90xWzgXqBUB2ENmzkp++VOcdqTPzuNLTxZKdUK2IrHq+565TN4a4ZSAwKWnF
4HoOUYek3LDNSrHmLcDUABj80W7zHRT7TeaHRVkztHN8z8F+qG1SwaLZvQLpP7OiW4HrCrXVGKu0
xomvGBJAEirfdod1UT6s4/znNmLn0WhkgYbNWnyOne169hsxooY44YOBddxZFxUjNIzYHusIkmcq
CDbjUHVanxL42PtcAeJSxK+mluAYX0mfZ5eez+88UQPeMJVR7Gb3wUwVe8jGBYVIsWCZ+EXYoAFX
8dD7rlbc5Fe1OjGvtryi2CaGWKBjm8tHPtE8xlWgGjHw+hXiMJHxYe/jhcmU01S9lltuWCbA9FZ3
v1ja/hCwKUaEIBvUd3nHmciHfABIyh0ZEgNkbkjEfWuVBXVqboJb/MtPj7+DcEWT2N4Dv/YB5yAz
AqaStz74OmMPetIX4V3eJaLUz+0TF4lB9pHS0/kue6ll/VH0cENF7N1/oxnzFi/CLmDWqTwXtsNG
LEWaTMq8fajZ0EIOjfBQ+quH/kbvrsdCukP3PP+hdMG9Hgr82SQGytB2206XKZbG38SH9VRArfZP
itLL+GW3E03WSSKLfg1UWXR4YEUADA9zDl+4kvFh/TB7Q2pGBOTpoXMftcsUbHS+h5uKUkQ5nmLA
eIKNmI2HtMqGMxjODo4kfaJ/Q8oqJeBbguWYZ77IejOLlb3TaoeLlR97JOpUMkuBwUNA+RM1Ai0D
tMgHYlCKoLdcNQe6VJTmhvXWS/aZLUgQtkil8zGQ5gBSeuFM2Z33ewgHB+CfVvThHKOdd7Dt7tD/
QmtPWuqCjbPJpdJdVPVa0e34uaf01rQBY530UovhVB9risv2iy4w2rOlBdJL84h3U9bDu8lSAm5W
pRH6tJ+3Ik6nNl77OuWLjJssMbVORH3OtKQTh+ZQuCsl6xECqKUGVJerTxKmbrPS0eyhvrg8VUkw
g+7YVl3Z7S0AG9OwbamZ+icFhRVQyy+jntmZqR4NjlInWIadlOVh9JIeYCjb/P15PhhWMH6/7Miv
dzWMl4r1UBWRxwTFD/2E+pjQhv+2/ZOT/2jYm9HfhdjA7/Tb0B4pbRDntICFd6ZjOvLw386oWCUR
vigrRshQlZT/g1R2V7i+24ftqO7uSENZnPVVvjvtR4x7qSqNN8FxjJPITgUoq6sJtRzb2erNpt9z
dBIDw71xfqCPUcqP7w33aLLEXR1CFdB4ve8TwoqmWiPfZDD7s98d47p1zHytWWZp3seCer7NcpfM
zV+PwcM+Q9FMDMKSwJMGe/OY6KLFSnkJZa+g6750dWHIYuwLKnb69PWl/7iYNEE7yPMSP3IypXqq
LGUJ6AH/+U3mhJuzm8Gqya/OadeXWoTJVcOmYjcQJNXQxLQfstosX1L5ODzCossmGaFr459kfaek
MqDneKMOK93b7NideRvq50oyTM8RWk96WTWtNeQwZ+3k1Cns4OGkgQ/lR0H2wg8X10UhMHvRBCVC
9ksrcgAeB1uaAegaV9mJcDQTPlXzxvfxmSBk2qVBfvDPPzureolYuHXo7KZ59fiZP3Lmwe6k/dTx
1D4Ys0gqE9CdpKjT6+ZpsQZ2tRk3vhG6aH2kaaXOxquKiUhWRPRFNDk6k3tJPYz6pAJQfT9DdQPC
s2dZn5UV61lni4jAyZOW3H7ej5p5ld0Lu2F8+d92lfcYKCwoh+5hu/0qKUIhuXmEy14yAoL2yDTN
OzDSGB18vIz6JiBmvKkshXbJAPOpPv1RdlHLhl35GyC+WLdZwcgKu/3JszoCR79UhxO4yx3/YoFl
5og7axcXhWRq48nfyWG7bKsb16s7ZRMGHGCe//rIg2n0Xm9PP1o9FZF8Pu8NzvwJoo+FcAPdrzYz
RXSKe4fM2fBg0ZaZ1hKdEqatNls4r9mVoZqOOwjjPgdBbbdKrst2fjU4Zpn8hw7HQlD6Z62Y+Na+
GEiTaSNC5dZFb/q6/LJQR4r/eqhX9QqdFqXykHqmh07rYaddLveJEjcIyWmZ8kOcrLV5Uz4JveeH
ad+9vtk8yQc51HkTWujdi1qk6Y04yg7LRI1Lh9jnhxTg+O26traPmZVK2YCCwgnAY1seHsvAJQ43
ei0ci+TTfIESdEk7PbJGYLR9vfqnLlRzi4S78EUTuiWm4KgSK2Nyvkfk4ydUXWlGKJavBOs/HaJu
aC8x38S7clpvr26aNWw6uTtF82HxqvEY1zWUHsmx0LVJtuHwI+dmSYb1Tw0YzShr7Vy+kM/F8S2J
1cZDXK5awD7DQ1/rVPswIojg7gDaOjBxH+xdNU6m2x/dwD4+XlDlDPRATFCKcyksZ/SFUKY7wS3M
3CUb3RZikFmO+LduuhCt5/wZDa1tG+mwUJHPiUZsemgBMKhUFcrFd7h0PNWRsWQpY0T7XEeHuw1I
BFT6qX42x4vUDDeG815BhVca84DlHR5XHTYvALsqT4hthh1J5hPuMgIZEvH9PPbky2/eAHA2+q46
bLoKmwnVcODZD6sfxOtTCb3Q3cFAEt5ELlRut2cnVphuI9giEx/5u8Qd4Y2lnzvljWW9ATIchXQw
cZuHfTr3htfN6fpDlq1msIXA8h8xeQpYaeVYGXrd7yjWtuCxp7xI7zpSnYWRZFEPkWhiKsYtdfZb
KQ+O86IlJJOXqrUOE/r94BLWPKJtNwwG08fWOBK2P/Bs3XiW128+gxkjCznVgAyUS5SoByz6JFp4
Od/lj8f5NqxGPOH0mc+Mf6Zt1Cisw45u01dYLsVSBO1cR3UcuVXTpPdpp78ihZe8Z22qK3oa9Isa
ktwnnAwtQextK9/HdNkKhApuUSA3leDKIexgMDpEMyiC7xfwQT/TM1nxxPDS/TD7rb7wAUdHDadD
9C8GRWdI4eTWu539bJNkU2/OfjXwLZ9dUNvKABPFmVInbFI7o0N2lxgkhv6dYLRXAKnxRV9oy45z
qGgDzsifpi4C+3nY+veBLfAo85HC/48StbMRCkTD3luTgZODlrE/ph+bJ+Jqnskf8tVWanjW8BmI
UvYrHAC/4o+3YXIw1Vwtpc3n6jellvf1iGB9SRs12oQCD8VGTDn2zRk4pH63iDykGavLUt5oP59i
V4Pb5Quhv4bkayQwr8RtW9/YLwc1rJVtFevJSWYaLTwLrFwUnKJN8CfWoVR5hLnWoYDoOqPPRWf5
pFLsH6ovktpBmeOHhntBNHxGnmn9SE6+XRwi6R5KCrBNWfZkXsKh4uEo7Kpck4OnN2Ud7aDzdk22
P73iBiJgSD7pGz7UnSettUO1s4fTsRDL0kYskWDn/MPC6OmqX4myygR88af3dsqVGDe8Lm/LaklF
iwCZm0ejAavOYgrBL/SYtZ7vrIiS8gbPG6zPw2TkBYzPTylm9B1qP8S8XWSEmukM03DvDZr3cS8O
kPtUX1EsfYBsPaCa+/GHIkwYxn7PqdqU+H853qGgl31YjsDsDWkheD/hsvIw3mKAbd0WRzhUhnyS
UjmgvOrPiAOHyFjfZBS3j1l2qy8XOYoPShclEZ9nkf8LDYOlzKDW3QoIg3m115tnSDO84qVyE+VG
ugyqjFYnz8I3KBG5whiC7Yr4zls66vjJs6pc78upgH20uM5QJKSDas3FIwYH1ALHoSIeamkMUSrq
ZIk7jQni8yFdxqOzXkO+TR4guIB3heoGuIBm+sVjFyqCvQnsbTEMKqIEmh8FHKWtLIcLmb7KiejY
8swxNGTeTHuxCUtG6rTjrQiKnI1Q6DvAuAHbYE9YiwDh+viK9I9VjkMTXHltKPOxznkGQF9CGVaR
e1w5d/5lJPPI5Kk0yIFEgdShkRTAp1onvgIn0biJ2u+aUYbsxAUcZkD9zy5pboQ5iyaVDjUtDr/o
X4wESa3x4tM4DNrlVHS7h4jEMjBT56eoqOEOfWFNUU6WJsqFHtYjBXquceWoYjcD/SFhFxxiUr7q
kI2UytpPvhl7NQouUOmwNiuiuZ2yDTU6eD72IBq1VgdJbXZRGt17X9SP78YuKT9zPscufYjHnAU5
H5ArskP3CW3EEc7JBWMVcz9iM7C7CSQY8IbeniDC4BB+xLOZGThvrlathLSoxa7awr+RrlqIqtO0
0t6WA5c1e7uJOoIubaOYkKwVp0mkruopk8nik2HGUaVIXdwA8DHQBJgqD7vVsMFEq4ynBgC5gu5e
++3sFM3J3rWRrRR8xLOyq/EEZVImxXHVRCcHhMO54/QRFG6BHY1PRQf4IhejkaZUSjfilrMdCklJ
xkJe08swgUvLKNShcmqOuIDz9pYJSETSGsgoLB7utHmodbn4O4wSGHBPbZdUlVdKw63Jmq7Lqy/r
fnuQGYfv73KqV1AXlLzfUXB4vfVOhs+Q+1xrXtuldoGEX4QblbFSCTas6Ansm47av6lrSA7I0o5J
kZWWLNil8Un2f6SbjaQ6KP5U5XC9HITHSMGpXsgt7bIgD1xDobsDYgAIhc4laPR4FphGzFEcJqJV
MxyoNBHioL8OaUQoi6OVaUYjMSYFylkUSvqn9WN69NUCwmIrcFQezxTS5QmHbEKw3geqOpCuo1Lh
PYMUA/hKw7r9satWlRBDFuhIp0EkFSqTPnPvJb/cHmLfikfqCKtOK+2dkkw9FsRpcRcmFHInldNB
bjfmTZcU/DZP8l2UGGF0lxxejbheajZTYTC3VnF/J2bPy5JljEwJRozu0p1O7N3hhqBACGkpP/T+
T/qrJ56GeVmrQvhGVRnJVxZtA9UweOya/SFC2m9rARJzWeD6rMTshmrRk1KVtQNAREFWhx7uCRYv
bfFTFBbtIRELUYj4Ku6FQBDBXrduVixZzkXJZLrgcbREmC1SOfh7qH0EX3MHRPg5e3COoFTvW4mV
14rBpyJQsCR/A9mBa+3wLQtONvcOZRHls4qK1v3hBkjNCA7HeijwqZxL9h0G4dHkb1YsfTIW8GDh
Z3teUG6761YM9+gIwVT2ZtmovJdbXLWKXtwli6uJuRm/jZvUrSntCT7k9yfdFgkumeooeUUlm4YP
sfPLHrAw6YACbHgv/RqbgpFDzL5rgegP/NfSRwUXY8QyV3OSUYy93F4lKoQ3+6CzOh/XvVBtWQTQ
RYQprtGVdzXKhDfTGB74tpbNFLlCFDus0qEXuWmP4uWRCOrdKVJ15VW/nLtJDK/fUzEohJP8z44k
g7pdJ69Z0U3hOwNoFngKRU9nnSM3M3f3A2mTAjSfBc/qfK/ZSgwfQLhXHpzOcDDBAd2gygdhdzoz
HISAvJrZklk+jvWW7ibr6G+7e1kpz5JjJkwOSCSfgewyg+BmrRPySjpo9hNrSLPLzkNVvbZNvw49
wy/xVlC3fwV3BkPftkydN0NkNQ6Qbs2H/1icnox9CX9wM+TwWenv6W5UCOAKzrjJcjfdim/t2F1s
VjL1GiuHDNvFAKZMbLY393iu89AU4GmdhSGcMW7eoU5cvht6pAY6fyOSv3uLdaVNCWxb2Z4X9eL0
ZzjN6vUTjhNSUzl/bNQpgRY9bGt+YAj1mjseWyrZwDPMqMKoNwGXjAZ8HLgCz4vGOMSqTu5u2I/U
b21UATpSOkqHDCi1pVZYFqrLCvqp9JBPWL7/G+0uZJyyvmWvR0aQL0cR0GWsj10I5y/NBgiLoLo0
k/x/6vkLNNLgPw3l+UDpHu0lsvKsR/pCmXno0RKym/sfEX+XcexS8K3FOZbUnHkRXv89XgA1V7M2
jD5meg3xaxJX2cQ5pAW+EhvBoYW0VcKo33JYc8T2x0ZUbaI6ePnnRkFbEZbLYUJpvvrX8+wvW3Gl
zPondMILr+IK1GA1ldtVfWDsmqnsvtYj4E6FHRY4MQHmxz07H1S2fNYXFiVvtFvDR5sj9cFJBcSW
bKJhPAyZOGbXeQaqeFTXBc10ogAXfTQpOgXSH08TqqN66qCS5zEplqx01+Jh48Pmh5MYZKSiT+eW
65S+JG0elAY/uzXHeCN3sQJkd2KiRZFgnumY2jipMfXnOAGhIMuJTO6bBPKoFrPUqN/cHwJjlHfo
RRl20lmxSCBJEIVOxuoxv4Vl16tF9AvKyKYicEGn+XOeZJ7ji/1dpsOjKG8WxjDds/4OVn5dYlrD
ebosq+/DAEp0s6NtoSnkAB7nppGPHL6yCNJwgfQrMwoef2WzRPZLKFnh6vJMf8wV1NtU9Glc2FPY
zUInaF8XB5KAKyF1pw3Xn/s8Cat7g4wrFk7oHvood950PczMwt0LOrrTV0KB7TAuIZWu/EuXV+CS
ZBJOUa1TxsaVunzbXRkKITc8Bs0VJQXwOPVq87O4V2JvqR8riwkdKMdNzLata8hzgIOYRImJrW1o
dXkm+pMida/MPq8hXaxQ9DC1aAM5m5Q4EgWsSqwn8SZtUXi53Q0UGMI9ZsTUFB9SHJPwzKmjLQyv
YoiFxvC3yb66gS603bxayVUeHuk/og20LKooTMDlC5LHDfQXAC4Q4+PCzRwGmWXnLUFZUHhglGuC
JLqA4Iq0MPEISkcnUU1gClvtubPtBbzLWn8x/5IMI419tzqLhd/b7MnPRuQbrRnVSlMq4hhdGJ7R
f0pvkBlb8ktMcGXtqUmPZR3KvidUzA2AWLG8r7vmKgM91NjrqLGzyEMsSf3VlUyOX67GAlHtfcBE
vIhLhk3j3FSlFd+VivqyZJ0LuPFmtTYkkhF8q5Wj5Oz6gllc/ou5MJ6lz61HAsjN/fJA9bCDYhqN
aoV41Fr3qbMa2rOojBVqghyrWZqzYwCpFOnJ/Q4F8aBYa07dkv4n9XuW1OVpa1PNF2t6T/hHrnDu
HDTyyRMOqqZ5FL5HXxQrhLBd9Ggy+M+K8eiJTi4xE6wFB5NqolHAWWC5AtKZlOR5k3vDHp1KRQue
OVFsYyM5CikIylo4ARmK4Jban4JX5ToIwgVIAXBmQxyXuwlHnGSSYGXl7Zq2dR0Xbr32UJULo2fh
zLfdmco1ZtLQmBn4hKxA4smN96UkY9HsMOcCy+EYI9HX1kRrBkgJ8j7XGG9ZGAvwv5R5F4QNB17r
KQdwVoPHB0N56ZnZZjBDusQQjyr+x/ClFKqhjkDK82Tq354s0WLHtCBbZRitYvVel8zIwZibmUqp
jSRvg3ow2TApTnJI2129gNcWAOXFD82zIVdpi4eonAa9ShKvQ/xdQAouZA1UTWBMKXwbNveOEByd
fJm7MQuOzJekGwu1ryOTEPu343BqqgZheQ75eXmomhGvHrv/jou9VjReMmdKvkU3CxyJleqHf5KA
8E3lLXXU3a3Ht51Ytkj18stsXxSzRFjhmcTlVsdMQGHM1MzYRp38wHyq8GWDNN+6keYzOs2zMQH+
TgMgugpnfmwI97Mth5OexuGJSaDzOzc38pESHn9j+2xQxRAfzRY/m5ZXbUcRjWFX7aKjyGBFl8Ef
Wf3F7CT/XgRMCj2oObEV9Omv8ChBNnQ0f7jmwUDwkTTjb9Zhtu9EMbIfMNt42Cs8g+odlwXq4fQc
wKCh6m87r5cb9OsxuK+wx0mWfV+iFceHHWQtr7AX6ItqhTbW/NYF0iESpjyzAMtNBJU0zDl124vv
ufsxCx4U/MU2XaU7vaa7/H7mAaaDK+kijhkJsQUO9gCVp7xinsRoqQ/8jL09yrqTa52u35GvmeHF
abzI/d/JGHVgmxbvSk3nTU6/mxqWCk4fxxIJzPAWDXf0lFfuqSyE9bdplFdbiabGsgqdlYgUX3EI
/IxUM3j+wNLZl2nr6MOeXroLmKLy7APvlMNCGbuOuGBvinKcHW44Man2Nbqnm/LjSz3LbSbgUh9Z
sg/GCjdamQ2gI9eeHqaJRAAsDLtVsOtqpyo2mAtio05snbSk/tGlk0DGgeIoRmxWhzwLW2AO1gBx
gm6CoA0CYs1pZ7pKNmojqeGQ6OXNg1oxtWeSgSMZ/DfOiUvvLVNM+B5W/l/yrGJdTaL6nBZyE47w
iC36GJdSX9/Z0yYIsP2N9iakSRaxlz3U5YKptDjDCnssccny3speC6oL95qg+vc6Utw5I8Gbk+Ga
ddUOICn0oerW0Ax8zvEcF2yCEaJxhuDCnHm6A7ERWjxQJsp+ZbYZtzxrt2afd50tO4FV6t+SvzUc
kcsRSU+dGIrzUhk+ZYhd/c/J6V5IF6ADLowMJ45X7815uPtvAPX34KQGY2PmWSuqwNJLV55m+zIS
+FtTMvwv9bO41B1P0g+BvoeOpam2LpxQ7DdSmRVccU/jBxGWoKCoL4eJaFdHnU8LpOzjZ1Z1JhmB
zAI7iqrIDnAVMyXZXTofwCivYTIAokr7Z35mRejW6Q41YC8M2SGBGndaU/Jb6T4Ck6SLl5nYXGen
Jlhfarc+9Ae8W3/WNJ7DhBE2FsJFIdpczGS8FfEVOoJUYAWFS0BRtbhVowtRA0dFvpK8ZBhHaIsi
KYNuZ4qwPvWGXv5mBsq8QPthrg1VhJHl3WpylSXkj/LyclaKbBSqArrCdgUesyD/X+XfirMozUmd
E34jYLj9ogODgeA3L/Clhrn9uO+7QZoFjDueurn5uj8yi95NF/crtHbcEKO1Tng6QHNdtKixAIJ/
ma4TqRewV7DrmDG/yflN07iQeBqN835RgBxxGv9G5j8L1otVqi6Vtl4XWeazs7Y14/Y1+awgkIyX
jF+BHu/0gS+unjUNKjdNwnIWyH+H+eL72dI4s1qxFHMyPin3BM7N8BfLFfKzMVxQCBR1QbIlmjYU
e03rny1iPJkeXD4b+yVkaMoE3GjQz+orFUJfa/vB0VXQzX2QTWGkTQBvNWM1PGDr+n7gSwKJ463Y
YFPHfsCbK6LpLAARZY71S1tJBtbHh62mYa4RNOn7rSpWVARLPaxd2qunzAaoENjrw1dgP9R9NPUT
GTXeafUkz3CmnvbPPY4CiV9Cp4jbIZe6flzhXrAam2PS4CH3/HMxaV03TW2FIRjyHzigcN1iA+ji
/5g00WtEyLNEKUA3IBasUlJK4qkRWtGtOsszCXADT+etqxQhxjig6CV1vdITMox0jFnngG+lgMEh
f3u8TNb2D8Hs/Cc52tUFufIA/ufnvw6l5hJq7JbW7c7OxG7xU4HpkSOqM9IALRECO23iCTrn9Q/V
m9YSMzCK7iLS2Z7XjBZvNQQXG3JoMfvH7yXV8UM+hSJ/d6yUOan2jtu7bxEd0KAt/3BJXua8HfXg
peGTsuRvZTfD2DzcganNQLmNUAXc5F+GELY5hCpfvKkCNctznDzdU8Qph6C4JiqCBiXXLukbLzi/
ePK1NQYzQl+4P/yF5Vi8PNdm18HWVL/10Ju/u+22TPaxrXqVb7LJA+kq3z0RHkle1DT9V3l+4CMy
78B4Jy/AQ82shk+63waRrG7CGQmOJ+uHtC07khtU4g8omTLwcy9id2SJQ4UUYFKap+czrKiuSEM8
0iomuCK6aFc3AvDRBYGAjftY3P33l5hYnBEimBpjc/ttAOqplxpc1c2ID+xguHYLDlzOc1tDUD2w
Rcz29Kpy1c1mvO/qI+ozh47STDtqjLFZ5IFuE2FoTyENvbdg7Iu+ZVUL1z41n0agwFXfI623aBi3
zsQuOtuU6bNrX+8mF2YS9pPL/wEFefCh+dgxh9hiVIwyE16IcToNMFPBPeIDbDK2aXo2v48cEAQs
BI3ArebUqTtkTHyRQ1OgcRq2zOewFQWx078B6h990ZqB9TAPQ9YYbmmj0GDwJbUjgWl79Z49oRSm
2hHSHE/hXYZJaaOZHzm3RNovho+QJqp/avUD8zWWNKeG5BDEqvSAAWQ9cgtSkdVnl1LmzZs5T8QV
r/YweqRLSLfIx1Cv9/0HUnoZmBkqOcC5boDYPC6aocQr/Y93uFfibSYLzz278NoZLBWSpedNLtNq
Abv7bjvEvOlMamrdP+ypf/wMRM6BFbec0mcr97cm2JqizXvfdfsbkY/Qv79cq+BkonzPMtysj1Zn
PX971jCUdlp2vp5Aky5O4kjb+ZpMnMu+ewZANdqtJb8Uj9XuEZvoEAifLjJEh1K7bASFRr8i769q
BKnYotSeBsPIiwsOZwlPFZpiCuOrwKZ8sQk55pAuHaRFk1EfyElbIXDFezXef36PZfTY7AZHBqfx
3I/CNBScQ/EGoF2EQMYDNImISy98X0gsFFbg1IhdRxzcWyzz8WYxLg1s1f/hRYAJwRRy294+cpjl
+v4cxPR81eaJ5+0MMpx7a2mlXcjcaVkQj2DeS+KDBT+AerqhKbgYQlQMYdmDgP2tVYP+1vYL/rKt
cRlHgtzBWpDiWFjTacdNk9I8ckugJ8USsiOzj44t1Uk1XuVL7v4dftExnW58iRo8tZUMPDeIP7Ru
R9zm1ecZ7rjMddk/7D/fOUVAz5LMOrls5FuNkVqx0b+R6X5vhk7+lUjdoJ38B64cLBEYy88e+f9n
vCBF5PS0iD8yFLLpfb64PrxNhq7vL9s6dWSBIHKDe1z5BT82IT5CWrWYEOQakSr9VapWYKI8xb6r
h9a+y66CuF6G/36B4V2aGOZm8hNifheZ/NPbee9dqlsmAuEtkd3DLKby8BXAwXQdNgLcXSmWObv5
6mA/rHRs4ErZUfQUNINz83ZxySfzJH8FyPp2StUzGnMiPMHOc2PgEprPlqWZ5fibaRm4psGDyNM9
+lN7Yv2F/EpRJPZoND6VYp8egcKarTBI2fUkr+vjX50BuE1l40ZeNvJ0K13DVOiTvTP7VWp8bzcV
3n7n4+0FnoP+x3rUHstQKqhjI2Vm49C/nzUpdAUaAPovsOD+B+bGZEHmYK/DoQ48ivylrE5UC8bD
ObxLBxU7jU+VbrQXTfwlScAFdF/Mz19t4idGdmNYSciKaqHI0wZXqsWqQ36M2ISe4kJ9UWA1MRnM
syZ1oolqKe7MU+mJ0Fj6h1JZfHj7SCte44lFH9Lm7y9sy+D2ja2Zt3mpe60endxbYFs2eeWZulmE
SkPyHJwB04oofOtkt/G9+XlDKIu+E5MgaFYaqpXO5YQuEVKkO5v9vxJI14XRhsk7bO5otZDVqAxg
gXElgwS2LEt2XnnL3fdtpKjzh2TkTneVOzjqqw++lgzXChEdzftZlP4RfTgaiGukuUlsfnkEC9v0
8sZw0DWfe1L2zNxB7ehqtyvyiOvBGYhZ9FpirD6c4wmSs0r1UewzSC6aclVgoQsr89S9wIxoS/vU
PeNZLmRWnXF/vIIBKpYWFP/S9LwGGRhGB/pnD63eDh5Ke9R+WwigsYeYlAPb3SgfByrne9905Vvu
Mg0r4BVUoXj0YrQ2t5pABQgqBw83/uRHHe/WKyHHDVtUAEFJ3koWnGVf0u7LRxVtfZsaxPOokuT0
AK5jBErQNuqNKwl1H7qbtvjiQzfKNeAgbSvrb4UNLzQVON8F/iqwmhJfsg4TFMKsXSeSiO16NNqH
g21R2bYrnNQlE7GIR5OO+NWMED6QPb0SADePhC4OJgL/OCn/JBmjEGZ5UwM2RbH8ZTToKYMLXx9D
rq6NlPf0Cd8Qvgy2zJdhKORMWn/0CvIEx4usCPUT2wzWdPLbGl4rNPSlCVm38nKiPmvyoCyMwjv3
3+KeHBYujZsHZhZw0WgPN2ddt0x819pu4msKf71QiiY5VvOQJOXMhcXJBliQpuZ+j9NHW8cU16FK
0E7SU2IJDfa3+fxGlZGOewoey4Sx7hWT5N9co1EwY2UDYnGMYMpebB5hXEy1/GIk+t8u/7f0zfef
EKQm27R8m5wlUkhqe4TLLs00ufPd1NB0Ehqryd3b2EX984yXjxQAzm9SWd3vNWsw0rZQEQJIEZz6
hAcuyq3NxX/JBkq0xNQ9O+2Bj5qkY19Rj7pvtc+o83GFej7reY2F78qvICQ9m1I6ju+YBueX0dWy
wAdeAJnIiFZ917IhaOA6hdkMdbq+dRw0NBF+CXof5Tz5f84qB0GAbA/PO2hQxNE+8zwBhWOIo0/X
cEUcDrO8tyL+vU0WXz05m1np7BpBovFw57etI3Biu6RMIxxOZRQcJttt11RXTGhr+j0NoCoyLrca
pZwXAPXfwMe26aAFRGwPdSzCUIZ1LHfwzqC8ey7iCKouiz3FyyTiOwet4WdeNp+CNJ8+Bl2+lhPS
y2vmLOGZ8vzTaR2gmMZ9lN/PVY8kb6Ow8a56RQcziZ+i7Oj3BdpdR45KrdWAXwl9KVk5R0BgI1sL
Q/aTJgl4NvusaCLKRoDBZYlBNEAZvgQEoINZykgKrUKXTNNADRkPD0PUbCBHucMANcLSIak6fESG
V25RkvOw1suXOCqRGzgn2sjrIwvk2qKhQNYm0rY/xmcbWxR+WYD/ytr+0hVrSFkEesreEivm1OgA
tUUFp/xf8IDj77ojFCgLOAOCaVj8naLrOjhHb1c7tFFPgzna0ZDVH+GmCisrS3Nreve6LpHs3S/+
FOlrB6bOqsPOur1V9kRySau7j04Dx7JL3p7d1BINodZ2ilEbdpIgcXQqT0lNbNiYp94clF8ESNmE
9WW+e+gLUoz6DC/EKwfd3BmIWUH2TykQN7txPNdQf7eH8ahb1OfCZG40JbXxE9jOaU8VWn5ZkCGi
1NnhL5RQFY8B7ef5Mspo7CDNn4Et9sPFykIlkC0URxc/9sTNg/byVoUujKdIFom8zHn/me9B9d5z
ppr6zMnfwMnVHBN1yt9Dbq/gfQodd44pJ/Yu4fY9uUAOrMM2gpLXprw5rhojBjBo2RRB6SFt38xA
WzsVhxodCm2gAfMLjlsB4fxdHN9YMkp4wVR2XqmjT2Dvr6DdZbOjnXikWOz4dMooQ6jpoer2LzhV
UV57RL2ITRJKdNd09a+7tzNq59YsbYamXTC1LwP0SqjFhNwfnq2O/T8lpBhX3IylrOBlhqSoe40S
NCNHEfIRPg6LjnrhvtRT9Q/JNvKguT2sJ6Tu1w4y1VDwyGt7+SWTkKjNSGO0LwYSTYPYePRQjRoM
IZ7rB83aKxG0beZIjoJIUXXWE26N9K184i9T7jhIgO2HGMCm8sIcZ/1MbCd3zTy9Um8mdRn0ZnOs
6L0SJyH4D/AmLoHODuhUof0ETasdVGr4L9moqczjQX1oDEzDJTm/yPLEqYPjxZA9CVK37d69Pihk
lnvTa3hQ1WO0UXP+i1fRgBiwRacmDG/CUykHPw+XxOeFQT4rV9pBQjznz7302yqx9p85rGL8Q5dr
n7TX31U/N6rc6Rod3M8ncw1CkZ025oXuqMfG/qaNLvw+FDOVJJrAoltx1gN8NJP4znZvVE7nUT7P
lEEfAmozTrVJYWTR7LzS9exJnq/iGn2T9g5tnYmlp7MDzYDnja6sHa1rg7BLsxG931gOeL8h1e0k
W/BqBXpMHmRWEUlBwLd6f5leF1KhUlsFB3/UvJFH9FENPdHSwFrsndqcMTVLJF2KT3t/mxH9uWVy
fVhkKYFOZMcPQCJLDrlIWzeI8WoQJcS0R7ONIOeAh1HOtqXoswAvdoGQiR4XmWQAmgkli15A1Z4r
boQ0z5Z8itzPewHG22q8P7h72kF7xIPMgX7ekQnSju+NJNuoOGJV8utkJmmiSXkgpT7OrJr5g6S9
zs6yZawDzJvClPCAbhHz/gP+Bl8p91PhTMHp3IhZ751mhEYoL6TGdRjytA4vbM1yrfNSfQ+KjRQk
IGbeODKfhX/0ALgKvVrl1aOUt2GMuXZq5bTFe/LBzbERb65yCQi/gzLXWOca76MAOY1xwZBApt2y
ZugHYhXcI7cGfBnibR9SVNhEdvleYf/WEECdssiPoIyLqGbq63hrMlKmR7sQsuFh4coSccjPjJCV
6fZ+RY1qZzbCv3EcKYXtMiMSfE+RokW0H3ge8Wm5Ttrn9yCKQaQGvu00j4aDPcJ49MgKbKylW1oX
wSEG4A01m10hxTeEO0Lqcyd+A1eC0tSW4RQZI8nCJURJyhJSeKzgjVeWQpR3cW/UhgbF3iYWUZ9A
fLHKn+k/5/E+5MHswWxgf3LQMZRXS31n6mCT4Pu6ZVV/5GyLlcrz+4BM/GaOvjZB4MLD+jyj8oiz
L8lqFFw6cxT+9Ryj9U0dwuvmwKZ02P2Y8d9kGv7fGW1OWBkXCBIopD0vHhL3aBI8vdH+apO/550V
co6P+53LIuoHjyq4u6d4lUzofX1bLg/wpcVrHNi0WGJLHh8Fv7bBdHpJW9YdlOBpLzL9coK7vWJD
dMfDC08L5k/oLNcimdmZsSx2hXIhERExv1C5m662H9UmQoLj95rXhOP1+AtAJX/5hfDLiuztV9HW
aIfnIBjwbhHJMuldQg1P13geg886yyREyYQn1J4jLJjkzqAYe1+pLtPdYX0IaW1f43XgXejkg+Ze
kCq2jn9M9V4ng7XY0ZX7blMd9/NPJxGuge2HIHc7uVx7qKyc1lwQ2AaEV2cmRczHiRnEFC+sEeoM
h3QwR5wBwqX6B340cXoJqI1VcQkc7zzTPPUTKqKC2aYU3I0S+59tbWAlQJ9Sl16PH0V5yLtJSrNB
EZiRYmJbPAB8t6J3VJ6jpcAdITnmdtBcCUSvUQ1LfLfeMYAWT+AKF4d5wZ15HDOp736Jc85vENa/
ILUmfyLpcw6j+ohr+scp7qaLU7OZ1AG1Epe3p00y+5NndKQxDWGcvXx50BCCOyKL+xd9YIiLB+ID
ohqjaElVn0uP7U4rCErpmiGNnzH/xhdGW/ZtRQikKYmYNXGorYKVBz6MVX9M78kfZU8BPBmkUXn/
8c0xumjOnIAZaFpiznZ+NHC9ESfGlDVu1WZ9X9DTuyWE4jO2xe2ppWj6lC0VYynNJ92g9bzMoEa8
h39wrjPjZ3FBHSqzEXsjByqjrVtaCewSS2HR7eI4v+4MPUQGH3lUfnd3FpxNf6CsFQbZV7VXB9h0
rwVLojiDM05oTNXYb2JnJGwsHU/JmOq+vXAM7UFFlowpFIQvukBBJMudP/p7F7rrPRfx/eQ3RLr9
SGYcnSdatNl58+xw4Dx890o4+favChhYmaWd+2ufKcSMPhp2NUYVeTmEE8ic0VSPb5GABf8kKz+h
WwiemQFtRB2KJvePXkxo2Dz+ZZxlTqgv2Eou2TbMfhEp3lfNBCawSFGZE9LqvrHasW39FY7wVWVU
h8ZSbr3YoVTpL7Omu5hh2M6O+fpZ1ZQ43hPlBKba9AeumZez2yvTe6W2/FUxV4NGnJFZHZ6pZHID
ob30W6EIpwZwkzTFATcKz1Co0jYk9NfvpqhHLurhl3t1zQ7TMbqxGwbbr22s7dMfJHABYKDaU8Yl
RkEuwLhGbqmDmbaokuuoQ2FnvQChsJRh1ZR0zRWguCURuZW5HAg/3TricnjRhsFkB0AaSUqUiyOO
B5Z1rPYU0LNSMstYjeXmbDLIy4zMeros6loe8g6jS6Joj2mgtst6FRtZ5+mOAaeUXxRZqRTIpRzW
LPVEUDgXwozoTdHLfxheLzY6Fhomr2nokkGLaXRBh7vbDeglDoDOLTGC07JcwOEnDT1i1dPNnIaV
NOdpIAOkj/8GO4wc6C5jXFRVUe3k8bvJnXoVSPcytKxjUnw+OUBzloTxJZphzLY2NEXhEAW9pp45
gJ9cSeeBbXtE/bZ5feeoiAP+sY63iCFFTrpdxgTh9WdeFxQcoZY4umM3yirQc3ctnunQd4aTfAVm
bTA/IE0VnC7o2es/oJadFQfxcuQBYmUBaCq8ouaIT7d8QNv9dL5uyaRwqAdIGut+9uAqFAcEu89/
bnGUhjjrI6GKp067BciizM+7MqKo/Egq5/hVrukATtWHaC9thfEFt1ieFl4hbxJUyGlo1cXTq7xh
05tVcAe14UD2teqqslW3xG+Nbj9JnTmKiKArMlhkMYNfeV6z3W1kVYmkKFifB2dYUds7acssc3zO
/QEGvyoEdof94j9mI5QS+tEO6TFi8qNkKxsG/p4u9cDP/tgk6l3qhuUH8r+HvX8IQaZ1vHwnbAQ9
PyL9kCwWL87yQFWWgy4vwZUtb9FMr+GZ6jeVvBcSIocLdqQ/Yn807I1XddXJdH4XUvfwtGBr2fIo
vCTHp/jvDBre+ct8Cggxkb4cbZ+waiZV7BALIc8uo58fVTZvjL5aZUtj3rwEifcH0eh51BHoiCMH
UIVlHsFN7krGGzZLc81OA6Hlw1UzKANFvktCOmY36jRBAqAmtKOIjDxJgoGnc8JaYx27YRi3hfgl
Dj29mOT19w4C+ZKe6muI+EX7K7L0CmO46hLI82CE3L5BGMHn/FpTb/olj2pbD4f+86WZZ+OeBqg8
jSnxfbQZZ7lIt7YeBcT8lsK6qPO7pOdsbpVLSwWcqivibd/HNRcChVCKpXj8DGCAX/3kfYDj7OdX
MP3dR2Na6RNw/kz0OkmLmuW2buW1ZmrVDwRpTX6jljVzgYuimpKW4oucp3jLOLNOc2YcG60tWHgZ
rcRSRU2F4y+RQ3nvJNdLOsyQfOogzEJDwbS7jZC/9XjbiejtvtglOOBbtXK0+Hw0pm6Ry94OZ48V
m72SqTkPke1S8hH/YJekC/XD+iLB6uRvh6xszlVOS3qlgQ3YHKMc1LdFi9tbbNWaDLnrdoGChm2n
bNaMIm6uxnuFVotDcicDj4G2buKRuwUFqeqeFBcxR0mI6HUAsb4YULIOJQs6a52k4xI7rHORxLdg
USWlYpnAJ0zF+OIZkgJH7bUtONLzwR0DBaBjtVGv83FedYRz1Rqrzc6ID+exzOW1TRgJuUpehZnq
nYtt0Rkj86I168pjwi0HAznjBGUZ9N9LiP80hKCtl0CewwJ3KjrGCMe38Rhntdv62MnzRbK5sVgL
yW9iJoeDAy8Ev8lu7qiPJ1S6Se9q7wqcFJFRGueyMPk6vzNs4+U9hmsdDzHxpyt93i07YUkUwSFt
1XSotpk2ODQtrncv7rtIkZIRb8mXLbUwxl2yTdAxvWs1xhJk/mlo+v/0P+nr7+2P/Zd9Smuj6iDs
N1vCg4sKz1P3PkXP2j13i8nGicPhk/ve4e+7ezoSTqD4fbsTyTq2EFWLMYqu++mlDi3BwbFC6fZP
N9HbSps6xIgE/LHGkFN3eskOqCpMIvnYLUz4+URFOHYqsyoFo0JUrgkLSHFeTIAXhaQTQB3SbzKl
wdJWk8lC+o0PJHlmqnYS9UStnR7vAZvlz1UF+1XGNyJ9S8MshjHoD6HFQFMYO8czpo89sHNyNLlt
IFfozQTJy3bY56vOUbbwD1hXVNfnxS7w0JLOCej1PbM5HghWSHXK+eBGqlNIo8+T7yHQ+Ni0LEr5
7jm19Tah1zzK9QVWc7pbcZ7dqmRd79wFg2HQLo0mV56uMGGVHXw+AFXOHq9YS8vcv2YYOZxpBJ2y
+NT4eycSzDjxH2l4HvSR4rcXJUG+xoPfijBIENbEv2if3xgPgI9xlrnUnqDc9LafNsZZvaKEq+p8
mnSyIQhYm72cXhq5W7TAiXsvd5RzPCdiq0zSksBXMbXduEu0lQJ7W4aVjPO6iswHnvGLSrQeEMsl
q7lJ5ZQAvfQ7zQ5OMNZ6rIQ35WfaXBE3ON+w2woVIRBkA3H7Bv1xzzOUo31v0rPzXVEle8r2P/De
24GwldKORkgfuxSCrSy8ekmGep7BaVdzWTFPg0DNQs2y0AX8Kd73ZVhZdU6njIFyZol69Le58xUD
PYGoKpQlZsx/KRAN7dGog+Kn+8zYhkTb8GHeG1i2g8TwzfAoezpnqUjJM9sG3BrNc2J/TPdBW/jk
Rlo46M/BuiWqFOTOaxWBM+FZTuM7dM/qHjgHaG4blzAsN3XSJTQpsdTI7mP3Atk9+o6rNx8sJaNI
PaxnO5Z6ABVEQlaDL2L+Thv8aaB1XkTD9C4oIQgmHR6oEGJf9eMCp/P0NhjC21cGq8iuN/YfXVvA
IwxfN8FMecG2jsGSiVNm4gKNiGUuw8ITdFOCsAj381stOTdv0g8hv+TjevakMEiqbADneKiqD2M2
iBGmwEsTzS6jRn/qKR3qspMbh0LrZEk4naWYJj4q0PRJu8xPkTnmlWSG3th10+F5togHxvFhF2ez
YAJRSyohvbUdE9sa69eEctlTidUxRPkZ1NXmjYayf40zbs54T+E0R24Jl2wCNQrTxofgpY78FmZY
CjNZhvdCbVC1dpYKdmLlQYJLOL/JvKSO7UEIMvrPzBsrijJ10mW2Khwi1CKWPb5Hs68L51PZL3TG
8Ovq3OvJD8aH3JE2fUOBfqjXzhVNJrrFZwSE/Dd2QlDBQdz9kmghIqQdKtN5aYvCE96O35arXMPG
IX5mx4Tkfi0WdM8y2v/QNZnc6u287m/SOWfyIj+5PYrg7B8Ozwzth99lkK0UkzbYiIrwCJ4+mNVu
artls4QclVgAnYAqkhYi0L+MlTWQSots155SBHpeYyzCyzK4Qsk18HxAjpuI1Vb/sqlFIgmN5q9C
CSzGjCi12rCHQujalEElwGhze/uZX+yYNZfgL0RR88cBesLMH5/YMphKQ6s/niZn/lBNG/FDt0DF
GmZhD8JYOTdb8SVvqxw59lZbhKTYviDaPUwOXbcoi2YxW/49mDpU8vTkVOkHhTKSc9FIxQuotlcM
+yOxL88kgSg7Ezymglu1q++Kl5W4h4kLF60wAJ+QoKxT5sAhI+1NU1eiyhs3k+WKBF4gorMHqlgt
xiE7qWHE45CYVHxNyYrAMN7kzxOuuJyE1wYbzTNp6QKPVdLCzmC2qg3LK8zXOS0sO+mlTMYc3+9s
uvQG7xOrfn6tkqPEnMA22wrDU/uINpQuNkTS+jN8QaA/Rpobw6pFf7WJBFNRab95wNFNH353vfLq
CG1kReTmqXDlFiKpvRBCPRYAZQZCvO/izKryROZ9Y/7wQ/Znet/YYIja1IAvIrqlXij1hUgOtdE0
7yl/SAXFK0uRVG51Pg2sYbTbw6DYHDWaTbDZQOOFMDWiTJ/rd1i/Cz/E0YAdcfAKafh+sbY0lSm2
YH6G6v9x10tqIJVelfzckqeqSZCTdiGe52PRAG6fQ5fc59zZSWmpY818dtgoNbiMEGlhnRDhEwQk
afbUXMQsbcANotyt8tPQsBz39+0fQhZu+OTE155Bi9/UGr0mBRULPHTiQGmEgYlsspwp8A3/6mNK
kxRfe9uJQrmMyz2PchTPcvKsO0qVA/KFScJzLRtrFXpDe3xF7isyBvVismwruqIeeOnepqwi21/k
/6sP8XEcI24lAjOQLrmnyP9epWLC2/8CfzO+rakYXPKbjQ+mRN6YvRaEfJJhmttw8w+P5P037s52
gNhiFhZaG1IOZ7ZRRXpomPFzaxvR5ZGYyGhGMCir4dts+N9KOxAUsZ9XIe61ePUFqn/jmtnxkqAj
LXTq5opCQmVm5ck1vYXGsdbKmUl8n76sPmskCirgqMPWA6zxokZ/vTJDZfNUB+N7+/ulDD9AYFIV
gKqCptqwNnTtqvbPyq8H0fzXbAOgZzkO7HtMQw8ZgOaCu7PvW4NeQ8YIsD4kbGwSxVK3qEcN8cob
7Qs/uNI6fTHyqQJkDfeLEf0SoVKEpJX2A4I3uqZTyyAIE3rAfWt9IR22sncwWYv4sNZRBBwVTaVS
xFF+Qgcgd5fYJKNvUdnXtzfvrKP1jrXs896JwQUYVL6SQVNZukthovBDCD5FWK+n43qUg8ETqKsA
yg2AzD1opfAipekJcMIy7liryklesJnoQ0mVmVR49OkVWagqYs+tH52SLk9GlCb1FTuyqK6sPnZy
3sWfQA0BIr4eWWxrEyOmxuglwhIB/40vLG4x+jU82HfYW5AeUPLEh0avNrfwLCt/v8oXgNIzq+Dq
LMAjKMIPr+cxjwuLQJVoGvE++qd2UtxTiEqnfZ3QnXpBEQBR9DpSev52RzLs8bZhH8QcZwu6W/su
o0sdCXg0KlYoRJqg9AZh6OVdXEeLmjTkw9BPYyszNed145vqYEwrDChyrUAh5qZ5jbQhURPRk9hY
IO0z8fR4hs2cn+27sHUzwVdIcetG5NAjrLfqzx5RLD5rjR2Y5sXfEhmmrcg8WkHp8RGOeIOTtIWj
C7fD6EwRSw8hBtFtGF9dF4rKPCbeu6emXqkXqnQ3uVYAk7dJ6w3OsrNTAlcMieeM8ZrshjoWEpfG
CkCY0V8fuAj2iStOOb1n7GWR+2m4w+Cw+cH2895DJztn9/4F8SSKIDb9LFHfxZ6g2ybtOE1JniWr
SgSlmp5mT/tRB8IYlTFp+wuYGq+YDb7hJxd4UosxvtwkRZhRuilHFPYS5godpjl1DtqVJ3/z8W9Z
F4U6+edJuQre4UyX7z7lnsQBX/CET6Kow1U40/Vaz7ZwnmSfP1A0MPsXjKgrSuqXvD879HQQSTXc
urpIaEcPYcuz11FZvFfm+yfNngayy082i5nzQ1ONNM7YZEyMA7EzqkbV+4h0M2oMPg+nx6qPKEWq
5Kv3rLywKAv/mQx3JiC39K1bFp5USRlezqshphlTray4FvV8acL6CdC+d1YaTd9lKgiJ6GEFkP77
AePvDAJITrLU48FVW6sz3Pv4gmBIUxWBrgSng32yMorszYvFHV+ZpLcJ5ivME4o+VFW7g9ovUwE8
RqKc1Ogm3eb62ymw/LMR4f1XMiUjQpikw4Qnnn+nmw4k1EOamhr+9bH5+u4XYpys+G8nZS718c4y
tz+qIuA1U2XW4kqpQEk3liFIiEoz6oxfbKAQJqDayUXR8Z6WEc6vnfrEkQ0VpXNIYIYfrBDSeF9w
rN9/6NxEzpFT8F66BprKslNPtaFQDbEZxdjDz+AeDi5RwUlHjST9288/lRd5PkXvFelj/mAH9FYJ
TJN3yvQH5O1LKCiGg5gh35Izc209ko8rwfmXpj8cErAOZzv9w7MnbyUSjQ6DOFLgLq8FmU1zmCb4
gcnyNk4bT/DSydIK+9uVoHmxQs8dZBaiaOqWU3pW3Gc3d6nFLV3Cf67a+MtHa8abP1FTksyJQxTc
YZFz8nlHNdr0bd1GgeMl+O2OUohHjVV/v7v3nKWvn26Jj2jbaUoyc2jyNUl3S7uf4PRYtNTFVqQX
OqSXWUSNxHjxMtWSw8urz0wG1WxJBRYFMUKwGvC97DpDWbXELHZVfrMcVXkiencUch0wGEz9yqq+
Nl4q0I63ZDpG3ZktBTRagFIEfvJfypQNKsinKDS1OGeg5UmK0nS9V9MQkpFYstd5ETELRhJCb0aE
28p90CzlaVAWObZruqz9WP29M8b3oZATplWNMJ7HTLBUwJEcaEfI5xxwwL8C6KYR7bKa0t+WQABX
ZpSVX4dM/WgoykoCeXUFgtaINiWsLGRdtBAyWeGIvd/8LSk/BR7xgp1ibWk+J83dGP+HHbOnJPLY
UwfZ6J7aT5icB/G7Yc8C9DZ88PiSjUGwWXSvQjCRfxTaZdxFhcJ6fcPDW+85v5PWs9XxRui1WISQ
6YgdcejIZZYIFXGg5b3l4fNxVkm79J0ciw5+VtontJGDqCpHgkdgqcovoB7JYScbnmo61gXGIx0F
2ZxMbyaVK0Dyc0q0bP8Q6djTdFpqAXLC2nlCGJ0w4JH8DUV8Skf0Ctpzvv8H2zfcMPvH6fHE+O+V
aOUWradbxjgXkc7XhRHiHq1H9ohvCwxTvnsPwUEe5CZz6G/kmayEUQnTH1VwYxM14MTyHMW2+pd0
/aI3KSyPiADA/rcUpe8OLBek1BzcF7qVc+hE4AHbRwz736nzqIccw91Lwor3OenKtCi4EIj81lms
V3JjoW0oZnmgxW22U0Tk17Q07Dp2eHJgQqiNxz+m6O0Qaf35qZ2nfrrfBPgFAQNVca+F8Xc/yHJ4
VQCY6wUkaEF/9HQZU5FV1giAKN+oBmVhoBO7HBnimtwXS2EwyDchbh6gzWgnAe1eVu9l6J8ltpUx
P9HGWERZNF+Z7SU0vVwJ/CRfa0ofM4bDEIahoTZNPwlXVbCKjUiiC04iaVPBPdIgssCeR99WRmUu
elr26TVbmVlAS849a49EXoOorhC6OOVK3Uczp6EDcrfC2v4CfDyntn8/x30hPo7RU/J/TTHpO9/U
s+wuNOWxDp8yuixQfgu991Vl9C8/mO03ZFVY8daFI7MDDAcl4D2Vok1X6D1xN/DFZKrwLQ/DqpmS
fZ9OEDC0JkbRF9Ucfl6x6RJTKVS44Z7xwH1DMFeQiWVZOyThCnu2HSLux7GVpKj87QBMgwV/rl/9
HqZat6Yt/IWCO6iCxGU/nEx9tY05k47MIntf8reZ9c+SAj98DBW93tPc81cE0reh7BNq0lYFtSy6
Fsit4A9A8kEwtKD3w1kBBjSRqB5Pkgxj2PSuQ6Cpv0Zsnl/XtWReHPghOpzYx6R2p7sgPLSf39Pu
hAxr+1brPy98+6aFwZgxp3LQfD6K5YrWqgIbiXEK/HckdkL0wzNy4j6hsJoykjnbxqyDIKdZU/yj
AxwujPfMU9vnKfouQQEefp7dAtaYsN84SfdxhyIuGvImRWjCrpNAf45R+5pv6Gy8oEWXwYbXBxnO
xipPQPSJ4KDSGHQhwSH8AxT7K3ZoJCPv2YUMvfOhkOEpPxKg9q0Id92Xky2S936yCoCzA0xJsjTZ
paHWj613N36YYdbWj+LYcv2gETVZ3ZitEFRkeYq1lMVh5bN1m56wTLhF/WckOku+SAiNzkHEiL1y
5JKgJezcDYFvawmzA2na004YDymCgbWQlA8NZKStII7Jh2K1QBTm2+Xo9LtHxv3OW7PwqdUlj2EB
J/BUc0C6cv1Zakt+F0vjwFtAUse9gT0Idu5gjzVoRYxHkhVPqX5O+xDHJXZT8CDzBg0OjxNPM988
5+rxNC8IBEuVHb9Jw/NN8Vo7aivdvdIta+p4blepf//zFKPnZOgwIvhfa7zgRDeH8XSyx8q8A53L
f/xibmUxvd8gIkrkU1Aitd+Xwx8N6/kQ8sbhnNe9XZxTKO/+vYGzIRcvnI//wGLXvORxXYjQHeLK
vxNCVDTPRnE6Kft/XeCCYdLbCIbpdkjSemTaGl3h1sMRxd82gTkh/c3UB63w1ZiPK0mItqZaRloW
AZ/zYbnwBCrqX8RSdZV6QK+Ai5nRAuVlzNvdSBAAMZuSSn6cJLPC0kHVxm/MsfDiKBAcTL9RzVRJ
dbY9ecw1IacrfTI7Kr3sx/QQOYa3+AhoLgcrNbK2e/0IYoLFO6SdM8GGm1NDQOq5R0g/QOIfvPtJ
JY0yli8tp4iLv66rmOnJE/qDPEvkw32n4UHE1GSgXTm+Z8O9HJHd1vemqlEoGS0verYPFqDGKtkc
E0CLwJJsGbS6vJ4xWLF7yy7G5Dednw4FH4Wv3U2SBmW5Wvc7lzS8yaGSfIoXx4NUO/Od1TqexDZk
w6JidbAV1bkSbrE6TAsqlNDXJZvUaixhWYx5IWwJUgMQVf46/kIsLNhoijuVCmfy+WqE6Ke6BIJ/
oqjXBEdUQoMdSXZpj65oSnbNjtbRflcI5XzLh4lVs/fyQX7hny8NMaHsaUJpVhle7FOxdzZXYhzo
IVrbERLdJ2q3wyXcdoTbY52H6b8UAB9IIpQr9MXEPoW/heZFrYZLgKx+0QlxZKy0kY2QsXuNwKZ6
sMG686wELQOrxNgXj0LS+z88+9lJpev78YdumBKenQ31+JLDZ7+wyHsSi0l+4jY0A5iN0fEa4pwZ
QsdahoL1B8PZs1vMLvH3xIjIMsS6zIlHmShP5pdq0aDKlD558YZ6V9UQhQ/sODrCTXSu4ANq522E
vFKTLsl1AcscnNXxKka1FkFGtsz3Pb3vKfqFbV9x7NtoYKxSVM1FzcBwX0XzB70rb3fKON+51OOh
jKU+gtsVKufgmPs+bhICl+bujiuA8PAwdhO2qHEKiqe7r4wVefZfgSE0c2NdOzVPzwo5PssYad6p
YdBIr5DKhWYt2s7KdZHww8x93pVqWh5HgiD5+0Zl/IE1U4JpGZu0u1jKjRxv0k3eWyqx9uR6p43c
DzmxEUaePTQOeisQFDiyhpwWHvnj5JdeHcCHGk8w4bQixPiAbL6FCL8SS5k1ejExXt71QgXRHHTj
+5Uhtq5ratVA8BSxaF9rVMTcQ+tvh8RtuHLg9MlK0Nm6GtYqNW66c5cTEuknA54Lrkh5KQgLrLe8
KfXtOLXO/urlOto7QtddV/vzyNdCa52+26zCwLWmAUKTkfCO88BVrUIre6ToDk8DCNLYkL4ygUEG
QMHCYDshjc2X9J7Cw8gnEtdAhY2u4BTTObLKslJNL1e+AB7EOhdO2uiwZz/0m0pAbLOA8mIbmwyR
Rkvj03ZNp98GOMkHUjFEuCCHrjb2tpKg7uPiqSQuGmvhGmiBXSXo+gBBOnPKDuFEDVGwnK8yzlH5
nBEwODq/gcwTgAoo4K8S78sORaBOaKi9b1hqx2T6N0TQr7DI0RqWRu83C1rgTYDiY/GBaiD4NAmh
s+eK9TtW/Vuby3j2+W9UAxRVmPKPadxYzJZqi3jHNMnkHz5WHfrU9HO0H+IuKYXe598AB8YMzWl8
AOm1TLqeKLzciB8VZomY136iUUcNTuJxRgjVUwPYdWI47h46exSwe2UQQh0rN07KuenHeBmAk1Eg
i0eYyd85Ztlf3GJIbm+hWopxAX4NbAWs2lCUjurydm6Mryn/jR/DG4iIpE3pxSHT7jYy/Bsx5/nh
qQYVfus+CtdlgeneV/bHafmSbo9KWNfzxMlZ08G/PsUnIwgxuv7baLgpUdAU4MRHvQp9+4Vx0Oa7
ejyLXfclyAOuikjopQXdmPdZ8g2pWyzAmb/7t4XZDE6/TDUMmwAGk0XlMfW5Cn4oc47rTr56sO0j
7mBOIMFHuweIFVAUYfczCnUybLktzWspIvIG7sFuqHWTCtX/znZFjvn1NBgsyExw5JrtBDh2wHuB
Tq3A6mYrmCpiEZlTkTh5Iz6vO5oYShakpDpMbg7PVdJkp1NdJ91xOQrbfYu3OhgxyZWNnHHSDRT+
40C5+jYf2V2I5AXT82Dh0jVheoV6e2hlnoak2LeeztCn62/F4jfkP6Fx9XuH0kVIVUolMuo4U5OI
vVEXmDbZoGWTgJIA8/sU4a6Jq1me+rsYYkj2PvxRGhINsAhpSX0i3e5BegMbkm+yzWewHUWwktHV
1nJOokrRvxer9OGGiDyfW3tGb0uwSUDit3Xq0d8+4g9XNDaM1voJyf8Rk/RB7Muuu/KtpqNEUhzo
hk74SrCUavL0/ZNCEkA6HeEUZrwqE+FiEJYACK6DypqyIA9wWKMkc8PjN3D6EAoC4+KRf1yep1Ha
2oB659vMqEvuOnxSEIB/t11aMrGgJ9zeAx+L+9orkGPEcriy3kJAKbIJANo++fQpD2bIqpEwcRqX
cjZfu+do8ltd4IkhrRTofkrHxE4ONay+wtwFP6SfbxNaB6v+/kWTwwndZv96SCWs/7filW4zuzkt
SR8QZM102lCwk26h+LM6F/eUExo0Krk9iDHt8Mx9q63Z+GRUrc0GQBBpmIR02VJLlK7fkiO1bk1O
9pTPuG3GN08XQ8V9WvKlrPWvFQxb4uQVXcvQvDrEK9o6rPGKLhvPwKyS38VTw4sboKfI3Cf/JurV
HyRwUO96BFQgRKy6Fi0mK/xv9tXYKdllMUkNtxfCZH0vkoGCY0e7eCjXCsmDXcHX/VTxUegITPSZ
ikNaJk/h8FUr5Ijyd95W/QD2Oj1a6/pIEPI0dfq6pyRaRQ3eUJ0LZk33sKG2kMrdduhQm/zORR9c
pJGsTdliE5+cXlMMQHOrezlyYKgQGXrQNcqzmh7WFMjdLExi46AMAF7GIn9oTGpBbpZMWGkzH312
ZLFRlF2QrzaVEBp/fKGIAG9OoruUgYJzQ86EFCZGhvS8WZs8VhNQepJk6r/IbFxMsRQTQzO/aGXx
RoWRW9cnznl5JpdDLYQIc/DHD9ek/Hhs9om4UhxciBVSjPV4zekT/5Llkb6Vbv0ldZm1hiY5xSfx
zUtGEShJ2T0QKTgJ95LmKE0IK3smXlOJNUYo1o1+WovKN5jciGIBIy8qnWo3k3DcfTTUZKmQJ3Zp
O9z+LhK2Ij1o9rnIU27+CSBlxzqNaCLL/IoiHxf+K613Or1e6w1GMOB+7wEMlSTQp3aSHusVGYsp
Xa105qJ8twk4gW/uElrNMw8WyMRK8DOjS/VHaYPGjDfAicSoOCdJ/hbfjrQ9SZW3g2udo2/OR1Bn
0FO8s6w9CHhjkpPg3bB97LBetKdcP3fDaXs8h+fgA0qn9b2TlOjt+1RN+8K2cnEwHLtm/k84xBVy
QGZl5MCLvHPAoKYMwy/RAF6IYiSuB3UXzeN9WG0TykHL11FqUOG6Y/Mq2gTx3Ksc1ei8eYuUUVFj
OCuQcrN0S79FCOUgfbnC4UJvz/UXx5qg4vFHU3djc49V1rY04Jwx5yZBVoWG9c7qTTdgAGBm82YO
Kr1gqvChYUkOjJbTjU83l9QPs6fO3rO0LiVcrq1+qyALL6eCXj7mPlDawuMEZFrDFdNHC4oVIRi/
xYKNRLNtne/On1YQLf/erAaLguecEO6NinoMBa4tWJ/1ZNL6/VJIfk3ELAnX1dwk16iUHAYpx9zr
u2ND6WDWHE/e0S3lpwcAqg35ceJEekqNor5wl3a2WcT4g6iAbimowdnc7DINv665nOnDDUfkwvMD
Ab+fygSmcLGIw9r0G9bc06Di18uJjuYGDnENPAg8r90uOv8jdsB9Nvv0C6MD+EhF81CG4AWg1Qjp
FAMDazrhqnhApujS6AZ0i8ohfreYr6npIi42pXl4/IQxtq7EPP8WJRvuZgSqXq/02mDnu2BVBemj
dPA5gogf6esykKP9/wc7C+i+qV9X2+DpUfeSEVyOnBG9J/oBT0EFGqtswlH+Fk+KY9ePpyPlop6A
Olsl0TRk+CRvWXiGOE8muNvHsw+IRsfoZJzS9qPnMBakLjas7wxuZusURwlyFYJp10X6YAYkBUIP
87gsCW3mrB/zrkAyuzen+lFsRQYTvhhrXKqkOfkNhdDCIURyDIIdmAs/xgSpb55el7pqjFB9VeS4
Z3DJaUsTF7ZBUXFy88dJF/dbg/zOnrcvITJLkCOBB1ZAqAHyMC+pn+xyIJSv8rURl3aVRpV3LG/1
HDTNb+oeaN1BAc4CYxregGwwFItP6QCFSzAmNkbbFHVkp2EsVTVqu5D++bly2htQblwmds5XJ67L
veSCNhDrKnDinFecNlaQjFHWmj3yhSZZ5h56JU8OOYV/C6q/V5PMvV65dxRht+okMhd1hkHZfzUs
7nk54emMXtX8LvJMD44/K1/KHjixl6LHF4aYnF2s1FfdisD9eHSnpfEnpNqmQ0ZX5nQRGzMX2cqt
aIPcazCjrhSwTfaYF44rU25KpYoYbxm7N/5VV2+ZsqAb9F6hzlC1YYU3Y0VSEAP6wSX6O35spClA
rt+VO2D3xeOzkC/2xOLyE9bNOLZt3z5ncCeoAY+uzB7YRsaSixIVXXuXL06s70FBu0lVb+PznPGD
UZ4UzsSEuxFeuL2ZA4PlN+9qoeFpFdNwGG2V9I+V4FVJnqMGrzFPlOmy8zDfJjefAff27D/4O56Y
NUW+VkYkKxmOD9D9Y42vcHpOcxdXEn3PHexkJCGo3hIYqzh7oasiRUrjAArcVmhxtR22aXYLY16w
E1hSJSI+UkR7sfPytU/HIofzI8NTH5pmBGvHXUMwPtGokxlz8SFjZabuf2oz2Yh7KlxYB5s+VwAT
QjGGlOnUibbsd68pyugTMexH8FnCxgvH1Lb5aR0pZjk8tF4G7yJ8MS8fTmxIyWrCr0x1ltbtsoQZ
4xVs37DGS8U2wKbiTrUpllkIo8hPgXfR13SnNDBhxij+obF+IEga+dmvVUwTxb1j7GhMaDaniWH/
6NwY3gR4R4YubOC4ewaJcgx/XtjphZj80B8VStbyuKxuZichymMWNxQ3h/GtrLDsMWBXXbKV2e+J
DRasglhIisiVOa/zP7CuJrSW+qu9oqlb8k+BkIz12OvLD1DB6BhCF7f/tWP1D90lDe44HL+XaWrv
og8z4QTOe630sbDI4XJu+alPYpD3F+jOuwdpcbIw+VQnwP/8XlRum0aa5x3qjbNiHX5+U4qRlj57
l+01xf3iqVpPVYk5SszuxJKvFykhcD3hOHfSFEWVYRxpwrdUtRBn+kygQwYt3Sqc8psVPy3sWSLq
OLoFS/BdZhOuRJQNEGV+5WlRBkPPtSZ7ypnc7QrgfrwQFih9HcHJt6MnxwsKXY/WoZ1veFumpmYi
sjw/obuuB7mvZulJdmpKxWlUqEfvb/f4VjaZiqJjzuPUUyD7p9hHbC/n0bpHXrj5w4gLN7+enK47
Mee42eA/YZg3v0Jga7CLv2DM46JIkHo7FR7bL++VCYFY2GRXmYqA30dw93ilenjEVpF6lGMTa/4I
lX7SmNovTITlkQEnMDMk0uBBJWbfChZpEB41g3jeNEMeYbxA5f6++WaHHlL7vfJQ2neYhIIkR3YI
nj3LlAFwUX+AZyE+cX49xPNtkx5i8IAE8QW/lqFEq4z5AFPahx1V0NqZy1gH+4J66c/UcgiML/t7
G6rQW7FxRWjSeZi42RsoZWsbKuNC8GmpQRLSb1vFCKiLaGW5ye8PafmwP8PzaGNEdRawXRAZDnfU
JVV7yfuxVuaI6ttjBbxTbBWvwpguXaa4SCEBJ8OEYvhLKYBROyoO9l2VKa14lokqtvC5gEJ4k+em
xNKVjZstj8G6Iv22qmiodB8rtC8gbUMhd6GSNHTNVFlH/G92K1W71ZX1i+ROgjpdwqr61coQh0cj
2wZaWkA6VCjcu/dHsdJEOZ3oO7YrH7pAJpZ0FGE1kFPXuUGt2pRFYoympMgC6kcdoJYT+rg/QKjk
1aOs/YvNeuo+Y8fszVOhOje3ihIBvxy7uGdfP/L0EGVOezP+TQ7iBho6JXE4q7RgrF7v4Um8B+Z4
PR9dzi5lLOm5Yd9QZzT3EewE8JzeLmGyuC/YhlIBlmaZlvQCriQkL1nz/w5S2lqztR5fhTEJQPpK
OY+fHJTdUn8h2lhLCbE/Uced8GmZ2CANcba+xro8DSSBVamrn5tRKd7ePRtJYr87prwaW8G9By8X
GJNYj22cPwX+XION6WQZIJy9KB65SbZLVQp677ghrtwvjiZULsUc+439yXTydhHCE8504DTIU2fD
grQcEYYLRzgfQFVp3qcXjT7VSC1Is94q+PYx4EA96i7vyzGtH3z+AztZhSb+kI6BLVm4bBVrtSg7
Q3fSIFlYcoW1r9x72VdMjIUnT6Rx5tWa0RjagqkyXWMZnRpgdJE9NrRbdQXNctCyn+aq9rCeb6Rp
mslce6FT748SRSevCyrLdpWTsOeBH56FbMDYyr2WYqHT3JHqGF2Q0468c5R2Q2sr5TjbYkosv+fj
T49SuD1lMbVL/cVjwpmwGWrz+0QkXZs/ekjycgl8/g22sKaJ27AZMtOjsH430aOqsglcKbQcA14e
FidtyzjdjanE0Ch47KICEtxK9M8sVe4G1qyDlCuvqvbJnAdyM5J4xaLZaM8DAh/l464j6wRwWR8Z
ObYOFv/7+B6fZQoZgnL4y6oJXf1YZVDjHVhPH6B3hSEAj8xNw/zqEzJ3LGhIDea23SY6xXd8KzZT
pf76MoaEJs5jSd0KeiVscUtBMUigcxVyskN/09ZrE9nrojt4do/cRaiDXw8Avz2PoNQka3kUfUc3
PWvwSFzHyGYiK2XBVHjY9CdJm9D/xIhz/0lwedofTVT04XpBDIqgIHCBtmVsKk6UfaOEP33Q6zTC
gy4RZJ/Zv8ezUjAKYohBM4Q3q4WoDjSOcuBHT2OQAyrTX8lo3JmQKKMUEz6XOXh6+LufoSt3vfIz
ZeWA1ZqOQHA2BH3XRMAEeyNbFDSsQpNulD+4aeFw6ZS07rDK6HDplhenTuzRp3A2JW7zzgKm/Nbd
OJ6IlnS/h4+wqQuNDIYD0nByv+7sOdSZaMT99GFKK73p4XPyPNrvYc5ArTXbnKo//722vLuRyFga
/lghyFEU2ovEExoM5K7xXpHtea9ckcWiq8yoMNjovd10P9CF54MQekaiFAAQUNnSBXD1ffu6U5lZ
TADDTXJ0ee76hJDNTiFSv6agFrn7l6IxhmAdmQp9Uzrzz1UbhDdFSGoBIuAAfXsUge0hreo3sIBl
E7UKa52y9HVHOlDNkayS/85nro9CxtIUn6Rpldv6sSOMxTaHCr0dvMW7ZmB5k/1xkJO2RmgZiXTL
cW24tXTNIsDbDzA66kPfnR80PY3g+XgyB5113+TAbtVxFsmq76wnkr4Qg0K6fLVXinkK40DbTbhw
pXcS5+DCsJXc6DBNuW1KBln0ikMEM15K8UV6I9JzlKEWxrD35wC6ON5v9BAbUvpdGfwdtVD89G3J
gwrNyfplM9shwNLYxkx/2bIPjd5z62aLqt1s9Qa/p6KK2aTr6yOYScknlbQt1WyFUCiVV248GMsI
uclFTNe3CBb1R/xK/N7Ynud7HKHBk9/JzrvQpK/8tKDaRxVeixeLu+0HPMNXuLvApWULkOOF78Bh
ui08Z+u0/GYM2QeBCXbt8yavtf4aj41FXbHKl0VKqjDWkZyGwzRndOoswMQGAgoSd68qo62pvXrA
kreXDmXLwsVVC4iD2KEzCCWMBFjhtlKU2pLlkupv73dI6wLRCZAt2TG7E3SP53XIdMZpgpGIJkC7
AOqKoKbg/8FT/xekJLUbqceloIyFYv4OnyEbPzwGFqOJYIdKM9wsFa0HCJkU9imAsx/ahA1lEIsj
bti0XIqAP9gfOVn2onlWeDV3hiX6XGE4BR8qU54GZ+gvdGS74JIRXXkeMWroB0Z6gSvc4QNtzyad
nUJTeS1PjAlJ5EspeF6fXss3Lq047DMkfLDmZ4lbb3I2omqmd080YFtOQzwnj749MJqxqvQtpSq2
+8BmxgPbbR6ILX7BUph1TCOU73TT/+aTpLNsdFDiwrGuF6k5eB9WVE7sKCjXXVb9iIQwxM+RvSku
PNZjrJGqon0QEO0Ke5mOFNffvJ2Dd/GOVkAenmMFTrPs29Rsj+yh7J6Voo8AsWKs7bmLcn/SxqIs
TznsvQRg8/TNTlyNgn8fYQfBLU+u8yA/6enSeThi45ZfgW2a91yC8Aaf1t/ybvW3rhiuJ7zLtUoo
kF2mnsKXzyFmziUJShmlq/YwFpDhGkp6n9F65exfsnb3CfIBNGrTRMXerNXHyc/oDJXpXdlCvHsX
ZdIqPGXPciMS9W4DfyiqMkIzyZlHvMUrGgyt64v0hCptpL03iwyCrcnnA+8CIm7bASCLiGY12jkf
b1j3PM2jEoNkK6bq7L7I076STCh6D7NNXpFbZUDHr2RbHRlkaEOMOrne/W1A+Lxea5auDItyZwkY
iFfVwZKpc8rN+8TVaEVHZiTtm2ERa7uTgAlJqBANqDiQjOkp9HgNxeeI/jpPy6T6UbkWljNHxg2W
DpQNtteUiEIn4dgMeDjn6Mzb5Cd7rgK/xBSbqdtzS/nWcglLLVpfZbyq50l9hnqgJesLvcDgA4k7
X1vwwe+WordYc04C2knIf4sFZHIjBRQjIOSkVzhENnVZSDsDsqmHBAtpYTViLwMN11M5WJVfJkBb
Jsq8TTJNwZsF1Ny6u2OdwIF0VBxkCCGVK1Iznr65LmhVV0Xm0jKnxAP/fQ4k5NqPOYkdMPTB6QDO
LqMWk0sKN3rn8F9rB8V8IGVMMLhN3v3dsinsolC29m5XxsfXnG42VciiztY/q4AT8rScL3CIjQaj
pR3kxg61Io1O0LgU/xZyP2lygOuyo8NPnO9X91nEIWHqp8TN2fpXn0IqKFmv4qdLfGcCQoT+G94w
F1klp2H/pLdpaPKFT60At+W3XgdgAj5GwchiMlNTRMJRFt5AMmHPs6xzZKfyKzHQgHP9+BfJ7057
j764wD2GCC8Ebtg9DdaQJPzmk+3X6kPTc1Qa4zkWkbhetNjbzrLfpf41DHajQLeGP/z6xU6Vsq1w
yFGQlp5LJvTRu+Eho55RBsKXATw0+PDqkQ3wkcZJisjgMXZUmYaMsPqNlzoSDPPyXf1V1RJdD0FI
WODO/1rvn+aVKtN2EDkbbH6w1TnTDFCbXsXVyT0IG88QyEySqNn6S6JLowgBtkW93EnP+2IjHwZP
7DatQ4Rx9C3at89LfEjuBlfumtJn8DDSxRUcpK+0UsktasAbCwdavSLMGcUWzjWkoEQVrwjbwG2V
dokhpScxcjEe0eu0d7D1jFGVLRdCAfiAJmODIa5HkHrRwQ1ziZPxNlJChCYbeVKmOUmjA2rmP2GV
ukRf1It9iDtHACfYQBhCaiknpSlg5MWGYTCO4uE4KFy+5SH7N/4weyen1BaXCCZN89OBz4JL3yXx
cxJv/jqPbWtR3LxxO/6cNL7wtvyoSSoaRQBk25aaxOQGajaPhaT1Dwl9PdqPX9UCI9yscfPMVE7b
yK48kwTdG+Xmbsi3HBfd6gBclAxzsjfSRIs8OvI9BkqYvEE93ar7IPdYrXqUxpotdbv34T86Ez1M
l5F5UtEXD/7TWRwFcgaslS5yMcuXn7SQtea2YP1IeV44QkrWWCmzXXuxuvXESMzq3rJIs7u2siBs
hqUlu8nDir2MqByvYA0YUMhfZCPxHXPfNqVP7qvZOSqD/z6idZk9sAzkUqAXnE8FxWgQNBNgzT7M
GGV/JxWcLfiP1huQKli55M+sHA8HzgvD7qaLlnFmA7VpMiJmgQ3uGWzCd9bsv/Uj+SMZEkGpAOxx
TfZUk5AL9srw4pAG/C56uTfg0sRgq2CMe84eI0ooNWV1HTah6SXiYeEdB4ueQbc+qcwxNySxrrh1
RA3O2Cn0QWEge0F78YUVR5tJ6MozN2V/7JvyTJbJXkkcv7L6SsoB6B1/ctTSicNAHnFGgqY3vKeS
AOD5Luzz3iMRFcv6p+bgbQT5vy4TrMtu3in1tTxCwsnDu1lS4uscqOUW0Y9K8i+r+c+/vEy2xNfD
lu+oMq5KAe1fk8LsT5H8snBdRsjK9nICT0RoJVDXI7yljwoqmIE+q3fXUuZGdFJ6Wyc9bdoeBOvg
8Wp6A1MQP1VytM+T7vVV7Gqx3GPEnbWisEB4lYA7xFgF6mywyCm57Q40Ymv+Yy6iT9UczKAjjT6C
gPa5NVVV1EVDLYkRA16s/0AUBIhA8kj7XLj+wnoENtYuno+pAeFM2Bap/TyE4eqLyGviQlMFxv3c
jigrEb3XE6oP3lFom5QkEreD4v1SogqB/Bd9hw0fLMWAOdoIj2ESFW4iO5GCBTV9St7BE97oe3+J
uP3nsntXq2RghUWmhSUMr/YGZs0RAwgJOmHBIi8wWLiJ0o41oZkmCsjy/x2OOpgtjCuKlUPxhBKT
GyFXN1+NGcAWEltnfD48+DgB7H3+MaJh/7n4UfR/RMSnlnDjfwEHUDEcw5XeadzEd9UFaRP27FKc
WZIHLz2J6HgqPVGoLc3snJ5jhnChGU8xiQmNgo0QSkrUFiQqqQz+fNBSV3aKW9uBvywkcP+FHQCQ
SNKd+f94xY4eiYJaiHJBXyGVt9FcJn4wcvhd94pN88F6tZOskbvDlVwJ3lrNzJolw0mpOPUnsN2O
a67sUmyAT7/xgwPT5nzyZA7j2DQd49rUxQKEY5Frev7I01cEy4Zl8czRIS4iyHVO/+tHIh5oJgoI
/bCKXuL8Zc04Usb9rShXwzBuCP3rY7duswiHAs4UvsCBC+fZoQRK50DU0eKJRXqbHhqUgnvDA2z/
vNnXxtROkhpT65Yf/Tj10RNTAIJkxGrF7kbHGVqySa2rLMNrzVU1hHtGa2hIaaGBidY0dYEbr4aw
kDwJ14X//b1PaXedSjMWCzgLck1p1202XrJNR5Egx/Ap+IChNvzLG3tR9AXfcfbA6tykuBmcoLom
GHE0nNGAlEIhGG7iEYhAXAvRQeUXZbBl6yY2Zg0L9B4tog22XIfkF6I5xci0yS23pCVo0dIKi0+b
iVTTqA9VeCqqfdjPad3ibVyCC2jdEvheJbjTo6vf40WZlns1T2q/zzjErNws/Z/QXKlgTZeLA4o+
WDVvc0S2GcPcYf5ntMtWW6aksKiFF6jHYjWlwRZKhvaWQwusi4jRsqVvdjuiEXxsfyNni5YEmI/6
gV7l99Ylp//VGB9PoxgBX6I7uJBpOU7/VD7pJcoC0bK8AQjHMSw3gsTWkboo98LEAc1CefY+2o/2
++50QM1nLyJjOGqBNlEvfdcOd3Dk5xNVPxwRDP1bckuT4v947Mo1vO2fnvDp/MjaNeTWg5TwmcOP
3K0k9fV5D1/wi3NOXFZ3eR/eALWTGpvhvyjwdLt+xuil6cwgoFDIwh7G0Z67we2Ssx33dKd/2h/h
1mBC+hH/b75DCl5s/+km8TYv0s1SMT8ExbSrdi6566SjWvYMdSu6Gtw1Gw2PS0doPUKIP44yON99
a5hx3QS3Za5tGOsXVSAqGbrcaqzUOK9GIv9EtArq92f4H0wTbSywEnZjJ0jxTI0CYNsRZkCNNkuB
OZdbjfuZvR7BDvLvpy3HVW2BswR5/UtlCyCsHREJLADO/4p0EhUnICnovMB8YUUw0D5pUGlGR5rx
yhIc6BLo3kaP16kCCjZB7y6ywYcRYEfUF7Rt+zpW0yapCiVA5kBPZ9jVecIqp6KKA0wdUcMhXeAE
78dyiLa5LGO/OpsddVN9Yb50rKDsGWpDtuFnba/GjtS2/hA3ieZT2lqM9ESpGvet1J+EBEQ/sF8R
H51AUNuLA7qVjTf2PLWuanypfQZLOGbjAR38+0X1HnKbPy7l99W5O1AH0whNpCUkE7J1O9Y72pJS
BGhA4Bj91EcZZnDllIBAZY3t/kywiS4Vqj1/E0oONLUlQMImzZl/V9AzDGcZuRNxXwEhGLYtVffF
kDA8oaOhSu1WjT9gS3CBKbKMTD6YGXKh4Bviw9iS97Z4gve2q4VD2YafQNjF71WFKFbIOrrGzwIF
fmh5GYYOAvnbCB9kZ8n+Bg3braDpfKp7rfihZdarQ0mbzerJvMk1aoUJP0AxEuAO0VCMDgrvBL49
BN8syQxV1+je5wH45W6gVRWkZrnkEkr8LT8EMr0lY0TebpCap9oGBUt6uAC91bKRo9J1cFsFaSZA
ys2Q0ETnLt9kNss07JtQ5pE7t+WL9W0naTCLWiEtamp3quJRZ7nDLnX9Dv/vADKCEt5KOQum0U7m
RKsO+WKoLl2BRWQPZD0PJrU5E+P/2m2BWYh3xpltWAABZGaUfkoLJs/R1dQ/88h+PX6sWunAQ7Tw
n/OI9f7Ydy1InViHi7aaHc1djB9tRHnnoWJ9ufrc9lOxgqEhmlhxVJdVVSlmd2RDm4nAPOka9fj1
ImynQDzy+XPTXZguaCdx3a8rP+EBXhNJSDD+j20qOm/8NTfEilopm9Bf+nhPdcSaV14CQpx+JqXn
zQVolhh/1AZ6VOGKbrqlWg0OG4GMxQFvm043njqTdIH68bnmBPJbmRJ2mkOWHU0nmCG6FGJbktmt
a4QDoSW0rxrSMMXkX9L1yTxMNccDWcnEKyRzqDDkL17565t+T3jrY2VHeLj/ynFBlk7peepmZ5qH
piYus/y6UeYDyc1CHX+TT9SllFaH33Qvwh5Yaqeb3KTTl8qde4mLf139a7xtE3lAoLBmJHnRb7QO
NC/HG7fAxIM5zODjBwiZOrKdF9AEx8AGnelVBT6aBZoomutXnXP43aNh5UXSvNVbaB/OV+OKELUa
XYaFbYGReAZrQ4y5PTZqOPOT+kZDwDglZafbiQMgkYo9dHLB06bokutxXhyh4hqaulunyCjWflUf
cLsL3wG7g2/HXAH8CXsaqlDxKI2zWsJxpYKb3cx/LHscNLF7+VpoJ6ZMmUc+OpF/gCkKANK2kumT
sPD1cjR5pNO5qM1OWon8dGzWK55viev60ksSNW9BFLX9130urRU8qWH75mMFHhxVtIfXlt3zhWRq
7ePBI7f8VR8ltZ3Fs7qnqy/02ns91i/S9eToMcrmtZOHO9Xh9UKciLK6+dvrFHyVAVXvNsI8Sq0z
DHeAjnbqX572RLJ0YZgeP0k04fTWClzmuWgQJV9QR4gcTso8MIAScUide1in3keHTZqfJKNLvglz
9hlXwmoxNmCWz80RYs3hV6RKBKm88TZNbBM6RPfYulIKC4BUJ5OuGwoMEfw6LWpVQDaeGcSp7uQY
5xFDm9p4SqCYj65Zt9XV48mQsITqPs5QqIKlMK4WV6kqfonsHdewcP3gzFBf7h3ivbUGH9PZ2JvS
m6RGaC92LKLPIwTWgxDmiztDJXHjvXjm2bCSW2LTD5u2qLegPJ5barR6UyVDcDpDFLDJfHNNRMwn
boIlMbCJPDdpS146l721Vk6isUH+OiSDQRffo8Prnt1IPGhKaqoGS30NZlrjQaXnPVYo6pQcAW/d
rFc5p8j/o6NAkkKU00aoJul6iHLYpsanlhN5U79emfdmKwbWlRmYsjKwl8AgmyUsh0+7XSqhzfPR
/S8X11ushS4eFzaRcCvwoU2px/d4BotdYxx037qMudoacakteYO+xomuXQIbKvXNtBqOIT8WhYo4
1tYV2VcYH+PiWssNdo0rWhqJxeoM7WnGQyAny38T4viOk9NwEDUvrMrvcMvDeNk0R+NB2HKBBBuo
DK3i0oasyOF65eB3xcsS1ie0DUMbBFVFDosJz1Dfg4aIgDj0YPlQK8v0RTNIPnXf8raxeGCQ5YVp
7Z89EXOL3TXI7bpiMr4tNFife2oyikLOpd5nna7JWTtb+IT01nnz2e79AtPhDLmDGpCvSk74F6fu
uCDTg5X9vEXgHB3ph2KDrqz1yqrFMpL4UbE1xOqGAZCTP8hTxwSb/EBKahdfUsIJzZmFZ/Inc6fW
CyT25ETycD48xD1m/9AZwcWHYe/esvcZMLLAWY3SgLtioF8i8sl1YWOm0rjTp9/wGJpfqUra1cv6
Vv3zV0o7JosEZfwOxJewU00STQNqeOR8HUWhNfU8yc+TMwBDzBd+mXTglXNd0rjLEUV95ARyi/pP
JoK10KJRnTy60EP1o7Iy3fO/wc5XYUeJoucapz5l1LRvdf0BiUUGgmfsBjAg0N3ngd2o1NveqoMA
qE4QMXrvGqs/6697uFJBMxSks2B1mIg1NLyDli4sqwTSWpiQHkqEHgdJzX9vIZhaE//saaW673Au
QwtbSrh3IKgS8quKFtZqAJ0kInQXT4iYoVW+59DhUBF8es4CtzHJFzPaZ7CF+FtUQ6kKQNV4tP6x
nLrVrBVXwfUuohaqlidPKNUd6B/5UmT7x2v1TqEtjKMbYSFXX2CryUBeh7HxjgrcLRBh4hQz41kl
cdXMLHBr45+fZy/CToysjECSV8O0Ejq8tWSwjpOiLYNTiiD78H7DrdUmFZ4ieenOXGrNpyxlmB3B
sdalhCaKmmFQ+euLkxD1svnHEr/eFTlI2kC1AtG4fk+Kl0nW55o4xwJL53TPmcyxCyD0yj62CMLM
epXPlbohfDT5MPa9Y22LR6KpytKdwbXmxmyh7O3MkgOLzXlyREtkzBXdMW7XEqygAiugtH3U7SX4
GrbUNOJ3Q3TnDEFGdbcTIFdARqeIZSZDk2m+t5M2bx3jDASjAULbfKif7aPSqCU3/wLIwITw1ep8
BFVz3SZZdcwTQzjjPb++goFwIs00/HBZR6iKj0uP6I/Nu3OWk4QacjFfrk28ud3bEg905y+uiiGw
S0P5SKqUWWFD/jmPyb8mppONqmgyU5jrYMEjgCpBf1hrjiDJMrxtzjv4cBetPcCqpJh/SmTINp5m
d5j9nKoUMQyFyGelGt9116US1SIT1P6P/i0iO/QWTEdBKqE/+5eZPSyHYR3GhRqvWIcIQNc9J0tA
uLT2aX8n0WcEUQN1pG/Wax0OF/6krep77M0h/i6JfgoSzihGhxBI6b0ffx+4XXgbR7iIRisKplF5
urM9Cy++9716nuRKb5w2MQn5T1RMOMj2EyH0PLqv4JFMqdj5wchtJ5qB1nTHqmfQ4rIWdSdnXlp4
mCUfp19DCpdDOkvx1sNHBLku/JZoBdpYehjDGGB7IW2EfVpG7TVuiFR+eZWiSXDvxgUJMuGhB1EO
hBduxXSraY8ZLwU/bBhq3haR88BcH/HmUZU1RBhRxqyw1xXpK2Fgp8PFQxH+kE1FIy6/NOFtOURe
oKnGSofEtF+Rai6L/MFYiutNokdRJ0b3dJXVNo8eXKFQ5xoPhrtji+xg8b/xHhMX6nBwNIlyEjxp
J9JtGUMFxrEb05EgQQJuFIQRGrHwwRsGntHwXzN1jZfKpCOzCkoo15a5Vc2dqGsS3KmOG5kC99oQ
uV66MixPirfWvVjQhs1yBmzSjRDDvPJ9iAhyOs/OCXDkwJrF0rObinflFah+DSL4DAyYyRgfVn5j
BnaPyXXXmx+1ZsAo9RxGIMyZexl9AHE9wy7Qf7GZ2pJXvJtvK6ZIg2rWG0qhMoVEWRp0bhJyrAFR
wEBNLSSAdLif4C7cqloE1HtC8zFxMMGS30l4x/1/pF3OgFWu0qdbkz7UX5Uqga2BxNRQSG6KtCd9
Fhy8pGUc/TnWQDlnZjQT+afjV2gg6q9JadLNNvXj6Ow9Y5EX+elLqUYnoA7zyAboWqg6eKirm284
Hu5b89CgcV2oGQfyPL4TAg0h9JZSQOvvrYo8Y3qAXHbEEydUb9HKTrvVbyQbHsP1C5HH+AFKvzHP
Uyns3W4DoZ3urI/Fc5/B1bJoCm1FVP1eJRHHleEMEtau9Ynb34QIbalLRpY8Gm2HZFIfMuXlLQk2
yXeUTbCAYgDXoHjqzTtj8/jAZ7D1b/KobSX6rTFKYaCTPoqVmFXci2mXRCpWl3ThOUFkTM5UqRNP
ipGmGLustdlQoevRCBzX0i3ROp/lW+PqGJ7BaSnqsCl2cjOBeywZlHoK80cNbi6N9PzNber+iOyi
pLAcCQ9NcBpEamUHgAKK1/72It7NTksolJjSI0Zp4x0T3T4CNnQLtzjEGmw5Op7BRSv1QUlLdxkh
edd5ocSl/eOV9oyiWPtJkaB3t3WscoOqhU/SSSfvGoiB94vbJX/HBFrWsHXI3yua5G9jQe2rSkk4
3eyQxFQQYsjaPZyzAaXfYUszSJAK4RmCPts+8mFccc3wfqrPQS7oC2myL6U9yhuKtEGWEUs69XhF
7R0kq3L0LtGMxAyGnXyZW/kBSfCNilXVAI7v2SDpyKow/sumXg1GJhobrdWHM0Lpb73y3VZlb5Cm
q0aSlytg6Gov2aa8Wha260fpdl+EC4G6DSg/raCpfeWilMUhmi5+Z6BClOtFIWR/zirB8LkdWBRD
eTagWtbP6wadQl5/fdJoSil1lz13EdKKL3APIwPbziJ1rBHOCNpr7KYTjNzt9SUaUh1c9bxiOOSP
+XC0+cwiM3p0v+Abyj088FbSFfxRTAgvAesdqqmOJbL6clm0II6eTBsGV8jC4L5mM7XGA69QEvtd
9n/1A9igXE9Cakb3dMrGsmJ2Dc2rJXXuFSkxjHNLT/xvtFC0ZFOpy276Ovuh95leDcPoh6VWW9AE
GmH0MPZS+MclJLlaqcM32UEpZSs7Nz/NBt1B5TRgA8c6XLWMf20KAuADb/D4ZX/sC/Z5+q2r6hRt
tZQTXAeabExyiJnHgaW3LD0eqD44NXFicZGrLl4bbnoVHiF+HgcJzZePWUccJfta8eF4snrkpx0/
BzmW1+Ys2/uPybqZmXNfrfabTNyRcbecdftjtr3z3XcVlxySTOpfbQbFJgygyFb3lQ4gzwic76Vp
1LSlki1MVOOJCWB4B27CnLqILhRAG8SqYWd2AO+1E3FFBX38oobppZG3KVTaev8um15+m+9RWpYr
Hpr4vcBYcBqyiRdjYQ310pOAlGM6t1vFdsAEMP6GHjFrn1SvE/UcbIDCKjmVhduBz8hQuONM5NB8
ag9e9PLPCzKF89dzbgTdjOmEKaNIvk2rXUTHdWEWH06PbrTHYO8qsp4wPkP9rw68s3pY/+WIpNzU
tpqbx1c4SbeVR4LVITPnyB4bbsLyx3KhCD9PjDAZZ2+Le6FhXmCHByOsF/yCdsyHTRATKHwEBo48
h9WAWK/2kp+UCnWSMImBcsSi1t1RTRR8mUpYgcbLzAtcgVRkX8dR71rKnxwTDjc/maXM0NV6Ive4
KMdVbqrvPde6ClPKbqCDQrlYAx4K6XKopMDpa2YYQpR47Cg3NDtwCJo2RhG3icHN//Ib0O74b4Ev
L1eWowYNsMZoAwMyU/4RDT2bSVLlTDhMbEHhOF3BD9p+4FgwN86HXt5uz4SNJGWvxX8E/EpbfMr4
d2iREyRKZXx/YKM+gZld6imYX9mtg5AK0Y95eNtyaZMq75lsgYU46akw6CZNeDz1rpt3QkWMUDFt
jbmxBeb4EK/3m45slFOK4Mzw8EcO1LN72lmAxfbuopA7bN7kqteIczAQ7RdiTJ1bfCIztffIFIfr
n7fm8fxLd/qt8OZp6sU7D4jjdkPxwWT2S3Q3NJLnpLhd+unhHVvOM6x0+7aY6YA1gLKEuOKnTt3m
kPIO0meQydkaZRwdHwkbrd0phvrpwG4fTBCGIftGTKCizQCihDzpejWvjbdlfrg3Du/9aTRbF3Jx
7b6/QyNUksQAqW63f3up1qnSO8bfkyoMi+Ht6VsXo5tGSOekJPsGsu2GoIRKJZre6Z3IhJr/31UT
iejDHMilFVkz6xm5xyY5+iZhgqjrqOmysk+nw4dN2Q8CGhP/ICh8jcbWOWK+PRL+IjHrp7S41fmi
Yrm3UbTGY4IIkqIU75bn0uHXR9wmzcMSeARdQ53486hUQOoese+nFPIybTA5hE5XKZVGs9dKF40k
ynrzKCKOm8ww1doKvgoUbYv0BbnsiPQYnzOzpmdViWKlwMioCtkI+fpUhXyolf7KWt5xNRbnsEGa
Mz2SCS7ED2IHTttDMBq2NSxqjktFr/Bg+SvgfykKXIB6d+AHdXPHOMIEFh02jJIT87Wa0ZzUzDdN
20sqX5nw0KHc+57+0Lriq7TsvTRo+yNo9vEoeICSv9KZgG/oBYs+TvsWJApEtggINk/JsCCePPLg
AIivGZ4Bb4yaSYCS5cgcumC+1MxBlNNup95kIi8MF0TAAp3LvENSzUjbhBCMjpBC0Gk4wC3tjVZu
s1D/uwwS3Zc3IFZBW7mUdiaMilgTI81DeS+EjSl8QDSwaGhlW7wo+KEHCaXwy9RbhzRsIOiNenvk
FegUklLzfTyaKOwKcIWdFjdARPKl+OGHtSGsK27TN29JtnwOiK5Vn/TjEqI8v84hMkPtUSCeTv2Q
vu/D+Dny0kojg8IqzhTOvyfh+Srbv8AyYoiF/HvO69j47jKm57S5SESkKZ3HRdC4yWzcN9G1DwcY
sx00UP7SlhYOfx6ER0TGC/GGGiYoPL1lQkAAIcFQ9EkwMEn1fKDruNFBrQiavT4h1uNk2Tj5jnDU
9z5LZHEchZ8T8eWTC4j2+lw/wf3clOWIi1SqgUYVgNqaoyh0IbazqGOB0vk5rRsRnGgsTjuaiQRZ
v5oMKinsxC8stvFzX/ACKbmeux8878rj7taEOwJFZIOzHQtWavMN4XDzX8TMd8w2SNqOhAoGo8vT
LUZfD0j1Y3+TIo/sKYFcY2mDOtRkXo+Olv31f1csGYgY/NHIRK7QAcbxpNjiEf219tUlqMmJsPyO
9l0Ht8Sv2Yn4toR84rrGCRLCDrMtMqN7VV6RvQw46P79WL/7iWv0IIW5BBcC6/olCzXmsnOzSQnk
Wf72x4lo8zpO/QodyFtzQhxBeNmzAzA3gMexbzRQS3502qxoMxpyoffFN4mcGuLrL5ZOBCYCZOLf
uA3P+glG3E2A4wCaGRQFeXZ5ctZbgylizUzS7c8jtTFdeh1sfgKNmDfojk1LuTV1HbhdoO1OfI4k
e+VIZ6Wwefcp+dMrOpWR+d9QTVvlKf8LEyGCFqxKrvqrquC2PXHYPqH881gUTfa8/My/9LVZdXA7
4Xo689wLHh37i5PY67l9wW9DiRzfL3LX5nqO3I5ZTbzAVnjMrXXolVqILxT2AXju7J6Yg+Ew6t/S
29bjq7uzsXOeyX74FRjIbxwt5ZbhygVWImYRy5+UKpY02EUGioNU8Fi9YCYvbd+/K9pNiTmqL1oT
5QAMfFLbRqshpmWj6wcJ66ft/D0LyOIOreEsVWSHL5n7VVo7/Y04UdiNEzXnq1wi0kfbI/AdCTGx
x7hc+H49ozW9vBp3isnYT9E1caJsBJUQgT59UPUSJZPCEykV14fmrxWz5bdWQJQZLmLRuaeMDlZ2
veuFPVuHYbJldEMv0gjb9EW2n8auUd0Rr5lxJpWfxxxoOAJn0se9nTsK3az9E6LW8VrpYktQSrkd
ZE8xN9yVo5r6kcAd3QRHSHmBXSh5nZGf8Ero21JExpHbQ2SpTNTTWLiJ3ikinyPgtQAz8bm/J2HU
NRSIyLms9F/3B1wHVawYidi2atcaSL3xOaLjar7FZj11C4f1l+vRdJ7BMeICYniphgTUAscG8rRs
/8fvi11NjE6C8bm7oZ0NnLN0sM4Kow23tAyWbMLFVo/kWPytjL7gjzvYxANlSdCoILN5ZYU8e82o
bVVLnGbRUXdxA1dBRWCha5AGN6gCPev6yLVTb/BTT57SdfVbca8goqSIiZR52gDsDDeqND2vo4ST
HPtOfFwrInCxdzKB3fIuIshuKT+cz+dRzbVBzkjT9HqNNNtXoonaG2prZNAyljfNTPDOmCiTb69u
cRPEMt1Gb9qQ/X0e9vNt0U8gaQl3OPeLQ3COiUw4Fo9kpH4W330rW9ZbLonmjgFHRsm3Bi1NtJAF
bL96sjTY8pWTqk8WvRPZGIy9IUsqeexhIKCRPJ8AUodwHOYJOwtvcZFEGthQXcrMNgAziWfRyxvS
I8ruSa7aIEPrVb2yZfGbGu/F/UO+9MPC9ZM5Vy8XrpjnxoJ/kqOVpLirJ4+74xWRkA8y1nHY3z65
NgWbRIlhU6uRlGESJEieF5EyTqyUGSxVlqiWQ50Dgi9y14+LQzdSeIBhnLI19aiUg0RzaVZOsVCM
TDfTush6w1V1A2fLOlBBZalT6NHEgFceUQWbTPhGq+cOpw97Wdjx+IpVhMsu1J5uxQZn4IOFxIwQ
8tgOo3KoMje75gkN/P191qb0fevUM3Fc7+ofTOaHZ3A1CmLglpqHPnNY1VYuVxj4Ds2CV8H+WBWf
2lq2a1z07FZD0y2TC/blhLUMefuZuWlHD26jKt4wSNlJUSaJfgihQVNqoMF7eY7W1BGgbrTIj32e
vP6f8/t5C4IDSIqz6ARfs51ylsX6Gm/ODr/xT7VvxqE/BZjqA4ZuIsTsRINvV/aLVq7k7R+tw3VI
QXGm/QbJs/I+JIUNPCep06qEG46brPfMDK2CyCyEO15paU8kKWz58DN3a8u2HDDCmPvjPWp8rcNX
DDxYvUricTxlGpeFYDrlAEDEWHQJ/ZVf+jQ6wXSOoaVQVwq86auFSuFWULkpxmRE7fvJHOf8dO0l
D2c07a+UG3s3l0zaahdt/UBdwcUsE2BD8sTCgkTFXhMp3z+0Tnjv7u56gldD5bpu91UxQTRTokjn
rFPQ6G9+f/dMSrq/CCSg+TfMROMgm1QQbh6gamrYcy5UmANSdPrqUAA3znc/qBBXCvuQS4oto2lm
pAhBPjJYuZ2bhePrxGE+KpZWd2YlmP97GUVVdopIbSzORVnK52x8LUxs/DZ/3EfV6E/vSCJUgBWl
oJ+gUSay+25aawC9JfNsPMJT03zkTL12dpjoQpF11QI/E7+oru4qo6emF68THNTd+8mLjxpbAeO+
n4ziEKX6YS4jSxt/Xzd2k2aFWps4NWv4A2IHWXoPP/bx871vtqPSyW7hjsmVRisN4m+5E1NU2uQb
OOAYjOey4RpCfVdUkwTld5HaXtnA8mU9TyeImgewp4q8lp0BZySd/isBQfsf5Ume4sioiTdzSMkf
VzYc4TeIVXt6saXdEONBWUheXHByxIyQZkx4Tx7IgyruJhRS5drsQvsWF+ozcqsRtaDeAyLTSe/6
nCPBDd7mLpnPlNGatOt/kQTkpe90rkeQ2pHf0zwB+HCwNpqzJuWhjQTP++vj6X85iJHjbFavk5Bo
P4K2wZm4LcTVcK7vronBBpiPRRNJv3PQPLITjgGVxK0uv0yRXFrA+is8b5Z/PFIGYqnjM1jMs5SJ
hkSyGhVGcWN3K4/YQTDD9OOmR9ZEXuVKR/fguvyBUlplGFr2I8YqYPSR18WMGCjqZuGSehF8m20C
2LjuAF8qea6e2eSYlT65rXmOdqu+5LJItRo3A7m3ysVyYb6I0pQ/CU+6CIxIGKozVL9vpfV9wQjQ
RNxb9OKZUcRshhJNu2fLGfUpZwetgarP3r47RiqxpaRZIbz52yyRuRA3kiYFwqhub98HfBj5xhoy
FFM7wyMA3sK9I7RcvdT9hVZ6N12qhG4+A2TLZ9UPw8bbX3kXZGluogUHCug7P46Yow4UX3Tp92jX
JgPechwTTOIwHfHy1FURYlJUWx4ofr5oP40XE6/TNIv7YfJDlI7xEUdcfknhAgg+G6c12ZgRrcks
+drUih85I50FV5+ZGa9OYWYkkWAuhMji/4T3on0lH307kS0ww+GnbFTmyR3cWPAoIVBT65t3dfgL
Roz/gzkS/1LAafrIdYhS6YfvDVYGforxc7y2N/pIxo2SjIGnFNewWDcXso7zQjjHnoED8dS0Z+sF
ByVIeEGYlMkXUrevIQinfh+V6Eq/lIX5vfDhMsPXrhSDjlmYGF3s0ER+M2ARanKwc3YXHrldxWbT
uRW31R8tHNYAKBSn+dnU0ZW+g2ecFoUjVSx43d04o0MKbywXlBMk0G6RyRigYH00eilE8CHHiuPw
0ahsnFpTWYZJsNd4r5Q1WmJHkYEA+ynNqIQ3hJdpWXtgbRuoMyxIZPfgPlwcn3cKUQkWac/nOnFF
4e9bSNz/3yeJPCfwZAZrdK5PApZpK51YiBKd4HA4OBEOhjRREhlkSFlTEJmCG8R9GBSFCp2mhxSm
OJ1npz6K528I0sfW4A0Z3sjGm9qG4+2fCf4WhjlVF9MieEh1TG8SMpryIKmMPn8tLhKalwS49c//
Jmbgza/5UbSteaAnNHlJvtJyLeoI2uAiK/gPrs7EsiQ9SVJTeR97We8ojjz8eIW+2VA+We34bbRE
Po8QxTLtCkFKWFQ56g+boXXSpj8MufsRoe3P9uxEtnHQ+Z+8r50oRcH4N9dCRJVooJGBTVs7vB3l
Upcd/BMcY7eyu8LDHL6biePdTU83b6p1owzz+9HOf3DFC9x0HiNn1pMbH1xYVcAsGIa5hcf4Jxfz
hCpawQOB/qOGNGloOwZA7vSLrh4Z9oqcRA8OersysG/RAvIM27UpXSCBW2rFYQn6zxq03KNHjlhj
YjiyFGc/ZZFkuUzdcH5Hv1VJVMb6P4XsP+CgxsY/Xq08CHS+IeZrldYQz3KC3eRCPPCiZKRN1ICo
fP1syC8sBKKeOrzr8aCPlBaI56z0dZZiyFBRI95z3C3FbyNVErCuVyAffnQPyghNvWoZK+ffCekF
vup9eZVsbc6CnbuRj/SE8ys6XszBRkD2obkE/8W5DBQwLYkiRCPV7USEnd27pEP/IEu+acog0Fjg
TC5vKqTggQHPBJ+5mexnVDaM6tFJ8Q7vTNUvsE5dQZa+0bcJGlNX4Oq6p+ojtoed04IUDw51PBrk
MDmxtdjzCiS48Sdd+I8yIgD3CLlJEtRCKBwG1wQfT+FeHUXayYspm1GpWctGFUsNK0pas1EM+FWP
N1Ol+ALoxniYKUgQpIMRV2nI4i2KYtLxGZnrZ5tAGjejheCAMHRKqPL+dYQaMojv7Co51JiC/Qf2
P1WWwBcY+Gg6H3YbTPmF/gKsj139h914Gd+g7FAC4iUOkmFWlRWiMk554tofF6w93T9dKz1cBSRi
J7/uapovMb5oRXzXLWZQULEVSbOIPT3UwpXHgZqRhOViFKWhpdjpvtyi4JoH2UfX3GFdkctPG/sa
lU+4CJhzuI67ecqIuBvwO3LjXoqpixEo20cJb1tCeEf9pwENjrt0LMT4SpwtNKcRrte5FjuZg9N8
2ngyoWZSiUO4lo+oWurjzfSMCVLhbD1g67cNjbZTJEepRpklcLWRJhDQMDkX6jlDe3eXW5oHiRVd
ZycEo0JGSWs79ob7XJH5E/mrgO84SdWmTKss/slZg4tP40lPMjX8RP9VafWwnDAXzSAqjKyO2Z92
kOpIhH6TfDaeX4V38gWoKQO/7QaPKCj5ZKyVH/AgafnbzxbC1E7I4GY29UD9Fp4hROC6Ut1oByYY
yNfU6hxY2aLe6chZiJH/BgndMXc6LNOU8k7oFR74xIuzEkG20ytQOF0BXuak9cmbItoUpUsYWFbr
oYi2JKPCVxUW3Dz2y21426jvjNT/V4K0WLqjLQ8QiTx+hH5lUt9CsiEEHi58DEKv5rcdg4dHScFH
isXsavK9SeCDSNzr/5/iKni7hA3bIV7XaxC4rdldq3dfYSvSE5eW3/PLTMkzUt1jIZEcfVQqVGLf
DJE3f9QwMLtFNg1rAj6ImmL6HysIopZxJhydbXPb/Mp4s+9ZjhGA7hEHjNzHqfnI6RPo2jpMDPvi
kEXlz5SV/I+YnFfwQ3R0hewzExklM6eMpcnpIB+Vk5DcRzK+NkjQN8U1DSEAcOqVDzvXFBSFQDRO
vyZfgBQCnQezqMevcB+hFhT7l8vgWVfTuniy7UBcSPCbWcjMnazUgGtnNmb09Z/1k1HBrtq7J5zF
ARA7COvN23Zz+VndQmP76qeCSmGqf4O4IRzr8YIMj6iTbZSHSlJv1VZNU5keB2aAKtRneF++s81G
6rXA6ZMTcvXF4TK4THWMA1Qa/1ApHwMHyYIeSVCoHqEUCRLtd/ja6wULWaVpMRlR6SNfMEjbfGZw
6Zosyy7z2/hHu+fEbxn7xqaycgChDMtKfgqkz4kJbcO7R5STbXL6m/NxtR1y6XHG/0wRBHR8NiJd
xwCrd7Q64LD+tbOauq2LQr3IoWqHSkyQWwYymvtgEBrzhBK536FS1E1CIx/BLmuExlw/bdCQ1KwA
0VNfFI7JLjnu03SlWtkTathr4q41daVUNdfGX6mCrkdE1MnpQ7BDJlUPVNTCByvmTzkdAYFabRp0
7vp3+ApFDXxkVAS2Nb4xaHdFZTnc2LtyMC2eWt3MAqBIf+v8URRzNjesyP731HMcktedTNhcvnSd
5YrB2P0Rlm4ifbz+o1vhdYDeHZ4Tw3EG9TqUu6IvuJZ5wi9pPpjyiwz44uhYLYw9gcMURb/I1Ubg
Qxzy3KnHr1ZzTFwPnzD46hneDXkrC8IJI0XfqrWEndQeoCXJSYagVwDeelZkW7Qjv03oGSmRPLUC
Dzf9hrtM7RPsL5bibm3R0gSmTebDRVUxGCmghBbuvYipoiebiu6PuUg2Yc0LCvI/CH7T0Y4//+ER
73RmWl9Rlm5+7KnF0IfRd663xMJ5Hgmsjoc2mnGjmTQmo13qW/1+z+YnmcNUTkulrYTY5BbanLtE
vusapRTmbvldopSjE0qDiad199AsBozVxx3UYI8UpuJO/DShRuocIo/UuQ4H4z5Wjav5l8QZl1Cw
8A3ROyzxL1BvCWG8uBW8l1OlNCHdG+yTkH8jv7Ss3FK8J6nFpoVAkiAgodU1Y27W2gmudiOEIzv+
iyYaEFDH0Z6XZUuUiZsMSY1wmjS9d7WnNXP65zwJru38pMGqjjN3NDHqQTFjlk8t122052zO4uAu
NU7NZa9Mqa2RT8dMf7o0RDbhsKZfY7EP0w3y6HTfEiUl08f697NdNOrtryuDB0NmNDqBPmIyFbns
4dMyaUqNsBUece/tR1+kT2uG2v4uNE8O9nvftmEzsfY4a8xSCaPIQCN6V5L4pz65qtYOOsXi7n9P
L94NLg4dnXUom0OciQnl39bKzX5beV7ft05/EkEEKJ6IPXtw3rsHA3HW2ywSc6PAxdMDqzk86o0f
nGxJI7RvzUA2rMVUw+QoybaMjHDgfxsQQ1LWs9ym4ThaZXZEICKgYX6uUM8jgaXsODTP+HUNJo8u
AF9RhY2dKkXCeJt8EoTbQRV8/Tf+Rvre6RQqytz/LobNuBEHu/v8eDerQ5PoGkuucIV3qmhxmujr
4Y4JiUXE1PPphdwmnDTNxxy30cm4gHonvjJxkOQ4orD9OuSU8xgOY3KuVYvy/F8h1sIWTGG5KfNR
c+4Fbm854JGqcAhUYf9mbkIx4d+e2sGXSAg2XMNeXBY3meukKRka/tw0KQZn1oqAGjFJB0XGQZ5R
+0E7j5Odi5krOmrAFRvi8rNZLNbA+vUTkqN1cjqXvVa2rP4h0lsl+PsQF8fx8Ggn86QRiTk2oygQ
UIhxCblAxZKH7KxG3m6m8VY5QBzleG3+QRctpvDEtgUJuUKfDaTqeg5Gh5QixOtg8dn+7uOV7ccn
0bfuKd81nxW5lvcLfAskX0cybA3c/G9rgefa+EUZ43MNdrh2H9tzJFLeA8rRPvTY6SkjOMt6RSqE
oN7dg1eF1yieyyqW+BQmvwq8Ybmu4LT0GvGjsFttxjkU+aCi+Ls75SXIvgn9TgOVM79WcRJ1CqSe
UshTfxmMaT7YFXZkkyWCyK8C1u8YhnpP5AV6O4++qUjWZa6aJVFH6gUHm/FBAY3Q4rJc/tX+qVS2
WWslDDdMXlnMzjxxsd1IA87JE/KX33TNrGfeWJM0kteuiZDWN47wElAB/5OGb+hNt5iB5FPRWi6s
61Qm2tB1n3O7iY3P3CBeE7BHUh/45lwuEO92cpI3Yt1CJyr9zVa/IjWPotyR2FdOKvVT+ZBVQ9oC
swM4L+TCEToRsL+BsClO42i8Ji01+XiOzs9MciFVcT/N5u2xRuiLouh9F+qRR6brOgSNLaBP7roT
Z25kotkPu3EHgrfEPQSquPlZcz8meVVc74xZPSyzBL9m36vJiGxEmsXzEzSQGcXuF6DIZAoAVloE
0gYIactcDE8vbrYARRynGqTWUF7PNqkKQGE6nshQ4IxGrxn10sVOKevmQrr0j1Co2zhlP+/+pHHI
XXR2x1XK/EMxuToLVeJMKhEtTQWeMpDJKaOCeR7m6lOy7qo3ZVM+H2IU49AxHhsoH8YdAyEsc+s7
3XRE/OoY378qrTi+ClyUBAaDMK6yENcMmY28wZj6DaqC3eTTEf++Nc62UQUUbHpruVbQHOzLZ3f/
9jnOCU+jE4xAW+8G5dowUJSFPLY/3oPNHTqq5v+0B/vbH8kNTnhehzTZPO+LUh1mlvVC9W7bTvMY
q+JkI3MFjc96zPyt5BZgCEF2z5CtQVGsaL7y63vQQQpgHOOD6OFcC+oUWGe0BNtrytWlRmKlvSYb
97rbICeaTO5fAByXt9ErTK8SbcH3x7qoWy5UBcLeVb5Ea+WmgV4yaYCJk9Z2YQvuMnfhBYY8NhDY
6Ak39nm0jwTrwKwoV1NjCrnT0xhfR1Ah7+/6lfTW3t4RFYdTBh1aENT9ME7/Tz4LxODgbFj/g3Oi
Wdrlk95AcJhhRVUxv5YpvPns0EB1sJmiYhMdkQal76TBvl1TJk6NANF1Ek8SsrFI8W0RKWbGr4lX
Xy6n6gETbKCG42IfUdpwhhIYp8qzpENg38voEeujJxE3JrSKeixk7ESLBF6+1h7eN0nGws3w/NX6
XSAx8uQqjta63Lv9ywvClEPmvirjtHptDt4AiuzERJdUjTgD+KewplgEIKg3DGSgDfMLYfBz7g4S
YhU+bguJ7eLO66zTAkSWMRs+UrnA//UeolkP1hQMWMCv7wvVLGe66t5uzxPBzl4qQYpge2XAVnhA
BDiThEuX22i1qeRXp7VnviEVoefU6yKN9ZTTITQ+wMi3QlO2x0xZaSxAcpfkbkr1esjm9W12UuP7
ycmTse0tGM/O5kUxJNzEZ+IuA9MTkdaI+rbe0O7oT6wAyvpICaL8jLTPujQu0Tcid87aGijEHOoW
cU/rRXUrxGZwLkWaLdCVsiYmEkvq5KC/l7zSnYgQKQP85G1gWrzs1nrOtQTcUBXKBFqFVlqG234V
zt9WVIvwKZD9MudPKDiTXvJqXl18ykmbnAR4W96gJG7uylGMCRZ+GLdoDxUZJZD/M0+Nconb4hDF
nDVYXHKrJA16nVMk8eAmhH+htqwxuTQ3oKnltZFUWyfQchB7rZXeodeNLQa6hEPqdUENB7JEdNo6
g3Vkq1bdf0JrHCo1Nkgvyjs+w97P5dzdJEyUChZh4B/7ckNtbTsHUlK8TQgm2ZfEmH6FpAF7zZcQ
iF/iM482Y0eAXqwBoLNLugSbBMfMi6KbJj1pwFNlS6ug/KVvSdG5+ZDbntMO9pHCRXneDxtHu75o
WTOv4T0RUQ6bmkowJ4PzmAPxwTj6r8peQTB6QIU4JSMxSF07wWGO9ULfPvCk8rFVOPqexNLZx4zp
mfN4F4CXIq6mnkoqhZKECrExCO+qwpf/02SV3sghXectcbnH9vJQqU/T7gddc0z7DCIyqLqvNOrh
kdUZyqrUeZKkx8hjFQ94a96D31DSrOqgEMsjqClJhujsMMkHms0C7GLWWkChd+fNCHofVCUzUgug
i2qClEZC3fOO5YrwJ0K6ud/EpcEK9zPRKXKnAxWnz7f/xXsaBeZAfhvsHCK6NiUIuokgt25e40yA
80OkA7WRXtsX7ZclZYgPiAM7zCXhHJvDpAgfhcyQfFIw8PY/Gh0jIYAqjOpY+0m6kz3XxAXJxRI2
PS4/fRbhCHba5aTDEguKxjEQZYaQ+bLhq6uKVhszkXzoo2uDsN7+OQViF1y/Rlt9SaEcEGd77Pmb
hcEhlk4TIJO6Fbsvs+FOQR3CbtzeBYp++M74WQy9KasmXZ5t0CtaJT9zCqMp6lmK1g3JTqsIbxI2
dIw5Hcv5BEq1s23xF8EfR0DnVdNqPZ/KcA9uxsquT6kzTREx0aZ5plp3CBrEFFYAXll6YBqRMqOw
yObi+9VBywisHFpypQ8M+kc57LwQxmQQ+s3+grEqrhxhOCMqfSIYReK3nuE0qV35wQW2GCsR6aLW
zoen72jNPxAQckj1XAUdWJe5TUBg+tcYcQTpy70STzeqrlcsHDKhfA7Qm+OJBUQR9n0VnuO7m1B9
m9TjFVZmRnv7kGWtWh8J/kuk+/PKG+o3O0JiLot3Ynh2R1Zq+7YAqOAQbY+DS2tGvuRW6FWT1ESH
BHA8fk0dcLwM9dTW2/vk+7f3fWdYrOd/l3J2Ub6aRJFbDVDZzu2/4QKrILn+Vp8Qsc0Vvj6NdSdC
Lsy974fZqtcsCM28dbpZkbd/BJKFD4+HfvQrvofnDyBHLA+mO13v2dth5JetNhl/AlRf7euHf5ZL
A9nBzTOXOysMg/dwhqK3SIfzGaREivCikkwpjQwH3E/RKgRQVBsys2YHe14IV8Y9T1Z0vmtBlgno
R8VXGxdzQ++HNWfHEYp+OlsmjFeT1/xyg6rS7troRvIeKNuxqnZmaxkaIUEh3VnjhtO0swcKjtmw
lu7uGyM/UInaS3T06gabWPIIf0Snah34AQfkxwRSZPav/l33Cq8DHofz6eWENywYohw8pmxSinZ6
towXkfuHaw18wPjgASK0TNz+X4osbwP0Vy9MdxJVIT1VHQEfbca2Z4BibiVkiR42d7npf5XY9ERv
ORykgcFZPK8eE6s3dhIvOmkkLRWRfI2JVk0cS/DxAH4Xj7KS4RwlGB4BBg05dcaUWk/l7CyQah/y
6+42/CXGlbG/oBWPFHzqp+j0vhKcHOskn7fKGvFIN+u+ZmWdzhjfg19IGxnWrx/utdSjPqy/9k6k
7IQE4aBTZCq8FE/ffMfzoN0d7uZ+od/YByQihUYlM3KbinMAELPDPknud9q2ZqSxH9G0xoQ9DSt2
uSVJYFol7Y2N4gutWrcJ9uOEov4qyJAQBZRaYSxBSYf38yeHXTTTb+kTyf/zkaL4R9mfGBUY8fz9
Nw1ET8kdoMf88Ml3Yy1xYhUK6LA9geVvAC9KKoMqVxKuR4BTVOYRso5bfqsZVWUm4n4dLc6wc3E0
Qon/9z4FcNR2oE8uEfhLPgn61wXwVwEwP6Tbst5MMjA9zfRfbT0W5DQmOKyVG+/x40HbmdtOuGOH
2hBuPC9ulHVLwiXryHn6+be141TZRQJtE3DG0nWvyD431zohdG6VEXIrT3qwQ9TV+Z802QLvwBxX
wVm73w5m+mDzjERS2FX1kSiK9YgZwTVCkiOHVj7fh94TikU09jB2CyuhQCgjtHRjISMGOQyM02CN
bHd02p7kowKB+kcydLnyoQxO28yGSfzYrDH3jJnVSKcFXEOrPN3iEdErHdZ3ku0nQO4DUiupIauq
l+VcwcwGesf+tHq7rwxBCPX+lC1l2n3taxvX4pfo0/MzZ42Q8ADak0KwreLbkQZLImY8/GdJRu13
/pNtFizr//u91KGTGkmr4OJBub7KUn3ptkkXZw0+hnaVFXPjIpcDSkp/PGYF97rAG2MlINujPU29
Hq/gB4bvSafpL3S7UZQ2pzS0M4S96DVuRBBOl/zs0JbrJdDpXGzFSVNtd3JgqAzObK+lLmk+9gzV
2rQTK7GOZHPFwblBF5C2esLzJIApoIM3n/h/8gjVOhEq5YCoitGFGywftfpva+dQLYCzqexWDvC+
40rM1Z69+DV+9wsha1SFilMCJpE8rS9XWh4/2u76/K4/qI4X7m0ypVayILEe7ywb3pSBpd+RwbdQ
UGZlr29w9o4ad6YxR04BczDPEISV/o3YpxC3Q+lsxULlo89BdmmlSb4ohb2YJgnlXPnI9XBJwvPw
/ew/qsuRNJR1tXQb/nUrXlwuy+hIn9+kfqsEEIsva60cFoCPKqIcjij2pwLKDTvWqRMVobyTEsyk
Oh5ZyZaVDDY/Nm2LHegbm5M0ny0PPRcNJeU7lR+Al+vjSXFAUJyjxy3AbvjqC56GvIrk+yXpNR5p
VyrpMqEYGLvkCbBOFnB+5b9SCYHVkYvcnTJGKm6o4Et/JoRl39PuHn+slkwp3QSk6mBlkCaOWwjW
CoB3Nzr0EiYrcKAu9MUzkmzYUrstRDTAtbuXxpZRbdcYystkyT53ln0jStLn+tmRHB3ktUtWBXix
9UlHsgQf+EnB4IP6xY2+e++DEko0m9rF3i6e39t3IvS+G0v0UNUaNvikUkG4qc+u7KSbIsuEakuy
n5y06E9KnZrpAjElVw+9u1NjjhixGbHn6wBfk3yBAK4Ib8y9bfAglt1HbFVDGzRQftdX36n7wMfM
r83gF6vD6ot74Y/YwhI47LG1h5jYh6pij3Tpo+gIUsl47dg0PJS0CeRYKEYaXtikA5+nBe2TmjXa
g7zHGMhVs48h25uCj4+/YiYpBn51TcnhCP0XgiJZmrPfHv9YhKk+rZQOfGPR0ckthaRvBHPeMeGX
p9zV3Pfc39M3bSx3iaxtrhd0nvkb/uIEeikGwte5OuRNrCV+/7SbdKrIrelHc3dxZcnu5FDK/K0P
gJA6y+LYKGRsq1RF4OF5dqsEM0ryW0fP9lZw/rCjm72BnhyCGBnI0DaLcvDORKG2ydnt+9Tj8K9a
BgHJL4isKFg6ttGvFRszC9+NwxvjdHITu47SRRHDYuRWdVu+h6LavM6S8iFMA+WA+4JAwKnRJYEs
0oBUddGKZhBQsgXdfsxQzIn+/NR7WSGMhzSyTgI9J89YiZwZfxEWtgxPukrK+w5NsHpL6bT7lGxC
x5c+BLkTa6zWRfXWExHKC63HKdYpSpyb9+sYwH5VZjXDUs6KmloST1G12xBI1DSdssNoewiVQIZX
OyunxnBhEy/0si2Nr+AvPT06Ua7TQ9STNFRzA7BKugBXnqEoBYxdU7SzE/8AHy+p1mgixBOpV83J
SPNO2+teuNjeZiezgKFah8f4BpcU5JOV9DL/B9stXNy9gqp98JzTKIeSxwEZ6Fr8Wo9ZAKDTH1WJ
v30GY7y7HoMGDHZOgL3/wz7E01sQTw0K5p9qbn1BJEzZDtDtpeq72UIxrIbNdGa04FvLLh4Rh9EW
mXN1f1R4SxqQLLgMC/XHR+/BfYJRRbLAyZfSl4DnPiM4P0KQy16y7VYnvfhbrDYUOfqztBkDlPmg
+92653geiGmUFSMeSM7JNArXSGqeYfatmKUtAZKVQNN0u2jVDqKUU4mlu+MwdZzFVPbzcMQmkrRi
O1FUSyMpoJlqJPAg1HuENhNOVk4aH/u6bpsVe75C3mI1cJa8tA6QIzOnOzPdz6oUoOYjxObqVptB
QN6sxRupwToiWf3AojEQY/dq8T4xiusw9kQPjtrprY+bfDoPEB7rcjTDq/NX+ThGulvbUs9Hv8GS
gZ49cXq1yYhsKC7I3gJ/vBGeyiHwSiof+gYWqzccohgHLU752/RWub8rSCKsGCX2Xy/7g1X4IdVn
+8hZPMzv6YUD6yYct6VrucS2O3CEOW4xor/hzouUtYn35iEH09Snt5qRFkQMk3sUkYPFFBtb0qEi
ytFjRfdLTDkxqBvwAgqCb9TJKEengCtcRGauFrzFZSXx4+uEBTOtoJmrXCe4JjJOGLZZX1s4yoAx
GKBvUb/wOl88Me6IzfzPnbftw2EZgTK4YmV5peQRMwtovOdGylRE0P2m0zpYrV5WyAXY122hnFGM
RiBPWy+mBBHQobQuCADr7JAdKa4NM37EfemfdPWWJaoen4gp51layEkcPsdqkgTZBvlPGe6bF0gt
lKsCZFO+FwFH/V0hPJXByyF0w/SsVw8apk+5oWSq3tiiUS0bysAURZYVisDQR/7tEoEL8pHQPht1
MbhTwrHiA/hV2Xn5qMym42nRviYEiwSBTsuOgZcQM06CyRaJ4ZCHUDQ29riH4Rap20LI0JhrPsRq
KbUoUybU0epc816eefq8/Ej5uRdgXA6Ok4evyBjoKSoIeTnAcEKSSG+th6BcZsFckFZIw81uhXFl
Ovg2ErQ/EOAvTO9OHrmf8IsX1ZVNX+nRQVvuizv6IpJNEDtuwOaYfmFdLedmHIJNYKflBfV6tVyc
h7wv9tCFL7IIMyw2RaDQv8dDPVSZiOvGML3HtbqvNsHsUmpZX8fWaj8vvbcOEtq9h9ZWuU0t1mIM
B+Nq0A88fcNp1LdYv4Z3iUqcCHBl/Km5cWOQTkNul9pk+r2L1yahhUsnOZYcSiTxHHgzwHzfzbZh
M/d2wevedZbrMlaBAmZa9TzTIDpigSuRNWD5pc5bSngcH2wYFIuk1RCn7Vivz0eGrt6FncA2PP+h
ziUbZReHoSYODlNrnWrXCyZlammPZwfP+Sm7UKz7LWCBk217IxtxZKmJZs4VUmM9F/XSlMU/+VYr
+UqdARvsY7gLK9y+Z002qfTE96cgxMGEljwf6c5oTQlJp842XCu7PE6gt9vA9cnjYqUVq3hguy3J
xqPVni+H+UCsw+59znyJgcTj7mQtJyhtZJ3zcs9CWM5sJW8G9xkqgOAtNh1DMKxTdU0E9YvDDLZs
I1U1F/8W8mb3OP8hQwirXfcXGkBc6hB0ofNiT1c4cKjJwqwVWcjPXIrwsUxxrPtCjqSekRP6+hJD
ZYfRi0XapzY3xyGmaS13DOhreVKG+Ill0+TFGQkljBjp3JqKq89ZMNS+kweWlRhFerABmc/qEBWd
KsZNGGGb5D0UItTkQuKOnpS3o4TayEjI3uekGAmUhq8/9W60JeGQNvk9VeTIGAB/gbxyZc1mTBTP
T+o54h4fwXZ4bVMAumnkVl/JPdHSI+EvuOo/lbczLC4k6yZMCBvXRdjAvHlaB9/Wci9EGI7cbgIQ
+p14mUzUz2nwzhv5u3Q+DviUAeA7bDhk75GZkKgEdxWSHkz6+yokV2Bq/s6tS1+Vi1rI+XXXXzAW
D30ZXMPKM4rN2fNvf6JGsWmGQ5hATgQb77/rDv8Vdi9Ce33clvKojuC3Oy//N+lWsdDfuqLgYqmF
qT3uJaiwAs0kwihmDMLdox6HFsFhlKexQR+G1iAMO3prMH0V6qnlEIgW3w1tRz7eDgsOFtSUoDek
eocQ06Q+MlnWeVhEdtPtIGeVOBWpeYf1C7Y267KG5NgNU4EgsZs9VCcurpUL5oypzvqt0E/ozntP
/NZ4ux3/C1cjbLOhD/GfginN/CxwSzfmIm/FXoCirBbXGKLRXTN1ecskX4Ic+J2TC5/+q9HfP5al
rbUV/OTS78uJd7OXpH/Uw8Ga2oKoWVBnykw9cLIY/OliiTqKJVPTEk3rahR9hb9cmHJoLEPUs1Rj
NXv6Ts+Cgl1o55V3+F5EC42VGApagGObnYyKmYSxZ9DKD77WIhLVikwlhJSBuZx6iA7PfUH4FW2Q
JfFCeSzzg+8W42rMg1+36mmS3iHxJilD2onUw7bgvAqjjn4qC2mICQQuyZmU/3Gv1YhlZwNs9JVE
ReHCZBYwfiT28X3DJN11UXM9ZGgri6kHP2HixJG7zIUuzj8zGDe7JYn2CYaMB4BJM7SO4G5xZYiZ
xVV6baIGBUikf3vidjgTyZVcsPMpjouQuK4OLXFqaLo3PF7etHQZWNI/XMppgVXWIBGs0NBMOeSa
LnboKgJkukbIBy8EG6BUvvMd2cjlbv7Bll1a5qQJGZdEbgFXfn1V0wL21DM8mnal3jA+bf/Lalhb
aS+xppnqBF04MqjfBo7nLpPov7hSAUVi/TpgrccRUwgYdLib8DLKevbgW5gKVaq+iz2ildBpK1OK
NM1dROSiACkIe1Swq/qzAJWa3gyaH67LIGe54CwlkEVUtFM5wbXmZOf2Iy9K6NgeewqF3UaLeze1
6+Mi9jzGr8ZgTx42jN/RF9tsER0yQqMhVJuUwqkLepWAN9jnRRRiHfFcBpkSFv6HqmHl61MQIXhf
MRk00pl+IXwS1LMzRTZBwMo5FjhPGjbI+99nEyNlqGVny/Fdb1L0QxJoJYUrlxaohfu6hkiUJ86+
Xwd5f1D52lHIQlvBaE/ORpz30WMrn+65TGVhiRttoInEGIJgglWwyy7hrg0uNzFf+PJ/Mb2EoYjl
0q8W1vg5BDo6UUh9d7nqFqflDSrarqKngao/M0Fy99MoT3ntBkT34O6IYN/szj8oWS70WmG9aEu9
3iYXuehjvNltwcONuUrhS86mpab+pdjsdSF6iPoEBw1hiX2ASiURmKo9wFOST2uD/c4BIVweUCZS
ZFRfH5B8zyCWFsFjI+lcY2QC71Y6H73WcbcV4mghi5hEL6LubnmJeKYV1p1YxGM69p8h1KEB1MOa
uoI5ap3cjfs6XxUa0v6K8wmZoETOAyuSXe2CCXJ4d4s5H+v0ci1388/gzMYEgTKwzClCdN2Gox0b
XxfOSgIyOiEBREPbFxdqlY6pb9WQTxywzYBNm4iSGKZF0dnIpQ36zb5M8E013eS5fwiRxaTX61k5
n0HvDg5/R2BzYQRY4/iv4c10gcxOIRYYG3MnbwZHmxUXjgxx5yXX1SK1spwCD1oAjt12xEuvYuus
p8nwIBE5Q6sn5WS5pv31o8agguA85E5ff78i7nPOU2Vig+pjO6yaKt3FVxcHJGyAHJmJ8eXBTZJ5
9PvvMxJB61LiCgCa8mtUBYwPf47a0OBjVYu6NngKkV9gHR7aIMnXqZg7OSFSbadz4iyr1VEAihzc
u1kzcx1tSS/Jr3GdLtdZq+W30Xi9TcbSaQ0YE8MFCVaF5otQ1A75SYxGpCYDTi6isfB72jMQjJEe
F5g3PU2VZBkdO34jkA6LCGuSbZkvxSR+W5NoDIQlSFCO6EFPj3LxcmOBsmoZoRWJ/DIel2mWGnRY
6KBEZSkzv4QrAFhC25eIUYtm0Tgt9YwNvGyfaQ5BCPnoQT3SASCdt2iVW/Q1A/vAiKUJsNDWe6oy
QwTcW+ZMO8xNbGGB2DD1wqdryI7rYtS7FhZl+Yf5HhRUBhPOgFvZG9ctynlZGJ+L/LvvyQn3mKnt
Uxsa9EpNC4O3iV7SITfZp08SahzTBbLAPWC32gpD3PQXmsePwskXBtjSvIwN3u2nwcwwaRk2MTM8
kFPAvvTtqjzx2tPU5kt8kMPOzD3ACWADvkmHHFeZ74WHoibAVhZs3ugFZKHEloaEzzQqfhC+5UCL
O2lLrgR4J3daQZtW69NiXDltS4emqotX0DjEMYUY0shLT55yfql/XgCbqFHqhxqMLWAYk5wTPp3i
AXJMNQsLppMuPJBkU/6jIipl4v8oa9kiau8wqHQ7fa6/LVvNSO//Pr1ZnyVEdohD0KNEzFpwkkfy
RFPlSdfVgYCbeVRFIDCqIN0BkwwbcDQvlloG0vq3Dm1G1f4Z0G1NykCePPs9khyuTpPQsJ/jJGlX
urIAimeo3QWhtTtCEakoYZlJiJNJS8/NxQBqNdthVBNboqN3stCdaJ8ekhzMpHX3zYhr4DXXEbL3
NMm5ZsTyYQZPFq3b0VmMYFdRPSLFRCVzV2CDWEKlFiBgxG7U0y0fP+72tk5sZBx20tXrOZ0zTkio
AScpqxBEc6kINARuyOxjlyT/1m6BMqT4zwnG3axyv433LcfoZskFFIMX3YsBpjCsq3r81gvJKDls
ERJ1L5903ys3MMm6TgnGJxjKc0I+u+I9uQNzVGJFvki7iTs2siHV7sv4d00DrbpdvLeDUoKvg2EI
vFQTn2EvokY4S9n8kUJQVrPWLPmZN/630kfm7OyMKRWHqVZQRAzDgnEFOYxxYWNmlrp0yvuRN7cC
m3n3J1LEQ/uW/uYaKGaRAZ2SYIHac1zAP8Tzx4WxIJV6+7FkIVXw2HPd7VuFDq2MZCxoVAMOAQ40
CuX1vrinBHc0reRrx+X7lWi2893WY72ttiConox6rK4ZIj4rmDeO+28rOpw3vq2uE4sQ1GzNdP4i
RduSPPyloG7aN9+CTUXQnJxoCIHsIOcGXUBl1h907YL4qwYQR8VkuEKvVDMJYTwAu/JA4NTtvTL2
wIAte6Hoa1Lm0eSKeQs60kLiwYL5b5Gja89RZtF8kmEl3jnu9mlBXAUb6p/eqZjNdh7C97gI2T3Q
599EJuw2q2DG34Z6VTRCE75QPvNurRBnFTpA3CfRE7/pNoDjCZ22Ndu9DTYv9JdEEVdzY7L9fAqU
cSpQLW8E9r5QkkVQfKx9QhbPC0+9XONPPnlSHHpKreKtqKH0lTsc5PQFbZ0/irBvpRP5y2DMfYju
wCma9Oti/5wrIRBxJi5VcHLh+ya9NR7/LyXmF5vUWup9px3razSO1rnwqYk54WDOotAKGxLvv6lD
iZ3hhZGTFRHxHPdPM3aqSTWwyPqWG5SbKinIobn653WI3tsueP2OYuPyHtCO5HcPqBNsthzqCpvo
WxeiIfsUZfxnkW1Nw/0SxeWC4A5sUlP/aa3dVqmrKBL+wsOmi8i1e0/o7qG5fv+fxalomefpq2v3
VUk+BznTFcLvbY1MdtcLfnkf/EpYAfSshNM3xdIH44Tcz8OrOGVnZitV6p5AGTNzKW/BnEwq/gLL
vaCcQ5sn6Vit3uXnWE0wUq3y6/nwiFMTX/Si8GxgkgszegTeFeSU42ajTDcZglQQf3IK+G6RfNSu
nH2aI92WtogzwE6Z93fLGtR4JYCWrfriVG/imzjxhfmU7RVBTgMpxaLVJGubLuLx+TRWj2nEclft
HDYegqC2hYjMfYenT34dB08UoYda2eYvMMAxyfcauWwuzy3mmhew7LEz/mX9vT8eP7f5UyINm68F
gmnjYAY38Rb7VjWDctIbBLTjT2gkv9LXhxXSV3aNuGj9DQK4RlnvVe+qSf0aT1RhB/+lngZU78SN
4lLjz0oItTMA+YKbetJaBpOepXp2WxHKRUjKtskwcKKoprJt7QkDtuzFcJBcN9r1SDsUPaPH4GEA
U/kXF71zF0Zw9BIoA+8Qnrb22Uh0CA1OLjSJms/7jgNFsEzHZe2RL8w58RHs6c6IwEC4eUedQnMS
PmHZWUmEcvFcXIt3AN8dF4+2Mg/bOCS/ujVT7vqpaximcRdAXHqCSgRkvlHeuYcKme5Si6ruohDQ
MyH8y2GZpNj5NAlOXpUKD0Qwx6m5KNUuQmayE0tDiyW4yrjsrWUjdpb3mESKT1SA1fiRYUrNOqCN
HTMFiG7Oau0qZx95CZklYNKXO4AcupmeOpRkM+MazoYZEUB6L0kcsp4OaR6rPbxpDGYUL/vT1Nm/
ylaJ53Fz8TwVdNAAqR0Dvt9dCxLJDeMwIT3AK8threTpv9E5KS3scfFq2cQHZV8oQkCWoa0yD6gu
AuYjMyukMS0/8CUtUIiCkL/YowFbTn6fnTwyNdNppkTcSDRuMgwX4/QknceRrVj1x3bpMbwXkbhf
fsbLxXdLvUiK0nDTuv4mw9RCok1iy8rRHjwpHOwxB3+bVtUY9U47YsiKIRUkYnI78qPJcFXtIGgm
yhZ5oqcvH0L7pMs/riTdGBuadKeIrvGQZHAryWY483Yee1Do69te6gv/g9eAa6YmUGmf8wUOX+3A
WkoQN1rdF1Vm/dO4hVkooC+k8/TyW1fT8VOXCljxzmt/V4+/efKO6/QOG7qf8nTj03DQ8vkkHXQD
lH9UOiOcxYk87lDFM1zguXiSsMqkJb8OUFwRxzfPGvjZOTyfO3nhsio+Zi9EIZWuL95BJ7DiVgQK
RHFWqZ583mxNknmtB8C7GPQ79jNmOkm8vfmgekTN+u5iYdZHMNIHmbF/2P0jLWSpoYSrstPgSq3R
7rRfWIkNSaOE/e3JyfdzxNnphKJ5TktFGRj/snB/ej0D57rbpDyVKbYSudiG4o5VFWrKUH7OqiJi
MW1hRlHkDyMORfQ5eXvKYJ1TF0SLe4YWCVHpC7s3V2bb5wtCaWhyby99P6FoXTzQe0fPgUzo2tJC
jc8SS/ugl4731ZE3zWPBu8Yoi2OacWx8ZfG4Mg6xQzlcsXrzar9HwVlaVKD03QElrSYd0pB73fSa
krbRpOiUP+ivai7y897Ujk6Z5SPk+8xeoFD5fKOmrr098twDxs58F3J8zhl/oU3uxFXNs0CrTx3S
2OlNZXDgDqoOd769HpKsWEL5kz/MC3CGV3b+bJNSHlcznkYAwzEQhtJ3rltkliN3au/M0xKcy2IS
KavQeLXNTrgK+0t1XDO+3H00azv0Ubotcaj5mLu+mMneoop0Xgnr5tUH5qitZo4NKUsaX7V/Fy8q
34ynVCsS0zTfEh30RG3T4pH4E6oZouohohq4ynN8LUGyeOIzx2QmGkChEN5AsskpCYk/+u6uAbFr
rcT/5mxTriHdLi5KSoN9AAKapFvzm4r165dU7QUY04M47mUKUXK3OFyigZjkmZ6mGSCWB2qt/+ca
WMGLX7STIHWjHlmZEEyBl8FHVopXPnum+CGyQf7Dn2Bs7/7DB1mghLXOPWnDtzjMRQ+Y3Xq5ZLCC
D9Vm5xw1Nifmb8uXmNxnJYHRhEW3n/rAovyl7pq8QrPMG1IJNo9PVBFMcgHWiTkU349hYhw/EPsD
TE2O+4xBVYJpWxMyDA4W7yf2GSJc/saV2dgCOXnbt/6QrdKJZ8u7ZbnbKTAOZ7Qh9T44MM9AhIl5
HZHhkEkOrSyHJp6PQr3H1C8i2fySMOWSFSPi0RhLDKE5kpYV/xb8V0AegU/uSA7hsDBa3DAT6dLm
9eL1BcVWwo4XUjb9UpObohS0wtJVl+GSQy/M8JAte9J4TsbfXxqT7U7Z+hMmPi0JBoyP5Bt5DgTm
tVxQPEmk3i69udYnyT1AmLWlP7hKHLhJYD0FUOzLj7l6ozIBriIHKNaUFKGZKjmgVqZqYbE4+0zR
ypM6OrEEKa1MYc93hP5jdWDK27d8Fc8QEI0njCmTzd9drjUiaYwP8YThbTYs4+S9ctbl6UMiVasN
cyS+i2wYjDS5fa09FqgtuhAVIf1jUyV4wA02TNGTI1gGLVhL24AjBGJxg3HlgrHm+S1PSI4uF+kV
/S8QOffJrFBzzVqXL2uc4/6vbeE6DYn9EhXX6a+mHngA/KjDmfRa49FfVj5XYTxNweHzvljpz/K8
3B2Q5KRipjtdYGA2yVGZpBSnqaKjCs/6RB8bCOazW7ruqHfMJWArMkGN+SifeelZv6QYz+dBtq3N
ONxGajOhzyL68uGm24KTxN4Uh/18mfuXHalUD1kjLgnZwJkfKeLpLS7ALWakRtRZ17sQ/Lg1CbPp
pqD+lLIJGlu3rdV571t0o/ErfiwYFdUWbdt1H+6/oS1Yvg/e3d4M16EsQwuK5tfuWcmIOqELalTi
iZoXKFQIVrpowTO9UfPGQrd5/0iY/Vnog3pN5hqSA9rkGHMn9DsCp2bfGnLQAVd71N7jZraavoMZ
Fu9mxacBK5A6qLTQ8gHrMuNoAHrLhWe+UwWEzW5YPRCBHuBz6Rb1bV57LCOs2L9tGiCruKZ+2PLK
ye72s+SBUUvenT7nqmlKpeQBym5q6CocANirsb5HBJvnnMlApInaXFukz1Ge6mDFfnRPW9AUt7hA
mge8dOd5nFtrTvyQC4cH1AVOSs65KH6zIIyFGCXGK7cyCJg4M0gwztaAh8x9YuyUGD209cHwTHZ6
azwAMa5Z6DTbg/bvfzB1UtY5M1fUCFoSRNID+GKqa2G0mP01pCHQpvqpTMVwMZvvBIAEP3Fibhqt
tfybV49bJvZy09YxtbpxGL2ZTBcfEgRN61g8hh9/tPOVgGmuAiAv4IRlhPaxsXUGr9rATbzlUwxT
qFjHcq/sgguriN8tsTUIz9f4HCBAuImauGLIewk5p/Ht+WQP/pQQnUkX+Moe5NPL1r/CZ5Wy+J8x
zL4KBg562vH/8l58H61hgaOu8q7J0HfCk0BcU9wNyoR2iKptsT3yTe5dA2kkm6O9DBaq9xSRwaJv
sczs8X0mW2UlD8+QMT2gKY3CPl2WYX61I4OJn8ZC81GDh6alm65GO4dTcvF1h/xrj77s4VxFw8pf
hG0nKbRpX2X0wQb24j4NzmZOj711ndzqIRbFDhVdFdP/oWLQjsxHI+COcOplj5il2dpUBsaaesyy
AOPmLn9E41pgJTHGVjcjqmsX3ncEfD/7KY2YrSOUYED4KVkqbqQnLKhmQND8wQGrocukBRzj4/tb
gDSQmhBp+L9rf6A17g5slNizgRGZXNLyCJY45hCg8z0Pc2qKPhvALsefB3ZwbGwAZ6teArm37Dni
1UG+fKSqHAZ69/+PhZ4+CUJioeD4Ty1e+HDsvZ+NMcdApvwGjlPQ3T+GaEslcJAQJWbaG43k8BTi
MOewsqGpbnLrTZFEt0Iymo2M6bi5oDVceBuxEHGbs6+wSq6PnWuPggm861OFnsjjXB4b/lpd8jwR
42Y4J72HKwKI1+RlHAHL/smbPGoSohrXqjKVsi/w0i396XUt0McVoLtKPVWIoOSMWIvl4Y4QLb8n
rXytApZV6lGRxUzEz0FqfKRuixsvHuhsi0s56jf048T1E185tXyMfHhIAK2sf861YkxXnQTAK9OB
ru7kWJd2+tWfNDKTTmDsVjhDElgskw9E9QXDo5BqY0Dbk4MZez6kNfYfGrT92KEtaU1ACl+hWVg4
r2nRRQNgeHuGkZNaLswrFRwGY5MMDNpAicIrwhynt1WxMLdTkZul1sR/DvAr3XdMIJ3yLF9EbNCR
ls7fYdf0YeBdMBjoenIzZv9RtsQcLEwBAuj07kHPyuS28jeVFHtJpApIzycqtwINpY52HP43bj1H
7Xzcv5gcfmjD08Z9vMbPQYpiF+kUzg53iqAS6PR42FpKGfAkD3L17rq444zkwmrLSWz/oW2qjECa
m0bnv6ADmQrQYZAd94pBusjCBT3LD9edH1Xpwrvzk46OrM9tH/5XB/25gUOyFLiMlMkPC4w0PQdf
CwfW4ffLCaZQQPAyHPRXsn6AMraAkMGmPaYm0i/ZLJOW1dDFO48KUWtwiZgxo8WHOHIh4FzMmVTU
r3fn8FyhqZ91clueyZyPysV3luryU9SAVCgt6OkRKXvXD3sKpw/A533SeSdjTh1MDjFWDON9p/s2
lzhP9aDy27RoDMntdpaKseIHKdfr3G+ioXluzthI0tYHwEu0ZOIVJVfNm7vj1KvHDczgT1+bwg25
vvhmJw6kj+OPuyFZYk7bNWUvhF55Nw3puPGt0yWfEZvihDpCWlUvSRhI/zr6M8Xi8KnOotf0wRpE
iGfkT0P9f/eB9PAjRnUq2HvCyZ6qt7w3eYvPeXj7ipYLO8jwbbH+vaWmGzjrxms16fTZsEwjf6ze
QHCOuNM6cw3O9pzvZJHeAlEm+GxyVLes8qkxlbv73HGtCzXP4cyfWSEL6tttxMWFC95UWSGL4sc6
2goyr2Xz10JW3wwWDlI/8Z/3+h7vJ2/BQUKt6l7oOMWfYMNcJce0f25/B7P34ldGj940UARktoxr
mSwgN9lncO4pLAWLzZXqsYUEiL3I+K49KiL0UC4tCgqp/vsxRrVz0aWfFGAznkZc4mcgBSuJDybL
jfAFAu7uczyoXvFM4j7rIGuJoya5HvH9lam03SpS78p0jS8Kf1hE4pRqfmj4gyrva4P1MoJIqdMa
CeLuglPas2WnO1SD8AcdaHzvvfkRpHpDOdL2SF/6uOf0AGMmwJ4aE3bOY/q+Mb0+0YLohrZ0vPLg
/cJmlUEtd3f2KQD86tNbiY0IyWtVlpDtqgEfvlufmdLT9JvU4T/MIzbP/YWs1cZ/BOEz5h29OpRx
qkZi3Nyt0PcllVWsqQwFmXUIXR68hTppcauRNbUEQVgB3sneYc6Rz8TRF4pEXWDFVw3+o6iTM08t
VuLAyQyfIuOKwAIkLU84bodsnvP4kfwBDsfmwQlaHCrK8g/X8mpl01CN99lRDqBlqQXyv05dBf1d
O7Ze3Z2VN6NVKJvUxBFOfqvtgmrhYDndtq8Mz/p0SuZY+YxD1rfMr4kzYwYeCMoNqE5fpAdWZP5e
DGLHqfbe2rMfjmHGRRw7VYdLwyffM55lTU8l8R/pdiiQROCem0G+2WPkXpuijusGW5SZqVRflK3/
7u0YZyzAPt/CCd28nUKLSUewsA3inXLiHvQ4/j657DRf0FdWF6N5Txc9Ge/OVwvApAKaJ7b31V64
VO6Z8z2HOW/Iw8ldJFIPoXxFK1t8EProkk+R4grHbD63Pv7+SXThZknNPSzr+xHLEN2MMrMiQIl0
w+cOS4oe9+T93pg7getufy3zl333bhk1TDefB9JldhzBKM7rpANRbgjz815hE3drweF+odn1WKwh
vvxwdMgdkM0fFhBG23MIHE13yMw7aRhLJA6v8SDxONhOqWkeg+Gc/bJp9bQSxlg4+tVtJ4NvZ+M+
u8TFdgCp34+PFrlqgyTqcJW95YxzyAIcGbGD0ONlTPaj8mCGZICaJ3EIkzkk6HAJjAMSXEqkvzlQ
2lyANLpptcaxmJZeP3RHrXbv0GOS2IDM5NOlWa2Or8EnWBwQceVj99An97GCmo4x3C4/ACva6OmX
L5TVLhxhnL80L0Y0o/vvV4XgsA8fq1Fs6uAcHBObWndYNX2tXvLnVqw65f9CUUbpAVh3vu54TZl6
Nc8MBdIBPR5eSORKrDMrOaMbqrS+ckud4aNf+Tu80WV6IjFn9s1bvGJ4X3wcqWbYwbFhcAeC6e+6
ubSWjBd83ikd7zlZnJS4eQZaK5MoXFDsvEeP2j4vTUq5v4cHqe4r76p2cDLiolqwKU5m5AfafjYm
d7CKR6cNu44oS+DpKeyxfc7ctGqokAzVKU15LH+kSmybBUTV3Dm47uca1kjxVA6kN5xBFgITxuW+
G0sBUnN0ayItpvZsADnd+5mMDAws39SJ+60k2NdjXCO2to50mCdPd+apLib0P6E/wyIDKsuogbmB
x1j3Y0QFd6TXwuLEgD3LbPd80lAwSxUp8qZM/59RSCMx7+1H/xy5kRi9/dyRLtBm0SxNmc9PujKu
NH5PQ0tBUwvZU1Fa5LRMVPf272VO7Sevrirucna4vKDvH8Vcvcp7aDNgRCEp6Rr03TuVsAHAliMP
SxcF+WGyl9AzNjMsFZv/JxZlJnARNaxP2uLULlLfe9hoXOODg6wbELm4dXhp/S733x88NRojPpBi
HhhILIuBKTG7hUE6wH3DiW1ES5849UZkTrq+mzIloTwkbpxRljhqA0x725VyIg/eaprk8A4feNYB
hTu0kEM/h5jfEsISgMEYB7u8k8vyCDJkPvdMepbZyN/nv0uKb2+BCIdyOgoY05k57ijuaaJa9TD7
ebXfUq5jO88kLOQzz9ENoCi7mwE9y2u8WPZ3hyCgLsXzMb2iHvWm92DRcwvRYLg5bB7xV6KRxH1Q
fTbhbw5BALk7c5U2ZW4SiF7SUisLpHqdDFS7iooeeIQPDfWXQJ16Ffr3X+Or/q4jAtZ2Ws+I6e53
1lBOBnwplzOredmmP5QYBPifmxloUEIL3iBxl5HaJKLWWdDDzEeZFT3DA56q2dcjkTgwzQJkPCFb
WU8Fx9kUNE2EldN5KC7gi0CPxzNHAESL1olNgjOeD87iUKO2gtDxVqJAv7QIrmBFMrKMP1176jaV
lXiAS/YoNdL0N6o908hfrtbrKAu1SI38uz7o97BrI6pmtkg22RKf3GPcZO4MWXvI8DGjLQ/HuuWG
dUFFfpjOyLOlptmxyveYczA62jAxADtJrqaJ6GTBmhqhU4IwCPt5bL+Wz1MvLgJXh43KFLv1xfrQ
fmsxUODWilsbX73hQbk0CenuOWNZBgkEVHpNhNwL/SyqrX2ALZ3FKOVJXzCpz8hfSB6ffNnyByzL
whpyYO5AgyWDY8qht+N43HboH21qYbGxOXZ2oirTfEiytdwq0VTE/YWMrZlqP9PhV6UEBKwnBw/f
8vIXPiQ9zBspugThlNpXgxgfZh+GK4xGHw94JvB0y4d10avsDeZB3LDRus915L+mfabIQdmBDYrE
evQz83C6quzLwwK72qiNbTJG7YwrtjcMljnijuIUDp5wryyzy8p+yzhwMse3s1uz/i9cmh7hCpWF
S1awUrRqMRFbrBkk3WwfS+HWElXGdsfAYtzGN+hXtAZRh+aeWAQDHvonV5QakczZs+WQDsZQf+Ml
29CA0FGE3JzVgBZOG2fm7ejkx1tGp5cAdizbqnpSTPQbp1+qSsDKz01LwDmQ9uIH9ohReAdpYV+R
kPekfAcVD2q9L46ppeuQ1oZKwB2BZwTD19Cys1wYdkXoWRjxUcWbEIDfGQte68Zo/Jd2hSW8uP7l
3D751Jy3WfgU3I4G61ShC53aPsQc85qqBsNaLemIWimDvX9z6AAJl4wgyrLJz4hlRvWbWLcls3T1
lbNlzWzXiYiFp9o+CB6tQQKombv0idYUjxAyDlfWDDdEh2y+IGxMLPHKYPLPkQYl8BhDD0hH6aK4
FyIyDJ52QPOQhi/lNOF+M1hjMgEmyzv189A5xdYGfi5gWrsEO/oUqWf66twr4/XKs2clXnihrhUv
7KWT805u4PRWZRCiAOUBByWlCMSWZLZZh/F/YmiAF3xpAvOpp4d9UNWk6CoAV0cXlVrYLqtVZFaJ
SZUE20raZi1oTjCXUmZP3+g9P3/JWiq0r21ZQ2uezrVe5s5APRfb4q4Y/zU6qtbOUqVB7FfGNo9q
BEie5crMDF/fyELbLwKmq9WRUcWytTXPZag8QYOR0JwOfE4CrVzS9eiK3AiAhP6zzNU4i7198uaw
ECi64SSilUGk7oK2bLgetulWEZmXqkMV8QmljNfMdjLyhatjPtq2GYpmLhq2xS/+nIw1MjoNNnVJ
xjV5dZrnwXBaT6Hopx94xs8hbYxHyZMN0V7X7xmLvrS/OLWy5tpMYZ1q26JRe7H/OlNLhYMda2QW
56pdS8ysfmkpb5lQxMUvt7FZov7j22PU3o8HObrg5LtIdC6WDzYdxT3VxJSfcjrOSluPF9lVQ8k3
knzadrzITfJ6m0jGulWhehTo05QWBFzZP7Ah1aG2asnE8LA8Ag/4e0PCpDt/eXDfA1RGKDI//TmJ
H9GSCZsekN9MwNSza35FpIME6M0PVtc73Y2q1mjh5zRxX1A5XbhdIAarZ5EUG67EhbMnM4S5gmqv
6SHLf08Q+9AamNWFTDgcGVixK5IAs3B/dPvCvWH8HbXXpbnuzo6ndH2f651QM68imka1K/uP4ZoI
8tijzYWzrgbT5q9QLmCQ2O7i99x5enhJmdsvmwpHdAv7GY6WNMHtrWh7wDS1lBGnZxHFeSU+bW5D
qs3KJtcZZWOp228t20lJZRSATuK66453kg0F/aSQx3+91AOPr1Ys0l9HgO1FICOi1t2Mfy0DxnIt
uzMVqcD3trdJCLpKqzBuARirw6lHSs7KZlPUexftLR8vBvEjKWKtD5n/t/oB7c7beBN9fj3vLq5U
4dB0npujz9iVdm7aqJCQicU/4oBv5ksTRlkfo/RJno0Wfs+5z6f+AtAmmqHw44SnhLGc/c9O1JoD
zx6HF6e6hTssnZaQWA1QeZBeK7tzpNk1Swl/Nwj7gtbSBTIrthDapYQ+RT+Uh0cp8067vK9VIPzv
yLDvsdA/Y6QDlES+Xg5mrZvYUu6HDJhv26Zewya846N/Ooxp6fdctaXJ0DcDWWgghsEzoj9MRGEH
wd1Xmm6eQI6h98oC8ragJx+rQUYQ5QAsU7D551DlEQ0YBalaNcRdhvPqnXAnkQYPHOubEhOhjeH2
cX4gu+hsWaAmPQl1vpH2qHV6qvnvTFzD/0tSYrVLJMBFoX+Q8YAqEue/v8b1qG3Xj6vQzEA2LCZ7
wZ/yBZc5f1UJpvB4uW31d20zoWw74/VKtgsMqhAZ9vpZhdkXlJXxNl/6XixrMXQEaoFCsHLUw2o3
X3l7nu+W+Dat96fjxRxSoPoOOKYiyrWNOOQpGSwse1nX2NabiJB66xwWcf9TV2+BvLQLPdNHM2wM
+YWXl60grFflrFo5mPTArlPcRqyFiapgqHT6JoyNG9VWuKUNIR4nbUGly3lVnrPuJX0xBU7ee16Q
4hofwI0VBVVJvPVmoWGIUqgKFJE9vGi9jL+DkQy6p2rh/qSlSEqNbo1u7vT0TAMQWaodgKCNAZVW
wXu93qo48cVTQlw5lkBhG7FiuvCYI9WGufJ95f6lyMnZvV5scHiN/VOj44Lq5cKHzouHlLUdiJSD
88bqSFvntzsYJ2BW4tPzrVG85rg4Jgez6nvm2tjRZqeWOx7O33fzHxpoRYiDo5ZtjpP69L3o3wIC
qU7RfGdtOIJI5yDjm7W5wyLuJj85Yz8QNxjKqd+JZErL6OD2Ps6eFHtVK5weXHyF8g4AOv90zRYP
z8s9tznniMH0d3qzmElhq/xTJeJQNEdY1D+RX0vrtWk4wwT3GvRjzoMDtoaW1/q8O9z+n00QrCK2
4w7w9S8+QrVSyHqmRxgBKJIGMPZK4jx0dwuMuEjPsr/L80BCUroCvxl+IKO40yMinFFIP9ZKBm6T
E3wxy2Z/BHAN4W/UBP50F/LjGIvCWm6SNBq12HvhRTCCkT3GuMCCKQdBqYzNk2jX6ALd/6SP/v+4
UL/WXxMRXz57bEL27o5hDQjQn7R325zkt+wXgfGjt53hnU8MNfV7oDQCz5r/A0jf5r0bFYFrlvTc
tgkFUwrjWqWgkfitF/ctbTAON7mQ4kyHr21H4N8Q/lGQPU2vZVBVfx3P5OhIvSs/XpU/xeQ2gAwn
YKYzcRm/N1D1nzZsfmC5KDdF1BZARhSrUvceNxFKcu5gDIv+ldZRqldXWY7NzFJgD8xYzmaYvW1A
4WvpaLs9T4k5RQXvWNwtPbclnjpjedV9fHDnDN5rgwzhjehpg4y13beUlsDL1ff3sbtK5Bw9DlDm
3+AtcmR/N+LpO3MxH5DJHg6QaAkXIUKyyEbrwkrxjfpj5CEg6nPrNwkx27hEZIF8tqjdjQx+/Y44
dBy8iu5dENZW9qcvw+PY1VX2f+WtkdsvZV85VTebZmj/aJTEGyHdDx4TeiRQE6ODilA6T2m+7cSf
6Q29ciJl4ePJDBWConHESxoAUkZff9do4ayhdO9/ZEDlSj7gPmhwK5grthep/8PmkH7Ah+0VyAUe
LwupvFfJF4Ops5Ua8HIzY3hY+85/upnypKbYNzVuKdXWc+NKTNBAK3ck00SDBZM6s+qQVI/UiKlU
jNG0+Sl948P5PiV8MlTymEM9MWNJoyknmxNE0wNQZnHuJOsY91OqhgDA83E/wrpetP0RKSQiez4y
3bXj4t9m6Wk1cfKZ30f7XC4EnVi1WjKFOkerqQjFhL8GbLgu27i0M20TcE5wXFSNJR8vD6UlUUgI
SbTfaB8d8g1W0vnMuN8BM7pMZ1GA1mgM0zr3FWZUH6iIZeHbF4+Hi4IK+S+zn0xtGSJFwmdPLkOE
Stg2uoMEqrZ//2IbXqlQEAPNp3xl9QrDWOizeSoBthSf1uLCWn5ZfTkv+RvWZ6bmSA+yZgIY5uRs
KgnFpcCQgvJesUHyG3oUMR1UGFgbPZXs6lPLo3EE2QWfY+zfIByC76FrhEvUBR0oMLwOby1bpi+R
namIJSalEu/HYumklf3RdjnJjvvpAhFb5fQUAQH7ybRViUwbpWzZLj5oKYrm9krYrgzT7QmJ8Idr
tIp4piFGunH5joVv1yBsXzOSw380feeotNOHjncdBwnrXJl5SADpEFwjGjRy3Pkkbgw1UKLOFzV8
kYR0aGoScqWSYzqkU7qSs0kL/nxajXyPtI3qyhKDrTMz6XnAJKbOflgCMAvX3QMNik536tj5gIIK
aRm1BDuF2x4OLsz9CdZMTuJqGw92DnHCLNjsbv31nkpBrPv8SBxkNuXxXMi8UTFAn7g/jnVj6xcq
ANnioRkDqJj2FjChxcI42ZEulS6xGifxEJhFAYtETk3Uwplbu2tCDFuxK6nJxbQd+Z3ZXRBkfXC4
Y5EPsrHUjSigW8HaAAJVH0dbgpHc7jWYQ3XdrmTfNW8jiGaj2o2Amy/AJt+5HWd2CE7YfE6+a5eb
hWAOr8GTE2c7lDu4zgGI48OOUVZioVvGneXNAPpBt6KNXczGjdU0x4WvLaBxyk8aJn58adAWrQbq
L47zxYeN0eEs0jp/3hl4ZMjSKlB8Wyjh6T1Dv2pl5Zkx1Gl3gRi+EQk51skIMN4+t2BnoUOb/bzF
2FfYEvBVLdE43ILbS8PZTwtUF3niv+Ef5h1xtzdYIs2uVHhQsdTPFCZGJ9wwP6k77ZjdG75FGYSP
iKqyIGzb//jrg1OXdUxny2CaRqxULKzszfSNRgKxaYDC3mNIA4BhEhqbdA+QGEO4XhbnU3+05uRv
dAvsyDMvpts0DU6mym4jqCACkWptnL5z8gpWMvV34pLxtFGOl75Ot5R1VaCAPRT6LWEEX7ZidLLi
//FGhO18FpwjH4s4AR71oTSp3PUFQXAwFpsJmPdaN0iBTgkkPuUucTDBtcp8uQEYwHf38HoBdUJR
OdrDCnjLNdZxxSEyFR0rx3WHiaC3FawPaA5zbA3MpEwGEw3DVVDSFN1aLPk7kKEnIcX0B0NAalVG
wYHj09t3vHplFjIp/vEtemLhqL8tKoAnSZOSqO1CgYcqnokZTT5+ue9nGLlWMQgqEKaPd2ARu6Sg
2MItxfvgEbYwdb3Z8cMQPWkhiNFJxBcMKB2ctenP4JZLpaZvfNyOMc8J3qnu6BOmNKet2kbFt1OI
9xo+IiLNh3f2D9+KhwKMRNnEgXqVitqeRhtYktgc8yNTPQe38drKZycJOj2Vqy4gGP2zhd7ckA8u
5F44aE8GneqmLt3eNz2zKSc+gE2A7VesjLy3hqa8LE0zW+h299kESvFEyzJVq+lbgPJ1hAMAr/Nj
YKs+DK6xfA0nd7fyv/45iehXhjIH5v88yGf/CEm4eNf0G/BGsirwAGlO3Wu26oda5CEewQIpLx0Z
k01TLMRBlLN1slq6Srw9/acJp34aKvlSLhM5m6+C2tLUTSQlifJ7bjCnB++NOWAAZrJeCBeLAldh
ZkMw7MP3gBonhGCSZTLRP8cvP/9AxUlffv6b8H9qi9m0hhWsiezZ3210HBJk9NxRFmpvMGD6ZOJH
lJKBfSEWldKXIU6O9kMy1yjAZy8h7fvhvdUriH8BmECrOG7nR5CU6+zC2jYRxkhkM+ScbKKburhf
AaPjC8eThAvJTuc7CgxHlAohbIbE6CydJ8x3XMvBBkBfkH+uJFCvOOGbbPVryqBWmNPIggP1mmP0
bDB59wjlL+3rDN5YZ7qhYGaQY4ByOxnAlTDOBzZ+ucX21ghVKaRWtK1CJROvLT8GSub0aMhQZSbq
H8Ysapm8/ETIpXIMVOygtm80TjeIxH8fBWSYTAf1YpQzZ2s2EY03UdEehJR4LB65sGwLhUSH0b63
PwT4gsHUUXvEcQm3jq+T67npLgjjwzKQi98wO2iO3IN1H6N9BCFSDycZVB9sY6IBiFyLpMUYNQEF
J4srlhfTsZ/Aaui6N3SdtEkRRW1HTD+sfd8iFVnoo9hTh3TcuQ7ZX5qWIyYId/7d2Y0TMfLOMs15
DTjSmZg7cJtbanM9+U3Rm5a2fyCasIlEaVpKwWpBKdBOqJ9l7bz+H4JU7AaMWtlnUaSkD9ajzVmS
S/I6tUaNv4ZAa7n2iHeV/iA5TRtRvAdH6vupR+tb1yUhL7c2NApE7cK1eoduVBzOyydRwWTr2Xkm
2RY6RAvD/ai0VQdgirdrCe0ajeYBlAHgVGAUlNeMNXP6IcltJcu7oBlHGLjH8fZ3hHLt6c/w2uyN
PXQir2E5iLApv6QDcyLxgIr6FIwHYMcak1MGXRX77tktiOhly8HWd4P6aMfbJ2E6qD3BJVFvcbAS
6yn9wshz75QrLEtYagu2hbgTzgDBRbYPdDU9BPYPCdz9Vp14Ovqpj9C3/deoDxQegBOe1R8/1RID
ppwOdZcIHz/Baqdxf/dm37rapHIMFwL40YllTmj2GqKUe2Yf9MYh696u47kI5VuU9doWV2JjSGZO
AtL4Umwjv72iG69wHaDcOEGMDf1/X1qzNn2BmdN215UHXlTx59Sksu9PlfU8jHsBKPYKdj2wVUAC
OrC3n56b0zHhx0mW5bEKa4LGmiKk5cobbbSS/kgei8CyuvBvkPWChvqvlkG3kgXzLFunGm8ZBppE
B+o6CdLzC3Z1PMFxe+3fJ4qDa2F9EL0OhcDftZdOFmx2CTYP1RiqdDNO9LmMOFNBaKVjOpHWTIwC
s1gktIh1BXIoHcnLq9yrJgUxPn1xcFAMRZzKDaogqS4WhxGTA0VciqstSpDSvF8hcbHJVJ1/v01V
Z3gGw7EG6NcYrGfJQ3iP6FB9T6563qgc/qDkK7oxENFNbeKPPkPMghXd9cv/yK5660Jl7cOFlfYc
eLXbOCP+GNMUV4e3Mo1vANNPZxc/ymyerhhzffbvpKpufXNzA6fyk/ZtWyAM+oQ+5PaLK58hyDDR
bMEL/mHZy6IoTSfhSMBmHAT+locByTUdvvqpbTeHHCQhCc/ShH9EixwLYFwiWEyQNCODIPlE0pAB
sHjGgqMFovIY7sP+fW/GP5lN4Qt0aEdS3GK9F1yq7cvcMhBMUzaENXQjW06mY4fSqXMsj/zZ3Z7t
A6DUg3uf379bXKQk3L4o2YBpVvU3GhgSYsG/RrPfAxqvdR6LMv81tWP+8ZreKsaV/FJ5gtMGMv+P
yqsQWLIQVAsx2yEOtcunehcQUaWTvbV2vRfglgEQ5tpHmsnNGoCggbFivM69Vob+C1N1fSkyhRKA
7N+KHJgMRl/aj9X8A2ZcGN37pcM0esjU8DCWcfJurSzPtweE5pu24b/WX3c7Z07e2wXGP1G7bX1r
nVExxN7g4dWx8AJKiuIh9UXsoaA91yzIX3WWkx5lDN0U+yeGiD/0Wa9cQUv48H7uI3KPT94qHh1D
gI3UtsTL6uvaEWRgGwZid5bimNi2h35rhdjFAditFTqttQrG02V/luOoYlLjHIx/ndwV4iAf8Dps
5xWQv9ktgUoTabHFx5FLBZswW0afNHbP8uIB1c9p2uf12tWpKfUr4yfxTno7tnlD9vShSE9GvKDW
PfJKn7/6te0MtsvBBbgW54EwKfJyaq5VjM+x+F1GNH3CFYI12fUpFRPPG3yhJOCTp2gw9FS1GgPT
rB3qq1cEdtBd3Yersr4XOv+H6Eq3cIcZxDesQXZVpCDeMBzpr4iIOEgY4fmMoGEViowjGktyl3JI
VssFW25JutGEYugQtdl80W9wkD3HVu7iyUi1Ajhf2cJxxWLYfp09bAgQ1NEtwrAqSIrxtIO6vXkm
B6rJafxhno1Wqp6RdiBlfyAXq91WZdcxIyE3IBtV+VZtay4sDnNhCpVpzi8x8oagTnBJpIlDoIBn
p9tQerMGTOQOeWxvy7uFzaLbatHtbgoxOIc8w5vcI4tiEXgC6923PGRYFRjt05NC5kYdc68GT3kJ
I0Xg2DyBOPj8JonP2fI1om9sw0Mbpvr6UFYe2Bi1IwQulXtwZBR2pyhAFuWdMA3qzDei6JUYRaPY
6130SGC+S7/o3kKn61n83wHDWLYs5KBuLFy6lnW8tBnKODIdL2CeV3gNEnnK4LH6pag/90XG8p7A
QgKHRMyPnFq6w0qQKC8aem7beuux1cDrxvW3UGZcXt2xesoXHKcLeqbqShfIAFEW9VIRJXE9JiJu
9aTQbbgfmxXEfwpgl0fqwdji2ye+zmhM5zMCxkzACN9HXJHirDaQd9RnrHaS5kX2kFNSIH9pIacO
3j6/JxN3sxDHLrTL6zm1tiI51KhVskFAp2OXBiUajaw1tnRMBUo7f30IVi9Ind+Oe9n+PK4MU+iA
v4c+tlraLG7UPZ+sc8K8r96zgWe7Kk/tphQGy0yJ5avWujNvXTAaEYluA5D0SvdK59256gsdpWf7
MjpTi3mdu+xmWXf0FFDHz0b4PlCWza/oeFwtJWhzuXrFLqYZV4zIwwPqmldooCpKmJ6LRF4aOCk0
rFzbkp1+MfKJ4XmhBE5ddfJkEnaytb/lCFmkjTbW6wgH0ToWK91FUNt8/ZgYpSCPE58FNy2siToC
43TOgCU/yJVXB38cy72xGFXnOEFmVpIpb6xDqBzMYALwe7MCNrCCcQ9AJgEqFZoDPS0GDwOjn7cA
0gn1CzNa/orqA/mumMlliMddsWGpD/iiUi7NGX6gtw1j1w2hgK7bAucNGm9aoptHNc81p3jLCZ7x
D5fUqe8LDclHBI66dcBCKsYFpFBt0d+PRaVNTEGDxxrDYKetie/Dc1LAsoFGVGmDeEYsvQ5+4iui
fAakh5K0buFC49JQEtParpU0qxDkn7+KQseyl2wmv/Ck7gJZxlCOalS40CDXmwcCZFoCUfmndSIx
cQvgY6lFYZBl0eRNKH56YrAQZVbafgYeWsL2MVv2DucAWjXiyWPRlIRcRuoLvD1jv1KcMj+xHqT8
3jeijbCCqEo1HwR8YVCKGpHJee4DpPSZRlMCJmI9eG2GHovQ6L8Caq6zNFlvmzNTwjg4C1fxM3FG
49ZYtsHijaQ+JZXEzsQJsWkG1+PEvwmuLIw9OolbRyOfVad4A3YRq8qU0HIionlRhuoa2sgM7Anw
+24GKLo3A8tM1ky2Eu4VitpfXZuq4O6jWqi/miL3iET7h5g0MAaV+E2qtENhVckiRPRFWqNz0Va2
8Ma4+QNk+OF+cv8gei/WeLG0DYERxBBsHRkBCAYw2wCLPYAxwUktzTXV2H5xtCcjGnCpNpOmQlMw
V1FCsjQv6rVDXd4AZ/sHP/tPz244pgRPv5nJmNFZGZk6mELPK1YqpeRLgc+9Bmjh5Wjyi4j+mLRJ
vC2FrrPxDS7LjCWaFT6H/M0SMB8TLaLXB5UIQ5Pdg7d6StKVasOUlXUaD+EG804wrz05OKLQYOuE
eS8rRpawjb8xWraGZ13lrXf+WP+FCSFGsU7bTXtPExf3yxZxm9GGpwwpVWhi5OL/zbws3WlVcy83
lWpg2ge3A7yTwrX8i6BSp0VJpHfCE+t8XLpjZBhW92UQftBTTVFLAVYC6ejR7V2hiffPJSEOh562
1Dp2jSJboeLULFy9OXauF/wwkm86cdUZdAiJbHp0TRtbrpLWiRsSH3Q3eKIZqm8JwunLD/ZNLvBc
SWJ4klO8fj9uV2tpUhdORsBNUg/cH+3BH34K/ZGGz9raPD1CjmN7OfvI+YIdzFDzLA4sBtbBPV/J
JL4M4xDVKqOz4WT65CFJfiuT+8oS0SQHqfAMBAxFMCbh+LIaL5jAITFa5CxSUFuXlhzFfI8U7eGT
tZ5djQHHdDBNUwY8C0KpTl/N+u4g2hiJi7LjauZtmm6xoyil3Zt5e0mzq5b8TWyAd3R9KxHfQzA3
FG+Hl1DoRva1jLnuhtmx3h3oLqoEaxLVdt15szFjcNLurPfNCjDPk1Mcu200HB2RNBX8o3SJi9dN
QaHUbCnRLmi6MpM7s0VUU5AhNvuLVvosj8Mb78j4lIEOsbWy62zmsHIi5zXSa+S46v5LOviMXymS
OqSNMknQK90IaHKJhLLav/IcdJqXpDqFD4JQ6W/4ppHe1dGMyePkbBNXSQDrzpZEJK4UvEy5IwLs
r4zTo0IkBKGlqD+Wia/G7bC2wS2w6ijgDg3dcmOOCvt2s2NfFg4pHkWMF+j5TuK57KnSL/orMVpr
o5WFz06RGRsb3oJijeJah6Wxp6hbZFbiOfy7vacgNeXeNm1azRH8hQsaiZ0qByE3lHS3pLobVGby
gHAejlSYZHOXyBLs4XsgVzsiqX1mFgCTkd0nCDxBU39bwftVPZdRvuABSW4paeyEb/qRli6GrqMH
Xi/3QiPe8X5yBqVIgGWmrXcLb0JbT7VsQ4VP6szhtq7UUy4wm2CKsVzBqSIfbvG6Xp2CFi/qUWkC
1EatarcAnLrnQgKzPblwkI5ovgFaQod+BpMEGUkSURYwZ+hyRDXftescqGn1NFasPABOASzdPk5r
ORZRvtLvfpc4RJWoSOq2XJ1Cpdu6u3UHPkDK2ArCHRl+HfhLP8H9eO8RXHZxnEnvRTP1Pc26beSI
4bYYe8VXMqVBKJiz4aWu3ICMaOSewqetnddkXrsBRAQK/qVAHp0Ppzb7R7sjUGV2Aw2CadG/yDh6
66KQF9f8S+5V8s9bTqB/K3uw9giW3tFvYJyJvKF+gHl0wzfzo6HINW9nMYlv4xGn9LOVMwDFb69g
wE3EZYg/+kVcyrJwUi0XP0fPIPdxSJb4hs+ctcP+uuJOydgK3HOovN27ZyGn7pnrq7tvLJ7C+799
NsUyJiTXZdqoZXTQOT7iOX7aqKiL2rB/QC2dkY/gS627SV0edSPedRujSYgJYg9lHAPwCEO94Z0t
9ileaVcZjuB0qiUNsB6xeAtvQF09E4xmXqVYU91dh26u85z4SdMNqEZeNf/DxEbtn0/xY4nZ4AoL
xGOs46sEZ/IL4e2LbIf+GrNe+kYyndk0rM1OXjzAMFq/E6lZa4W2ne9KvXSKG9UMxgREfLWAxl+n
5HOgDML/qu8z/9Qg5EM1UrXpk25llr6K7Ei4CtJppWJwrA0oTvTnAL/mmArR7gK6j6SobsvLF5v4
TJRVk06rtAGnqGp90vBTqyPAeITQMYOAPNvj1ryo5DK/5wZiEUG1pDhUJ97CcOtR1+fk2mtzdB91
3WY5Z/M0D6zWtEkn1QO2E+InvJrGo/DYAtV4wfyf1OXh14gGhULxbMvL56xG9QuNYvwB+EcMjSMH
qqMFZmxNBhV3wiITeGGZz/6oVtaqQox0FTsuopEr4h/hziMEgJ63vWGSVzp/mLaqU130ltfj/lON
n58ZhYsx70SrCSLvEAOWpwwrXakIC+8ip9NEnEoWLxSRwUitiwY4NjmqKO0nkvNrU9evw9GZMw4i
FO3kQCNSoD8PjoRxs1xMPfNE0a6RAzz4vOv+OPPCfHydoAP22WRi8DnWhkj+/zEYvPxbKFRXvk1T
UdkiMHlHvPkq5cV+p+pLqYT8NVUVdvFSL/KaaQzN7vsqC5OGVVbvdHmKQwawI7MFXVZfDkuZ5FDj
eW3nO8NHRwNJYjvDnjzrWXHt+qRWvhJK/xJ+VLqPbXqReA1RsVbMMB31tovJp2pcltfobrqzRkaa
rD/iCPZGVGePQGYpmZmA4pnr35bF0ALqxSOLHnfnGJbAPFH/xl1zfFKFzH+pNuqPhCLpZfEJAx+o
JVTtkl4drOJvGsiKr6tnocH/LP4Pz71itcuRks4/p06o54/+X2q7RNVTzdanuR8STZahv9IIoyCv
QLPt9FHuuvjR6bwdGfSDNXqMgtz2bCBLJpMFgVwt2JdLAs0OmqEJ1YQXQPqpm80VLIC9d8N9jEt/
cELa5tg/zan//CgyVdDdiVvqr5Sc0dJrwm8czyHBajzJ9IoU4ClHBHGT/IRXR9dsISRmDJdP69Ln
bs7Xe6zhkONPS8iGTKzNJUQEOjOj5Nm+3zUniuH/Nh1K1ewZrdgB2yTjHh7cLPLwYfGIBGEMH0nD
/EOgT7uJrGv6eu6ERGv6IZsL7xbgVJ4tNifpnnRabz0uK/oZHb0+zqlIiEw+Ph9CbY/hvDpQR/Vp
61XywgUk0DMf2Ly1egpZ/t+Ib3b0MWry6rNg1eDsqFMW2fkuG/XjdT5T+7MLbk4HyZth/YRCy+Gw
7NuGQ30+EZ3cM7N6sBtYc3h2jzHJQMlthrXk2APG3nqez8kNfykqqh9fE2Tn2RV2cO3qyaDJpdPP
KKO3JPQE32JoZ9XqWRgA6eonZuMkjl8OepVVHh4gwc4e+Blc2fSDGFD6b8U2+DdaIwKvw2hzA3tT
xReNqx8PXfjT131VQx94t/6NrnipqJOch2bW7umwF4tjFxoApxbJd/qTVgxaAXYPymV2MKxrDhbj
lfrDaeeyahiAk5c6mIA1RBCngVgmZp6DqsNpG0Ypq7pW4iMRgf0vRDi/AKzsHo+sycdomVnsLHDQ
xt+7fUnPpi5yd/ZlT1GZO0ZuNMjUhRmf0SQvz97hSa7isJTsgHecv2RS9V2KcNN9n07uQ2dlIb/d
8vLBKI/qfClhQxVYq9R7PHozri9ORBiDEajTrJxM5XXck4Bwl/0/C5dMmXf7YmZgbBQZmJIkQIgA
qA5bLAjj5k6+XHf4qTMhW5Clf+gd5EyqQPYuPamJoRbsEdf3xUMib4d1NdibDk30DhZdvMTyaqrX
5fcLYwmdl2opRGzhEl5QblGXXjFiZKyE6HU6eV/bZIhWH+exOC+RM4deaRA2XjK3JeibX8fFF251
eMhuTYTVOwlouFeXiYhHNAjsJPm5G1gW/0ORil7PQDxUIQkbN6zCZFbZNF3wAuxlrXYJFJVvYCoT
spnTLkBoCVgSz05ljMJgoSYHot1MCwHDn1y4mH3Pj9axyjmzw2prMEwu1TsFHeMYOhusvHpR4zew
7AN+H3xUXbjYzgwYuemaNTu63LP3XOJjS1zqnEeVlMr925c0NVS3Wyyof7wvThaenaRk0ZZ02rqq
PN/VReGLhcVGLGv9MIYhXnMLCM4vM2Nx84S9K12JgmoUwfsLGwadU+kWFz1eLRG+HIHQageY+ScV
x39kGb/CDntbvXSPaR/b4xfR02//QSiR2m1Sb0NaWDxe6etDi/U01Su/pMGI8YxsCRnrcSC+IDwe
IZQNrWxD6WQzBod4edryos5e4RYCRdFVNuu7A7RHkzFRSv0ZmxQ6M4vwnEj7v9MQoq4iSyObpw/d
w566eabnT8AMk2HeEkOhgZpRfPTVXDnN5FsW3n2n/JwrCcU3AZ9og1aQlfrCczWEOiGBqVBc+Y+z
wllygUGuiWDQGLnOWPjlnM02tN5C6A19oH+UIQAEQQzQfqPxZeWNuYsl8ZEvpL+FTUOg/mhP3spH
YSYY5H/mGZEGP+q01zKNlQ09uf0t2Uh+InVxtsP35S0yUxlrPcWz0org6fo3HZVzQdw+sOpu5I1u
0CuF4WK1Xlsi5yl9HtvDkJg8vn2LTZLUGgbSh04/reUCQVEwNXfZjcwNkahG1lhngPVOGvbakH1d
UJmPCeh2wAEa+tNFH19mZrcZuUSHLZ3OxCgfI6y0q/DLH6/h+C3egrIKphcF+Qp/IWllwE6dbjK+
9n7pTskN42iVO394VkpxGSDX2RdCt+BaV5QGr/BOBGzTmKxva3391OImmAZO/iBr5yj5Fxucm7IM
vXqC+QHYlLrLMyGei83UbJH4QYCokOjdGGXpBPyhp14pA0BJatP7b1zUKDKbIFTduiT0+jBrfiwg
KhbtCirvXCjXCtUcShWskZyFRjgaWym9Z9wqX+0SW0beWTJ8N2nd8SN2d05V1a4r/6h6/agk6N79
XyenbXic44jQ5INZhDUeFmkOfpgDAvOTowVpX7e0+dnBz2g108rNXZy9LKmg9gNqoSjPCD6SerWe
4HWTjDOvzrRlpAro52lkiUkOXnxPu/OJoJFajVw714Qr8MHoe9Lmgmz7YvduQBb1XoiYasVIw9Pi
yKysCFI3DPmUmHAb4QTIK3ri5dv5YevdrsbfJ1MAEVzZ/UmMYqTEHNl057YcrogCWGFTX0xb/eyC
1GQQuD6+GLMstFvdA98pQAAnjqPTECXLnRhn6bBgRno+OFTRqV+ih3U466bIqOhe1EAINqDbD5em
noeAeZG4iaDCucJut+5EC1GR5KukNPdD7bQMQFKt6x051EIxL1Vp+Y6FAK9XOPhuzGkinz4+I8xz
yumO6GAg2KUOYYjiTZHP0FTM1vrcVgISAQgagx3DBBls82qppMpoqbU9yxkCwxnIv+n4cCi79mrt
vkT2zccOSPw9boLY0ewcDUHGqJ+o6iNbXuKVXuOvvQ1cDXBOTw8F3YpNROio/YK9dBenqIOQ1xg8
wzXII63/M7eonRXzLudJf1IpFkdWpsPXWc1fE176mWX2MGrgIGICW4FLpWaWsP4iBHjBg+Icna6g
wsq8pe4BLAX+1Z/CSMcMMXIv668chh506pj9togBDiXe4yqYBYH5NsaCXD84KTzLLYRoDzF2oZNv
d6Em20y/d3ApLUJmhViN1lrIBlRyETS/kPVVJ6QAA4wHVNTXL4utZOJOuO+fmS9/9jusAeuabdpj
OkZsl8ZAgqcxp0Gr6uWiBkuxZUCPLlDniV0WiTltovrjcj81dD9HynjSaM7BjhyL46caABe7Y482
spIM5SnN3nHAEc/0WlEUZgnQam4b+iMoR82kDOwovl6XYtA82e0Ve9C+LGSCERMZtTzLAaeyB9ks
OaESBSo+qlWc6jvuUM4mnUkMH/m5Gls0mqDzurVuycFChm4/l4WIpdEa8v8oNLGAKsWDyY8pcogX
aFTEfXoX1EES4aLJoDNyc1FxjbrHfUtaNYCNwlZt7aH0hLEN/GiplKEe4lJh+vj4/LTGB0tOLr8g
EnRS1DYzTAjksJdhuyw0M+VJsl+v8ctyJYWQpIQ8AhXlMtAn/pzNGiKrWlPVC78pd1XgncIT1ngd
bkM/16JCNRhBGVdH9GfhkQ4zsFB+4VVNN94LNdK0Y1vcxZztxcGDsyf8haZ7VO2wrYlJ5zYzUaxN
i3YS+CGmryhuWznl2sOBiYU0TnPyWBhUKSia22rdGSATtQZH4XgqMm97ZAcOJG8B6rQTxNhxhH+D
t9rx7kUVI08I51ebgvK530x8k7F4wpc2sKkf/pqRo7lUDItelO4nMO8fpcmDW50OpY7FFSMvUNiK
673VpKymNjXCJsOheplFcshSl74O7tP0NagQ8fMChWCKAHRG0HascgzttcH8pJ4ceoYqMG0rPQGc
AIrIy8CnoxDpBKF+DIJopa1XJmJ9ZkXTsd3gudmVeGcbCKCSlIqXid7TjbWRmihs66hBlmpDN9P0
LP0oaMJFrsqsfeownA5Tc1jdZQuJGYF08AOg/NCG7X0GJ3rgwj6Wb7MzjXyi+R4PSoKL8KRMoxFi
7YLPcDcbkQ/ybBRbphbvjh5ORNIPkuP+AAXmrfpUaCQh9g/+8guM0cIfpoqlJibr4x6Io9/45dp0
IFlGFuO/BEFJ6GK5gQGIkjhJSGUBk6iOZil5x/Q+BFZXNEt/KtFHWD7lXGfK8uwQFYe7bXMTu2/K
vDqrP7eJpeA57+x/dOZXap1pizX5riaUXpUn6r82CK2PobyJ3A9N3q+it4wy+k9C4kPlqldShLhT
KCOr0e0IGDvhHpUhkk+EQC22rBYr5YRcqtDwhTXG6Hs/sN1ZcfR33k5jRHo8+nz3varR+dEk/oJC
Ocd1EmYFrSnXFhwQEzBjVBvREEB3TxTHMh+VauUu+KXzgTrb1WbPTCoqzTdjyvhaXQEshRXPo5Lx
4o3BwaT1oz4WiGAK7UXjBkllkUWAzZpbxcJ0NRxPwLaSSzQJVvXMatUyiUd5hg/JypalRYparCNI
899mE2oCoTLNeEwRBpkjIAnSejgBXJUrXAAbIjaKXGfppCGH7NGf4L7F9JtiGnc4OJSRkp/66JMp
05F22qX1bgn5KeE3542yi1lKKS9zfs9FSPOmW9VpxVyX0C7uS6ENm/4ZH0A0rWiR5vh92boVapSh
dWbzJl0DPDWHnoHNMzHDOvoe+SeA9H8EAEjKbkFvFRivsRLUh+pd6CF7sbdLRWQJ/aFasvt7k0IK
4z1riGMmLS4bpSQjT8p/zBj4VqZL9lplWG6vdIDGXm14K81GgEBwzpUmZEiXVFVupd6bn5OlgH4d
mAhvDLS0hrQ43NnX5vaH49tN8/3vKu+ynfVbx+c2qV308dfRiuAkJyFQpq+gPBNGsT0/4VhecQR+
QO/4CghONrpCTiI8FLNijCfQ63FAMOZaMxQoYLJFgSh230Y4U2KxmoOiqs09VJp+ZNL31c4baSZ8
OyFJroVhMwjQpBy51Kat+r6r92/S0Qa3hInuuKaVM0AX8oJd0EHB5KVCQT+zXjv1Ta+xrFZ0m/J5
kOTPrS6A0ZmaB1uuA+rAsqeWwxPwC/A8FOF1bLtQD74rmZrnrT0++ZQYwo8KV/LbG2BLj0RT8AZj
lSkf9fAb44tLCUz8VDbwJB7x651/WMsoNEfJF9p+K6mEaxSpvpQ80CjLbwQ9TF5OHVIuLbCmq+HU
xkybtmf09oQ6jgcVbQTRHaHnU+PUwWOXZVKhDtAIUOo7sDvts+a3LjfQuH0mKVDhLejlt6Kue0et
tukmX+ooUQrftOUOr/XoRp7GVPAA0A4GTphyApEJ0UzKdNC3TtL5vJhsMnVbKu0SPSNdPllE0MNT
AtnUeLwbms/Gz5y4bvc7e70PlklOAI5XOSuiByCoVl4Qwvsm1Fo/wanqXdgar8rJVGspQhFUJyU+
CgQot4E9DZMQStF7yy9PHuYCsodTWArDKDapgdOaQX2aow1NBPwJV/OZl6EmO1y/0UjzT+zfaL0Z
vO1G/cJlJ2nSAp5XHE0yYr7h1YDm7+VdaY541NoqraD9F2ENneZ3JluPMsPl/WHqipnqYPhuqpAg
eup6yUOCiIrCl8DI453vRKb88qNBGWDrLSMXDTMMVRrEkaTS0x+gvN9lRo8B//XjitTcouiTiSg4
q+KYtMJ2PXSg0SBVFqX4mLfobZl9So0MkPeHo79EHDaB00Ft0SSs7e7rXP/bak4Yd05757G6REpX
gJb7xszptbf1ZbcCl9A+IqypY1qBTkwYOwkKJwLYIEDee1Ty7KlT3gbqti9Lmg0oXxkD8ytVSM6Z
unVkH1OTOA2LHgBpQk4kkSUtD1bQksOObc+ITuVN101MgZw6V9aeWFjo15Ph+7TEAeMiKXqxz6De
DABYulaP5m3uzPpPEEyT1WYro+uLmUCeYfFFLISGC90pjZytC5JlA/9+V91gZbleuZJu5/nplVjH
CgyR5WMZ6cRqWVznodwzv1DlUPf97faB6AKSKoNZEBiu03IjQ3tWMHQh2OaG0UgXFjId/QrZL1cX
C4vvDVbFwKeNZhI4O8ss9WBCBDpyN9kKLu38bbpqimFJo6CoQYMIhG/AHYbVW2GCbP4dVYJfRVeO
JVCROJ9KwfbcJzA+t+JRNeV1RXFPlXniQKa5eJdXXQzR+sk7qyCF4cNTGGu3qaCkm//e+6q34TZN
AwUB+D8hHtp3Igx/P54PDxx0RTM7GWYRqm/hBL11qn3QncKVnIwAAJldMKsSiOw8sPa5EJLERag9
RNTqHmVqkV9QZxmpAxZG8TYcMNzsSccb3OOfl/GkmAAzVtr7GIij5laB4PiEBNcJRajyPqBoRCbA
CUMpfJJQfOKjeY0bMrVh3XAOG3IVGrVupUhgW81AP/XhJMXo8t221PCefPB9nBn9zfT+cZ6S33XV
COQf23KOc5qtfk/CZto4Yztw4deLv4zPPdkBPkZY8yHhxTZP9pHLIq0IWK+S66LItweQmwxA12sm
eAAQCSjBJ1uJUzA5eWP+K+3UNiQFSoZpY/jXzZpIjphNlKqwFE/x3CgddkTMTt2UJBSD6VOkVKjP
6Fy6ZRKxo1hp9+9ujLaD8UVyCy+YrjSu1hQgiToj3cper7Q6o1d/YqSf0OEloVpz+xK6LD3IgstE
YSmQ+HY6cSf6ysS/CcUqsnpGwCwr3qCBpVEcrTcpaVKq6aK5WZBk82lXTICloFFX7ZiK6ygNlope
mzo4mDXt1ppjywQjVKk9PB7+6ie1R0dYwzFwT2vfdJsJDRqDPaxsyOM/reRS3sIQUMOi+so9fhhC
kR++IUQ+P9E3OvgMMEI5bE1Pnfdg0J6WoJrBgjD3GafosITCJLvzBABYxv2OCVVXLL6/GNvAOqqL
hBwtf0F6MqtEzOIJ3h29lsbAooVLHTWLJ1BdTHWpTWKrwSfqwZ9E3XxKNeeBj1lwzkA4bMC0ogrd
XjkjWtQ6wdTWhgwEf0cIU/lDOnD/ZCcXVU/G8J4CjNuiYaNy3e+qm/4e2J1jJp3jPF56fig34Rde
QftweWn38Yg9NvFnvhsLQNEmInZHcsym/uaMq65NH+Icu1zZEfd2bCHvI9bZO988iPg5L0gaJ4cm
feJtpqiK58oJY34QS1kOHA1339Wp8JGEzBGf+mVj110JKwWZbv/6XxnIwoHTiH0kOqoTb5tw2HJh
7KPOIYunh39E4CzwGioxFoCoKHZfK4vCpxlX4XyrHHvl97vzlS9Wj83lCmp2A53GXFKcTA6IDf4D
PXCQStbuzEqqcP9AH9nbn4wRl/ZtcQJuj68eBLn4jlo/qhLHw7E47vGvJsnARya+ea0IudCBp+XA
aftwathfkIkIN/5IDeUk/KbRrFJ+4b8eOlEnWXP7nS7/I2zI2EbDp3OqM2xdhk33I0fwFAngjTWs
MRdV/cfEfGWvNbKe4OaCxw474UWG3Podw0ePCpBvTYTT7xTx5JxKUlT5yL9NJgXipWb/NdhH3nWh
9ib0vX8Nc3Ca5CDhaLe4tD8CnrgT88SQv5QAvEUk0iWprgIMPvCbsF1uyFw3rgxiw8+jX13wbI/r
j8QKzDJnTzvQEd4VqKK70hnfwSvwXNTP3h17+xEZevrRjBXlpryumoexx70EjMWW8q3w7PbTKpdB
zMEKFJm/DTW29xTOGjBZyX1HmIrJWdBYMH6vPyHnBRLvserIXKkeysaWQfgyZ0pkjOSOefhLoo+Q
XB4hovYFu6S/avs03wV1/bVH8B7OSjbiC5t8TG+ua15vJRD5BL/46bs1yLDiG6Vn21a2V2p8Ff3A
CsdjH7t20ga53efI3SGZF+UFN770zmUmJGVFJstJ8Xa8IC+7v60fhHvjME2bCiddvI8DEJ9tSf4I
6KSvOAmm3pALrHF2I/2KLjm/e8JHGgMB21aF/OFwMWr0W9eMMbgN1M2QvjzOtFk01bp8dzAxqaVE
VQGpDeSrNKaXgBdKRAKo9kBCMKoXiWgfcr6Ts5I85EH9ZjvYA5uXCSnn/3VVfxqkzUH48Tp28PD5
DeQWhHQrU/AgTdd2Poifpr70uFFQGa5FpxpSGH21YrLOirMrwUZTY05DRVKd/RtA2B5g8/1ZCGhg
WcJYXYJ1M4rv1a4IFzcp8dclfgWfjRuU/qHMDMIiSppFXHPT0cMrmANXsE7Ir/0sNxE+GJdf/f32
/s+DtHGMsZ2Fad0pbBf+kwjXPLS1BGLL7zIA36Jt83KVrBHAwJIPlGxWG2PxHYquPgHyb41lVyKD
ZQpNTxqxhgG4vRn+/O6TD06Zd8xOYd4G0SwT8Cc4DNPT8k1jrsBgMzSNHEjXbnkmAYf+YxMc7DMm
Sv1+bk4IIVxzCUBZtmyxzSe9UDvzkjkqhRkErfNLOrwq5TfXSarkL6AuanokU1asOL3XIBtJzO2u
+W742QlN+NamGFET3sfq71eCBAEB+waH81XqDPAXjKuirxd/x/HY8JQ/p/sNraohVqBBSCppfnMF
CehpU2I31cdUgXQmPmdrFLUYHlmfT6t4KdmcN14wfOmw5er2HK7Pl+qnfJpyt/709yUeYHOLYMvS
N/YRTLhamhmqWAmjkjpw8HXYBbKwK9iorKP+NF69oD/oUX7mqz24GspehCiEbftXdRYuCNVKJFeR
KHHKG8L8hYh39lkBO+oNouvSluU2+5nUa6UbdX4l8Oc72Y5Rkqxb4sw/zgCpL62sU4A/eHKfk6TG
pTSkaIjVaPOQr5fL3rwr5gmgUqJSzFxs4H0NNww2qUwRW6i2QLGhdd/sxfBaCwbLHOF0Jx4gzulc
CQde663J45fRq6uxvyBd7Dr07enwlK7S8WFBz97423CeVWBunKLW53VjZn/gra94cIkh96wtwE+H
uRdMUaFR+Watmp2Wfw7K6r1pkp3+E0DnQG1piyw90mFQm6MH+36GaKzMiIIlHkIzpB+RZTjqohVq
XaZSv2NsskWQIVRt69iLZcyY1qKprDcyZSr0GJxxajqDE8fPud5mKOwTCwJ32x9Cwo4iT0KQPA24
HsDO0fHTgdbj6QDJxyigKYITklVWwRLgF6jVClUrBcsyrNtKTNh90MWfvmatTIsFzOV89jGnRAC2
VpXJlaxXqCGWt1eruBGiwOmr+fRzU69f3PUSEEkuupVCQP0YRyUhe5aiE2bePDTYXak64zLqmjWq
RF/fG27dgaNHgb5Z2JQGZ5d++t/hC9MnWqNWmXX/UMOdgzbvLJnClEJXc3jvg/HuztJb0ZUXIZ8z
ILiPxRubwkyV/WzIQGuJgqeSfah7HTifbppbCmTso22HpRfDKwsdnL8+4duTeEJII5dtQ8a1Jgyb
Hqta5GhnQiZ9DGBHDg+B/90zZbpH5+ljtV5GSPwAeKtwYGc07BhBlqjBgW1dH048WRNFJG5Ebm3/
qeDS8DbU3XFL+lkdIZYKZbDBOPJJ1ZZV8XqxWDQtRaU6x+kWYy2zQR3X8uGTIrlHvETsr7MbQiut
4n9xinUrS/mKq0Dj09rLrSqL24G03DygNhUI+XfwNsDUJ1xDMOLH+fC39oygSBmw1T8PRTGickXn
aZ0J80kop51AW5VWtg8cW+kYF1P573R65AaiFF3wqEpLrPWVMeQNCXvvxPzg8airiSooBKvS71Se
JxHwqWsJ1Ip6qwa1b8l+5CyDu2E+0EgmXehgkeLPhejlB12CWNQqdU/9uysaO+BYjb8+cpcxhsZk
XzB2USd6YiRQJpJYPmJr3DvCh9TVPub4pah5Dv6AtBqLxiWTMSLqVanBgMHfBEk3eiZZePkR1WmY
UgJTkWsJ4YOyO07+3AMFzsPIW8WnImLfK3a5VlY86Kq8X5ikd8uS0hNLwOkjocxTd7Qi97C3L0yT
oo5YqwYBNp1avKtGv7kJbglwMHx5VC/yO818flHuWRZZdbQCmeDbQq2Tsy9yRD1YZuvime0OB7Me
6MDCof2iU/XZEIGL8nSiR7behDxj7aUoqhV7Cltl/1n4YiRHIlmPSfOyRth8WFDGDSHOQ+f+9vp0
naKecibnaX6FD0petXI966ezEiyyNre0WDi281pCKWiQcTqyV/M15BaDlo0pmqvGtSAd4ZmcZXjz
9pVhBm6aM0Bu+TyjpipuOmMIWb9kvpbWvHejwT7M64lNmc4R/t3vFaERJzDxFnQinj17SLyJsBPX
pEU3VFKbLWXwTLcRuUin7SoWMDkiY5sCv0Sks5I77lBXIk/ieNd6LmpWEVLi1vgRw+19PnX8ouPv
fgqFfJ7zpjiuIee38MfZPgIRq3VXZbeKhZw/Kqt8PD8P6KKBAn5HcuP9/Ky2U+MWMdgsc6fQcuiF
RiAHfLEPDh12o9p3weqt2GFZ6IPsrts1bOHLvbezKqP0XfewR9LR9gFYShJAt04zZ8C3ZxQ2IPxN
NaRG1uPCn1zQPnYQ9faGe5Zd+VrxuKaX758udij0DN5oq4oo+Uz1OidO6ymg2UFU+6IbNvnUwiBP
aGofbXzfSoqOQdLeIwklD73T9oNXnOiyeKXAv8kyYh+17W+l4SQLbc/2RP9ZLxZ1/pPtMMARMDTx
G/Gp1BEf4WfZcAKM5yrbtHK27+o0QT5DytlpLIVw04yRFrByFLYyq1jTXiBPOaWrjIe/cHrhoUJR
9KJmw6yewQkGM4JAu5ATfcoVcergLl6BXbwhIxM6q35pl2q3pcMxEsO5mpwXUawj+0R72EFtRluY
1ZV5QYuYrCxEdYxGI29Gol0pOMLHhgA+8rFmM7zSKfJHBkB/9QTkHRc3r4X3nMBz+QyUC3zNsnpC
5uPG0OEb702W5iH/8pXXHLlUoydHUfwffNN3i1A2v4wFXWxhvoZrIX2gz9PGTJqcRWgtAOjpAtbF
DwHnJX0v7F2+3HPYV+Z48M5l/Yc/LHsPX/khdEle7yCBgZiDRSW6J+NlinMxmw9VTHPOT0KAsf//
P1jdxWWW5O6JxlDu7UIzvF5XxRjr+DmZWr8KjyIsdgDyuDwKKQwMRgONqnDFhG8xz1L0PMRYiKNV
P+IgNS+8zTWf1kqtlrf8Qt3kC/s93dNZvdH5cLepD7/n384qka387jNevUZ6TdTY2uYetJyw5gnM
wHcDPKuTeHeBr326ArB2ggfV/LPR7fVCaAsF2jX9F6ri4TmYZItV8+EK1KgpL8ZDtCYXO2wbMkik
MJm8Vl+w8n/DmC4IZseSIXM+QLwuIqYp07rp3T+GxWQWgCFs0RhK7+tr1/dILhA1SuLaWWCsHkxD
C3DS0GBtKS7dJz9P73Z/a3AnYlVYXBtdwHqb/RaMs8olb9x3sgXZ9PFC0b/afWuq1aQPe5QwLq3l
RCFb5cOdTIUthIZLWIwzklwHpQoKFkIB+CKRsUz8rDjvMoyHrCuiwRMe7HBfZNomPT7iP7BvzRQ1
HLja3bxuka3OqZk3oWn1DNYl37Fe9mJGJ9T7wXEJR82wHeMJ7MvOZV+ZOYid5oNpgyvtEuvotUE9
MP7B9EnNtr0QOXM5UBCbtz5LahMD7n/WXb+oJPhUcecsqjD2gYZfKGtUfNjiSijUd5dMw8ki4KMR
ozAGeTl5uAdb5KJqOqfBKAMnOSrBBsAROS+G2qGpRPRceWBEguh3/HEqNrIK1Q8SZMabhB38ENmc
lkwAYAS54iBsw8Hsbj6KOKXR3zvyx5y+EGl4rpaQcDKsmXmpVo/jX+dkdbpuvNjIv7poYmoMzrzJ
TH+nxDPsC45Rq80pTsDiHpHCAxy61XlJFWJ47xIvu3cEe0pDSwvxns1IfwT5oynY2tb68riLqiR/
EaJEMdOYdgxB0kGmPx9jgkKA7Vrt3yf4sowsQMKN47LK84mH0DPCKaT6lA/r3e/PhseUFUzz6K0I
1HZHKV1GCji5f/a4AeIBsEjeanQqM0P/ptTSepQTLLHMPbXaJFk5GSbgvk2EUFTkABYSedgT/ema
KteBDaH47Ffdaq0nVZ8ojxRoamhO9AQBdgXEx/Bvit6PaMiV6zjH0qkSPxVT/wO3ieDDapm8bgg6
H7kKf5npueiuCAnh58xOmYfdyf/LbfE3EOhexLM02Ywkq1sSuq/8l09v8ugb4sCiocA1/rzP7vRX
RTY3avC8PIFz0rYTIbq0z3OlyjBM09SmlanZcea+OsHHXnJ4GywMeC+10njJM1jfuroaaPQP1LkF
SEqCRoHFHkznonZlGJUTbiOr7FNBaK2zBY7L017Qh8sWy8nHF31jMyeO83IwzkOKYbY6fdCZThdU
QJ+7u834GCj8Yf6z3qcNZPv3uK6UUCmHRyOCCcVxLyZKn+jL9yjyC1288YjfGu4HwsKjNXX5zrXL
+V0ZAujiInbCWNf+cUbbSKUGu0/IWbtMPFk4Px8WiUj+01PzV6oUW8g8lWKlTfRrosKwAkOz+mcu
NlQ9CRBZGA1QUBDHThqq2yhrMBLTbguDrYEPX0ynA16u9ZEYap/b/pphKgk+03euxPwNQjrQEJMY
wrSR0spxdDdgnxDAxPcEiphfxP5sbP+dAlLQCif6nc0VtbvdWnec1OOTE9cP+V+qkRKqMoyu/AbD
fzSklco1uNTeLBs+9ac+T08cq91+IjK1kzSSAmyrajsRl17wl9P9Q6JXhuzFGxDpLXxcTXU+I9O6
G19yI4FzQQHTykfG8yWBezTpGl6k+bccIW2deo2hSupNCCWen6KYN/RSJNc8AaVTTSTGQ/IVMdDj
SOcmgmbOTjNVVWGQHwbztftZE2JieZThYitOi96clq4ulwaWwZHeU5ZahMOL2XtNBb9MmgTOEaLw
sLYjHqGENS2T0caBZ+w+HjaqBuuXXc9QGu4OmZuW32jkFeAaRE4yc3NBGUZsup0SGEaSjkuoctSh
XYHz/eNLlkpcqytOye8VcxXCRTS9aovvNkK0ppXoY27X5m1TBSPmeaC5lnID/1kiVMnRU6a/90kH
rbp5mmbOnDgvq5GP8CR2DVR+sw1HZbBnEJUHZO2FTjp+6EBN4/M/NFStizebIKdlBSr9di8ZoYc7
Rsm2PsGHQcZhP2bAVT6k8XCEqSCjssEzYaDf3vYURN6KNADl8Sa7TIPZeEWZG+9gI46wknT/PMhF
FN/TwvpsuUIbVda9dI8NHb8Ks4al4UF22RYMpcxSRYY8ovpiXujeCli9TgMiiYZB6TbtwRED4wPi
KAIRoR2v86nYr+kDk1TxmdmTCEQKG4CM55aTqAJKaf/YUm8iTbGLjH/pTTj2RY472ndwCpyWV6bT
97Wl8+ZpaftOxcT8kYuwgbNiVIuwqdBHxW2kBIoc5tlmAwL9sojUQ8aolyK9jJSVMEaPswcm55R7
RqVaSpazR4RMt9iKOYXpL69/WSvaBE9p/5qAj/xgejqSSv3eGZ6rbaaLqLIZLvaBalB8PyoC2irC
sNGAgKZybxgfthh6Et2Aw5HS6qH1FJXrp6L+XTvVjy5KPVQRlikJkSIDWuK0IkhXrjV7iTQVxBxw
Y/oL+6cR0mN/dz8uf5nvIEAaz3LkdS2/1aI0zHAieeD6CSlbOIelbHHz1dYS1KH3IfRF5bTBBfir
hnKBtgsnfUOMPqU/cbOt0X4rEOds8Ma046vda102LGacaWyBu5Fn1ZQHHUgqUrimKOdyi8OQ5ily
ZQBCUvEeDbnfr4oHMD3wPBdUq8zFjFxwLFx5Cii7x7oNyYtqfFUGHFkdRRZpvrDf6M1T+sNFURqK
YbJwBuexUUKkuQ+QbljCVCuaOcQyedHeguzwM8PVDqPcEsLzoCc3f1y3bfFwSmdUJq1vSPgM6q/A
TQv4wYCSOt+FJmvuCIS8/sIGvn7G87qbgkIqFPef+8/FVKixFBY06Y8uK6/AzAWA83gHgKQ5dz7w
aUMOwlq2qx4d3nfIP+tXdHI+skfQXqTmsPsrap2Uka5DzHHjRzhyRTx3nK42zNVrLwdpIAHzQClJ
q3Cprr3u11d3FxC0GSDXoFfQTSMrLjJeOqBeKsXnokuH019ycf0O4W0sSRhwZdgj89GXoo4vFLd7
/2gF4USY0hQYwesL9YzzRJ7VkoAvSqeQoHEZrzpbqXQkMiqKey389yKMPQ18ms0S7VPozMZw0gZl
hDcL9yFkk3VIwcMFxEThBSPMCkt7C3vvrE+SPfHGioV2SkX4UQPk72PScdhzIhZHkcI+D6Mn6/8Z
n3wWlp1WGhaRU7aP5+htOz93cNub87OMvZcCbM/6kFqn0zrku9OAo81eAjE9N0DLFIDcVi5gUqh2
eMyDfb0hCPaUi8RlIvUb4iQe4TWdiLmIX6Z4sAx7vBoTNYAtK7oqmiGClqxxIsXMKoIyetDtcaN6
dixyIwgBYO68bx/UcfW2Q5QtUwFTfewxx89uu/MO2rZfvVcjhPVBNV565b9sx3bvE8rvJIdrIpXp
UFSbZECPRWga616b1ChnCVQ9rabDtFfKkXh+zIX1SjHw7kxsCW3ZJXqa3J5vwU1sJzF53ve1OC7c
/RNuCkRuPl2hpFpoRYhy3aErRl3O3H9c1mdkLdx8Bkjcl9ddSChsiQZ0ZkxHfVxlTsQq3WHya87p
fpi8FqT22KuqIwDNxdIrk8jHdjG09Oo1HM/f6q+B/R/qECu/ByCWMw+MtqOTOJXhtBZbOPTdxttW
WZsOtPVei33Nl5aD3DLRTN4zSL+5sM1pZllNuBId2dMsQqC3Madt+jZmnJNaLQQHkjMa3qEPvZNG
CWNtbNCsF4hz4nAgFZuWKvE67OzUzsZ3yyhC3zczzB/P5YqB0qvmmhAFyz59q+ujVeQGiXqCGmN9
Kzk97A488co2N1a1I65EjjBf4OMJ+ncikWYax2sypPnZd7HBmTu+7J+rVJt2k0HC1lw3cXnw1wdk
BqFUAvdlaWmcXR/Vs1HcCn3DAejeGq/Qie9BtloV+QkzIGTHeAc1UdriGV8WuIu/Qutw4uq9m34q
dtsDQ/iP/Gt2EiD40tHOGlnbPRjor5J5XNpQALyxiNYwCJwPJ758TGxUKAfoO9haY2fYpu7BENyR
CGg+6LtH2v9xmpSD0rQc0EWVJJNnkYZSRzwsBpN83fTaI+8N90+3dehxP1m4JcG3KCnV6T8ab2Dk
8qxJEJ7m4+fz7mLWr61qBGgloc6+pm/B44CMQ6ahHy00tGl8uqtkP6IXBTYH92EKzsYDuX9A31YK
HsqiBieaT2Y+rWJgvhi9U3xMWELTqTOp/3AIZV2tmlzoDwhVF7k6LScvVfVnFWhqTgyOEXfbIFlO
uQQHT8XAj8jM6mDvOUI+XTAZ8JSQT66aXvrQpuScwJixZ9aPSAZUSmmjRqQknarYXomNKC2oqjk5
mJIA/n5bwIZILwG58CaBjoGVRilqJq9t5eGqMSfYGuzf+PKxJeHKO9CZoNm1hOtQJWDl1RqGRcFb
OY2TmWAV/sxKlnXVcDrrEtOSfl3pj5BRvNGjPX3+XHPqDYuHpMOcPsSRE019w+p7+yoyRlodh1bb
pY3kG9LGIeA+RzmrPyxv+1m1L+UrP201osqYjY8tCgTroJ6Z7uRhqPhk6wsdi5Qcluk/RHSLbg0L
1+pb8eA67sDzSVlS8wFZFx1Sxe+l3oqdOgNvX/cq991J+IN4I4DTrqqIwOtt/yFtx4KzTc+uJYxv
haKIg7hJBxUZItqYKXoMl+T51b1CaVNDZ7cbPj1LC337ucO7b7pMyVP6PWYEyx4UW5ef033P7I7Q
707hRMJTp+YAa0cQmvrON+KMsk82kwt7iZDz+V1PEeow4CAgMF9zYHV+F9mrXUW2xMChBL7ECqmO
JpllSClSwkV9tgKipntWXFOW0ehjY6yt1n1mq/qUypYJ8NOK9ly7VxhdgTnBo7AB9OImNwTnGFaw
FLdT/kyNq6kq0zTyq1zGrzkZBuF26OysGxkBZZQilLW72NEUIzcpvvw5ZcC75V80LErImWXfF640
lVRDwGXVM1CHnfa2dC7q0pT/WZxvDzsTgzyJVOnyR8H7U8pekE/+iiVzdbbpKZGhk8NoePiVaZ0g
YuQ7m0utip2HHaazOi37OAgeYLPzPsZ6BFdW15fPzm3cJ6DaBlHxgx4cm5ppkDH7jADjZKRYThP9
E0Kgi4Bhs9HvRCx0FJv/Jn3jtqwAVh4u56lpKrzyORqwbsWZmAHE6JLfm4DNU602hV9ftT/hs12m
wuxsSwl954ItB9L11HfQrDwXHwiNiU9Vdth0keBkEY0iMELxcgToFcYlSVdAU6nTAAN/Bj/wQ3K5
wfc9kZVvnIDxdeuzaJ9DTMzdfThJI455uaOmt0B77t5IDGK4SiHp732wAbWLs/l5jSCgHdNDoX7S
Rs/0nvGAp/16Kj0LYEtvC/QrhPIUU05Jt8ArpWM5QRKxHEaW1sYC8MgVV3YlQvioSEZbXvMkUcvw
pvdYEEvAYwuqT6uV9eNU7lx2LZHyMgjoQji7NLA+xXw4ithv2awLD3QdaNrdamKEGS77KyThUipm
2iQl4yg3Ww7zH0F7/eAso31uW1OO/zzN+av+y3IjTHyclcQpHgg7M0T9JmT0uv6hbvM2MOYyt+Q2
MfF7hfgWUmeO/kvVtqCjK/5YhWVtbK2V2G6L6ReddUM+vkEls79d4IoyFyZlf2zEJyXYrr5xDX5Z
faczI7wQr98kqfveEFHqYSSQo1kU8l3bINWWIgX2BsPnKeAbDxOs10QRFXib1Hoax2CEzVpZp7zk
aQRvFwKWvj8lcNt+tmAvK3YW1AeZnbVeOB8nv6cikTa9aJzGFlY3kk0XQPULwL4JaJ9iYPUtkwdh
E0tUU63v46Cca1CW2dVV1ViYOqePptrwr6KHWRoT1YHFRhdtYn2tDMTsPHKk53tE5UG3kkF0TU/b
Rb6iuYzlJYxf8zLRZVfaTp0Ij1T05G8pRUiU0FUYFZLmVnK/FXM+PbsRRDfmO3E6UfSERbQeWxaD
IU7b1Iphzyxj509Eg3ooqM4+82MhOVKNFvWjNcN24XB4fw6Lbqz8SQTQoGvEOsmjKDAx+AFpUGu9
GZi5n7SWY+MOSmCsRIjcxneOK7lqhZK/sAeGVlkCFMRctOoPBYaXRGXLeyJDwTEHZcPOQoA+OEmQ
jaJeBVQSCWyGUVS9Iai1dMLtXPyfnbOwG7Lmmi3CckOUBZlDI04957eYpYQZ68kiHoE+oGCAJjKD
b9t6LPgeF8gTttnA3Z1eUag60iyVCWia5qA7Ptl+mO04etndwA7MnXEXPQC41AQQQU9lgSr5sHZl
7Y56dXQrDPeUhw5la4ZU+mHBvvAysPKEDmo/fJRkn0VbDVauj4QTlo7IB0wH9WgnCFpY9OJqPXYk
QLd91QWwwiIiKw3jVyaay3S8RCXhNa3ehHIukyh+dOVw/d+H62ab0Nz7JfgxhetaIU0Mqx268LD4
5TNnBEDVDaYn6iHTkqaoFbyESoh+3MzGqF42DzgW0QiCznWl0Nc9MvIPG2roCnFIqvhOWzTHoZ4h
45pG+dewLrOOGa0iTy7U+SqvQFBv63OUivMnafOd90N64G3PelelY2B1WNb0aR11nJMaTHB5YmIi
8LdJmCzxf+0KmjGuD/Cu7QJzjgn9K1iTm8iWWXSIksX8KsLGXoXyS8VefoV2bTauwZOaj88qP88Q
1R8C451zSPDd6wrVzV7wSPV2nzoePmoVQb/t6Sn90UNWIuSX5pB6EQXOf+D2T+PP8TJhdE3ajsPh
YDt0rbFr41hTyGtEmCywYTFfXk3vs7KGWgWPBNRwvc3gWB1LKw05vRv/xGEKtvzhrXidyo/VMIiu
zC3Hqp25W8mLK9wOxm5zI6HiCRqNUgdGj7F/yKzTA8XjRQZWnsDoIqEOP+lJqt1ZKl4HcCukag6p
JessVaHHuR/2AMCUbTMRDvOS/Sow9d/WLvTbWCNL44NAGMEwBUDl066ieOCkFhruhN3RFHS+XEvh
BuAXR24WBL86jqhHT5DuX3UGN9+NvsnvmzM6kG9x/LipF+maKPqKvIoiitrURPXvRQovY5czHZu2
jrQCycy7ZwnGwZUS/7DtYxgir+70SUkN3pjnqWYIYtt8VkZIkYQy1K57KEpsTGKohKwAMRUM39IV
QNUc0bIMTPfVut+ORtUC/7mCmKKLw/Hzj9mlUyh4Hu9tGuPdPLmUXvgzYuKU9Gqrc4kGm5v7NDWb
s88Kc57e/duaO0yimbQtp+EfPaw1xGz0RC4MEQjcQ95RjwuSvQhKJGLISmPM8/dml+PpkmoYkpIC
q7+w9tzSteU9vbU3KVhKI6L7+NsWCwyVChqPyoLpRErGRs6yurT56mzBrhda3jF9wu1MKvVRONpI
LIsZczJ+i3pRza0buudnzNNGxPmYjk6oSgGbY3d6fCKtAVJnaHkBUyY/aNTUZrQpPbtdt4YT04Yl
CZNu2jrm4Wp8/J0j/VdlntgJprBC9RILSKIR21CJTEBQjYLojDVQXKpivaIlzaYkkD25JYHIViiv
sZzOxRjmrV6q4+HkdvAO6iSAO12+Ot1juewko3wmNuOtLOqVaXVtUxmMqdys4L/gHtNx8dz2ubSW
4CNBpmi95iw6vZ2K4499IGrJxXJ7j87YNxRWRAf5msFdBr/IeJtFBCZO/RsRG42WKzMsfFNFoQVd
E3HCsksGZ/bs5qMaJgZJXw7dC4GFkUdSZ3mueMcJnPZ58Ux1MxqjeLDFgUtoctq34gIPMaHbV5V5
Cm7bAPwEKAbLEcTaWeUNE0SiySwBiduiX9iqfTtX3K7xO+hwxt41xS1JJNoUnn6Qwt8JH8asV6LQ
wfr3NaA3BNbetXy6rhpWNMO349rEDBCJP8S/Q7Y0D+DFVsHVEjiBZ8HLWl16K0pQY7+yLfBXpPMs
0lYCZFuDkFdf5SL/ORWlMfndN3teOfnvOsaEF8kb6zM9/9pxqHiUHlUXeXHFvWmR6NEp7pcftRjo
UicuNq3fT0FmyVC4OCGdz9p2nYEjj4LN7utC5W4GapwTQlRX6CBQ/R0DdQk9rB9tRwxmB5Dhycy3
h5HNoOSkIKE6c+uGhP2OeUD+itYxdb21HzFrLsdkUbDlHzHSqrO0ZDikVavEOOHM5J7VqJgxHQ3L
cqx3e6k+ngywe8JOaJkPVfgerm1wBJ2SsG4frQolkCE6qdC0jWOn7lqGnQ5ZiixEfxWtJfsL3Hf8
X4lBClyBcXlycqzF5Q7hUTNqnzz4LawLU7A1q8g0HFkdxwE3ehSQlaBFhycfyQ6diVcz9FqXCfOE
EcfZ2GgMnfz3gvKHES9+0STWWOruPsmWEOkY0Ha8dBaiF0xz2qZwtHRCcqE+RPiSaVyrP1mGAiNp
Dv9W1Tjvo99oVfdEzMzg5UmC0uxSZjRZjIzZoqR5pxVVeXeNMe03G7X3OhZVoans5Svu6V312/7M
EDxl4WXXP93SEMIMS87hE7+n8HC5YmcCiNmxJ/d6JDNHTrpxGhdw5a51NTo2KmizPe2MuZBRondz
KHPpLksmIA8EpZ6dkhot2YcgwSUC1HCtDvXkqFPLmQ/aZ2wb79cohqns5uudvcVVWZp6yrIi8/Xk
7nUYctAhd0zpUe8811vXekUCljJivas2uhW4k0y13LW+4x7M4plXIhmJligED79PqcETZyIpYIbp
M3R9e4sA8MV0ZQNcreoAxcVHtUjnBENbnnldCTMAqVAfTghEcyuLgJ6jiH83K7pB09jsNvbCKIxk
psOQ3PEiKxCOCjbUlsu39+RirfIuBanSnMoEbmmQwYdI4fuC+PzxSEG2WdcnpLAda6Zt76FcqZh/
WN8NnBcMD9UhumLGdB0aX4Cxf0M4xdvhiT3NMTRBNvmhcupZGe6ZCVyZTgRE0/ehY214tiN4va1R
uCF2Pa5vOKHr7WigEZp92FOy7CIKZbe3sjfQPk7OET4cUD2/yCWhyI0a7PwFSIEfS1lJaOZps7c2
bDQ7bXGpAWySAul/pD38/KtRRpfnilJq2Jmm9hx9YXwFKzCij2WgYCT67stku4lbwkWui2FOrBCo
p96OTAd4pi+Ue6cs7u5FdWMdizCF7vQiC+C9ElRYg6bgjAPwzL/JA2/oqSAqEPn8ftL4UOJ2cXDh
6dFZEwdC28ejd4ppYY0Jiopp9Na+4IovOr6TzfBanXW8khD9yB0BIJ64DYJ6gLEbbbzVeu7dPJ5G
D72aCctLRsilp7/KznZf+5GuzsdXEfIUhuUG6u4KEGnVXQzgsD1OC8nfNJliWFpuN5FPmcboreUB
3CGZqUpgD0AjKLqtpSmJuO+T0E0h3sUvmfDuLeUvQfQroiSVVBWqPnRavE39zNA1gwqbDP/KBWqG
oD+V4Vh50NiIte6illVMjLXwglh3URrnrXxMSITVslX3UBrjjiZXk1W9DNFA2m5I4BKXaNLpqUJv
AJ4+Ve3JtTVQvR7sWi6Nkg4KFU/6S9/rfsP4/qDnVpRf4n/ATFd9xfRFHDPsVG8S3iIE5VvU7k3j
WTZH2kCl2+mCQTBRNBC7wlSUUoJZJeSzuXVLOHm+7niwoI/EDm0/Gf9uw0kxOQhdWwjVvrqs/QlW
COl6kk7gpF5ZJu2JfWd5LG/Z2qUPbFVyVb+hJf3vgB/MGfSWVwbMROqFJbkoDVlKtzQlPBu1cUZ1
WUZ6JG1VoDQEKbxKEeWIDW1MfXFSiV/iSq+Cawtsq4Qe6YeL23K9+pXlPozhDV3LAbL0L+aSNIob
CEoJAqWcSewTgjYTNBEfnZ6PssdOL0AhMrPfU46f1btNHwulItnSeaCHlkEKPwRtdf8IJZWchH8F
XN/VxPAyeJ+az9NP3G3+HozgCv2mrqI+vP5T/QrdEYLibR0/JodcaziXk/eNXvdchOXTIsmTP4yw
NKd4EO3L/jZDRwcVjRGH++kLObqquaHObFyDCxCM1N2Wv/GU2ze6ZaRgPsmO3reajvZvdTPpXLnF
/vDDLvtInRp3LUeAvDr1D4sb9rGu9Rl/UONAPlWeIlQ/Hesx0lJPIur6wEGnFREb454Npic8/ndd
RkEQDoTfvKWxjhMtqWqJV2NNRjQQlYC16pfw7iw/pG/Gfl3qKoQraZ6lMCLEF7g2m5dCgJ9CxOLW
43nn7u18EuSmMUwrvfx572Uxgrm0Zrep7Q7mLGhfgGrw3dtnXt1kAHaDaD7g3qK+fI+8KQMc/gsX
JEMgxATtz51aU/vOIEbi0NGJQeF03TWi56ylSebLnjRWz3OP8BUIEDHTYWu24eUbLiVe1RhjBx6N
rJ0nfKmVCe+wXcNljHQGJqsHGFexFBbromPm700q0M5x7W9rJXrhTOUSLssYnd0lzf0x1yVBGCDE
MeO9lN4EHVTwBV+Gxiu/LEV8IMoTHF42Sk7ySQDn+0VqFc7o7ADeq20jx6Amvsu61WG9TMCMMvBd
4LFP7G7HHraR8d3Yx7liB69UHtjSuLkUQBU793Z9GxoCCVToeL8CACu2bQvuiEXnD/g/QpZxK8gd
YCqVkfsRsVJb90M/K521Mkz39ZrYSSXd9dFpjiCC4SX+gkJEtBZdbSSEpMDjl0DO5Xmvtap065J9
IWa/+ti+1Cm7NTuaOCA53cKburdrDx9I5XHaXlwQuqAJcK/yy1hso9TNSP/7HoRbRjuNTlPSQ5oe
4MkmVHkdfDF9Ve/tyb43dTWYwVdMOg3DZ0OMnhhqJOyUJLXqQNxQXRJu9e+KMvIPzQUacLQl8XQ9
PklIl4hlHS1BSN/96fS9rWt1+In3ZBqCTphPR1wpCVCmfUpa5IUOx1mJBfrQFB5vBLlmh/GMSD63
hmpmu4406pOMk9Wed5AMaRfbrW35NrJ1ZiTyNb2FjAqqf+BXYDFKAe2//FHvhvlVNgwm9ku9N50a
/ANr3fvQtxOrMjhT/qP2i1+8BzZ/WnaExIFc0LGww4my60CEwObc7GHt4bjzOdUMiMpXfr5to8Op
3s0YhQmGolJPAAHiu+XKNelDnFIZt6Hy4C18ds9Pf1mgMTg8u6DRv3QuF4gQklmPyMgFLfn8pc15
CtDdXkK0/Lj7cREFGPhQkVSQTr4fdc8xAyjBtLKn/lxcaj0yBBXjbDTWXLeaEdD3YJP74JsutKTO
0koTaBgNydE41nNbdjDguvgbGkXGeZkVELD9RZZyp8Nnq9d9HzoPkzKGO7B3snhyagJ7WDfTmW/4
RqJoAc85TxvGkMUHSV/VosmjdazxdFxgb2GFaS4SqFp6IzaJfD++Rl9dYXbKWRXMWGPtiOBWmdR5
s2LqJErtwEMdVzH7MNxIHCC2FUPan98sQ/l1Z6fE4KM6cK8hUuvAaLUkGippQR/XTBQxXGQ5Mee5
o5Jjuy0uU4F2cRI4I8goZFhu3zg0kB/dG2uCUKWkNQpKZi27uixxjJscV+sPFR7b5C/JXgF8LMY3
q1E1OxQNY29hDwRrZbb+pOJv6Iz1vOdfKwsdLT9RyPEM/QBIUIMzDbmUxzbdytjTlkqOiTq7Iz+s
msapf90rPiJYc5V0u+RUGYhXwdAU2G40PeUUz1WzO3riuK5Lf1jDZV8jJyiaDuAdlzaPRK5bM/zo
TgA8Rcjej4uFdVz9nI1P4ZhUkaLwwGtTg3cVN/fODrpmg65rK++qB4tlJQvY7kq2O5Vwua+jy8tn
OsfoNhsfDwJePixP7/GeUp4sU3MICtWeXyHy/ufgnZA8gS/XQDomK102s0qxcDUxRZO9gDK8S6jv
cjWpHFiSO1HUmukN/R6Zs8GrkNGL8sRfpk0pnBVWLg9RL+P85eOPhgl45k32nnPJBE3n5KCDCEJ7
6rkoLhtTkwv/WwHpN1u85d81Bvy2zGeNbLaLC10zqzwsLGl3DFluGS7LT00ZZpzZDAKZTzYY2Dnj
qlo0beA5YKl4Qpj2+n3roO+1uO7932yTidBtuMJZeSQij0T0ITOoMUtMxmY4l+JhSpjlt7dp+FZg
lJCGkr/jaCX+uxkMyL1ZRRTIflGdkRDnvIdrD6w6ZPn3isMx6k5vxE7BwxAwZDNfQ7XTz2ZRIJda
rEkGvJyLpZQVqERPfKv3UhsQsyhLF519q/GK/8sZJrIMBTjxKhgz2qLCwZDU2ZNtLAnfE/xG2sO3
F9niVLfe+8f7L5irMQUne6DM5bJX8QBoDL04wyz0oF5bhi9i9Ql3+D1S83BcsYlW6B8P+lU3tl3H
HrZQ2ojeJpOGp510kviN4Vjh5jAwAd7whWjsKhuyPL3rKD+w2v6FgWAnQuUgnSE7cvlpoA0qLEnO
dG8JtzFdr4x7vYWK+FYNaMOMxSfAgBfZWpBsBLTNVYYvU0vmOdSDR0g0xfWTUJ0X/u1GMf418hCE
Dab3L4X14YNhFotSSv2xevodwTBaPEzY9L5xn/XSHrOh8iM/WKSGOztUPuRuypXjYa0trU0y1AxJ
IUkQXvnFSGgm49HmB4B3EnjX3/HfMiCwBH3INNUNuWqt6I2K1h9C2XGCvPFeea5Fbv/VSPhHTFQs
P11uNWDJdUnyUkBKL25LyzQ0WfH7O5IzT63wHfjpmt7IC7y88a9fzmZWv4YMKLqkyC9KHv8AJgM6
oA13LSiRMhOL67ElLi19zlxtSM8ghsIjMsnmLGoLUzV6yXHIK9qIo8cZci8VQrlX4wK8bPMbyQRl
jZJfUoO4RS1b+OZyibN9bJ8KT7MSPfSWhLl4FVjyeSxyl617oGBYfj2dwyeha1ATQy1j3xbK+Z2H
88YVWN+AgyQ0GVOzAQkuRKofYPZlLOQtOK3NCOS7zH1O2BOkXiebL2ZD7Jbe9OMvt91rbKBb7aAy
PTO9ZO99ozWpL1tnDUq9+CoIsf0/Nh2cW//6jl35OzR3N5KF9UL8sbnFlST4c02RA3R2Lq8+A5uX
1q8pPiK5PQDO9+ly+D6NLHG5+JSr/vAzwuFVxSEi3+0uFZpKDEPZefObxL8o0BD9s4Mm4O4C5p8M
j9qPtCQRhLsL5Qguf6LVAw9RyCdXs7R+5/n5lyA/PIveJa7+SswryNrpJrjIlGqIy0ax9YMbylAp
t/2sjk46NgwA+/2lQJFjl06tMUtFxXEWGA7LoR3xSnzbXbTFKM3vKt/lm17Fu5wB0iU8rf0rUUnJ
h7DYWetLsxi8EggGdSfjnjb0t00Yc7q19A+7OI+fzcF0iab+VIp8vMzgAkN/HI33YK59fx4sYtD1
X7B03eOitTAvTM8GVd68xrp8oywPLr4QqMqssNqvF+U+h5tOGSZMkRwRMALSchMIQFPS8wlQAYW9
+NvODAjZjnl7hMic2fKn8l1qIin4TMjTImcpZLW2ncPiD7HsDs70Hhkqe0k3ZKrr6+Tzc1RwSn9p
dzeWATgLuGGDXMtoUujLy4/BLe1IClj4mG0A/7/dZifA38taU/FrfZ/RvMlWd9LqWiYvRvP6rYKD
seo6N+EwOQ7+w3A5DpLz6JO1aL40GIijb2ccmZrDrawXTDyaFI81qTAtv3ufMSFFvzJmxP+lD754
fEOo3DjQ6thKbWlbr0LpmCkvFmER/jEDoeOtIxm8SleziYFWEbZmka3yFlyzE3ulVGWpZbIiZV7s
5lwf5QjRQT8VCf2YrtI6l6VRoS8pG5d6JleZw54Ud/oYPzG7AWcti+eUSFZOEEOzeIEpXNDcYQfC
L07+T5Xhas9OvsSHjX9Sxs+Kxqlzsg/pNCn/6UFZY4Y/jSeSyLA1licazmUOm5zBGj5CaUH2HlaF
0C1w1QPEgunHSfqe3Hy+eWpagm16JrcW/jw/HZWMLijLwA1tTrjdyoxdTJG3CeNlilTuXiTnGB2E
73MQzWt4vIT97TPi40r1h8kE7qAF0ocz99o6J5WOD3Qk0BIMK0vsgxZs6qLdCCUiQ2SdjZK1lRjZ
xeHJllSKi6YB07g7oTzfP4YNv+95kCU2uimuKX2yaPOmnQqrh/s5KG2MUEhZLFUhkszGBdmTMXtJ
JXSiIvIZnlJ0GD/R2ndLXsVuFhfKv9rjdeXZCL0G/Tc370z1EUWgDo02+wu3nEeBymgZ39KIoxRy
6WJnxtWqeBGElXLFF2zTh0iKqGkSTT9lQwcaFoPLpz+nF+MY4wqpgwDqoc2VI7gf6yHMLVhnEDxd
bdL94d1SYZiAbLZOTVtxmVvkURB6G2otIvmHPQu3yeTxrICLsg7ifmEkzbvA4/bRtdMWoH1aRYa+
nzU0DkOO1XMhSyPLiwVnpImZRho72iCn4etv8LcKJqeJNthPjWUtVO1gEvXT66DD0hQLZjBtPH9+
6qr0L342znPkJ72ox/K0pR7Ut8xZ0MrynyT6ODW03j7uxm42/UotDEfnG5ZHCWfMljnUrp1r2tKb
ZKhePBcIRJni2B+9P6f7VUgz9Nl3+ZGe78ZRjPrk+GBNNaDX2iysNX4lhCZM74ieQG1C/CivwjPH
bGM9Kj6137/1Va+R3MSzg+fIMHU2DlqOlUHTJv6kCLTCvQ0viXKo8BwRRZmKRfCK/UvAduDAGb4h
Nekb2l2AKsHAzwPwrTfXKPt72pglWxeIj1ezpGMoPplyI5nBpARBuB3CBAZu7WZg2eodkoGiyJNA
bBsB+BxQyumGSSB62YG7SRkW2/sMmJJv/lVhSPFt2rbPYrsY33uy+7dh/v/CrYYsD77fNvHUpgdO
zPUDmSWqtIkiHrhJv6YMcBEDbJvLtOYmvet4WYcv2+GUbxwPk1VNlborlxe5tSGhOBVfK4uAnFCm
TjN94QSNyms68JmgeD/hfPF/Lx3WUeRuZIODaxrCuUWKcHXqr9lRFEjtfRbz/e/BZUgkfY9fbGIO
z81hmiCPZDC6lBK+kmEwS52FGCIS5qCPdOrgs3hbjB1gtfjMD7YzSF6PCyDw+pZB1VWA61VpfI7o
T6JmnYaskRHCylxxMrTESIWZkkJ8v9LlhFr5xvKUS/ir/sIGbeOO2lVzkkQEZJl8ZS+ov7Yo0tz4
TYqV3tkkmWOd6n32DGlsHFU23Vm5kYEbn5lwf5+ApC12bEyQzsRTqvKnT7mKDCkTFI6Noan9sV6u
dmWJReGuRe5xcwxv8PCN2AVKBwLDul/fR2x846nHKt9H+ZlLX2JBo6+onTEzkvtRQT9X3NUWcerY
1KlsigtIEXtVhBhEvALBf0V5/IvOBIuLi6Yjp68qISmk6YNz2hMtxCCTCm+QZnurykBKHfRZ/K9I
xzhdj4co5MiwZZgZ97ZqjgsnjHzQCZJWQhyZrg1Kcn18LmEn98q/r6UuHrcqGudsj7LnwWksm7/p
F+N2qqEkxTLf7KSH1fdjFW71Z5V/PRjOSEIQMmOtMGsE7NiRxvksNe38VdABK5mPjvcQAY+85sPn
h9P0XO46AUsX4bR8Cr+iOJy5DYCdzFUDATFcfD5U7/lgoQiiGkDCbIgERSjVMa7+Hfu7r6X1mymv
PCMMqj+8wMlI8KAlIcFLz9qS2pZR1IXdzZrsqURR7+qFa3sTWEokRteaUfMDFM1NK2i7vhkLne8M
czQJ7mzLOgN/jhw4MHwh4aIT5lpLSLOdQnf3afkyWGj9+ZPS6hK2DFIPLvX3G08oJ/gyq6DEZktG
3K5a+ubRDIda/UkAZPMULYF7R/CX13wqIV5nNDn9UJ1Z/NpQi82e7vDax2+BKhWW+hF7gySsNKLC
fKGjc9DmXqnehs5VgNy4I3EM+kS7LbJLRiPf0W91Pl4FMut5IwXA4jf8OGy9BxYSKtDRxNC7SMTx
nXJyBSLjI3+P+b7d4yqw/436xmd6k9sYIMY2Uciov0R2EuUQmdBUUhyjmw5X+srF0wSMDjwU+cc0
YfADCEFp+uBMAjn397a+GlLF6lk8pakWCHyoGqZZ/JNoccstgRSd/x3XSCVVWfGDeljqiZWo+COS
nv7u+QsF3A1lalpvxVTp5Knr2ghRxg6sx1DHCYKrZFJPnzenQPZItdsKPSTB51A2e38jfc2/3BBv
b/Z8/K3xnEuSrBRZrRv8K3z7TL8GCA6ym5RqVJYDusidjC7JPNBzFC+qPnhWeP5qIMnrnnD3ImHo
k141amEv9UuJF22vVWh/Ng83lZHZFEQJzC1MvG+SGUcg1uri27U1nLsQn5Fs0ZeH5Ux9QirUZBkS
jyTxea+6i8xgvIf09rmeAExDUzKeuRotzBwyXrOqbq8mZNJFNAnPDeuJEHqLko/y4VJlPZGwf+6l
u5eYAC4wdDxGjqo1x+xyzEyK9SaLEqK5MylzaKletcWAYpwu74dnYa+x6+/ax/TqLzmE+y/h1BFu
to48b+mcLx2BbxHq8+2ouUc9fQlGdHXOGN5Es/7W+gAxu3ecwXvVhYbAPBuswICl+UXp259M0z54
WTOjGNToC27t+djWLxKinDWZFIIyj6kXIH8EKohEHzVZJYN2/UYchwuLGUbjt3q8RuDJWlB9hFgb
skXpVINrCYGcFZEwHXjOMDAAamaIqYagq/OvX79a8x6lMlnvRYOIO3SWoEPxQxekOboeyYJgSPsp
iq7YE0tJ2en5EtiMesEH1W4sIW3hqN+NteINTsdFNZ5DaY1K6gNxMicRhJQOS5RnyPA6Yb7dyW+H
qcy+WXzVbm9K+JKE7F8M2q+eIdiNA7bHUidZIR2J/rovSW8vVE0fVg5WaHyi2yPe2IpSH7Xp2HCb
awKeCouyvVLr//QxLNot+vv0noeh+7HcAG14id5zy4hAFQWkfFkL8msN7rb7nv4ipm9r52vVvh22
D2ZtjRkJgl1xu5SO07KtqdyVmGwAbC8Wtp7BPZxbod7Ed8BKIO/CL6J+QZWI6oXxsUL1OOCTDyl9
Hi49DiILQcKMj+PTzp8iBBqoxkCfDyZgXmyL/aD584Q1yG6842JOSceKDIKBpiFdxhBjhqCXiasC
X1dxq+qN67kXPg1QQr+orWCMjHbjJbdRd4pItnChNM0WZrE6y/v9YEwGzW8Bda7JnhbvsO6YlbAk
Cxjjl1I542zart4A5mXo62bqXJpyhZC3oyaGdXp/kLia3M94ivtW9lUV4PRsDz6zejrRiVyO91DU
7ZHIVPpWOHXVrXg79iNrR5l2F0gN+h7RbGvfU1AcwApy26MksZK/qwQLLJqphciUSNrtKieMbhgb
ETpw6DE79OLFQ+IzkYRXn39fgh4OJpG+Ql+jEkpLVTgZIzduXcgZgTLdBbyPy2FJl2zepKPt6T67
0gsDlWav+KH67pNj5oSpmP6TZL8OLQAYxPAaO/yVrAFbAbsXmg4ZEgH1lChviV+ZuAtK26a/KsgW
AEytyq8I+1fdLaQ7nq+OtXTuJzHkY9DQvK7D0l7dcetJp3MOHu8MFhrgRZNT05KMv3nbqtFr+6mE
jnpS9oFsPTTBY3tqT+92hpPaOPCY3uZB1Wv+7s1ItPkPcz5CaeB50XBUy0W0FvzsmSMTrKGVR6/b
UbKBC7RBhgR2jrczgWtt9dI+l3SMXjjIgQ88obE9rylAjMHf162FM21cYAv5KA5yjLHYUqJXyqzb
sqlA2ZRQOpaI02W6rjkqGGESGi4ZRu77AQHqc4GQug40qMbuH4VIuhkfIeY+C7FcK8TwDocniH5p
qMUBoRF8bxaevXnJRJNFYb2BY0+6mgMvizGx160PF1Ze8lnbk2yL8wf2f3hUSNkiunEuM9WBF2wT
J5rOntSbJf6nh0nR8buBvqtYoPSk7D3hYjL6F6/thCNb0nPf5y5FdTxcvxh3gseXSLDRpu5NphaO
Dm+lPuXxDTbStn7ZwcCw/y6tUKCqU1QIVu2UwOYw0J2vnO6KwTUlZ5kxQ7BugaoxX0B/aprX7vDN
FW+k+BJydIJHFBIaO/GSTyZsTwfhNoyWVWhXLwpykr/Z/8dlNe7boGlXkzX0iK2oFX81H8/qno8R
Z/e0Oesf3EYFDjbZP0nmXkG4qsEWEbb2Z6w0HljEMZnehLjh095kZ3d47UaFAEeeOBpLgB3knjhI
G2vtcxXD7+bzM+TugEcKFRyD7ZtwkAHGlToug17z/PzZy5Zg1GYJP392J3Us/CwkFwKsxToA0dh5
07vY/r0lvY9+TmOVCznq22yxz6VkkPL4zZ4dJ/2FEi+STvwQlp+2uQBkDQscf8DkA9yPMqG+e9lr
z2ZMzW30j9J4YJyULMad/yBJPyj1wt2St/CEzAMUFeeXlIOeZt8MPEpW1rPZoXFjC/NG8LQmjo1K
Foyo0+sfU3ZxDYJq3DlldcaUdSTXZ056KtjsuBzGh0tZDNUg8XKH/hxRGhG8Se66WMxG13IxITjp
nSLtLBwGI4fTp7Tn2GOuBvjLvbhoWyoFP0S99qOnpmZ0bnQ5W/LurQvkwn2EZcXBJTWMRvj0WFBT
QxA/tGCPNhrSFNpECRP4hRE0/nQVq59tuqO41kWBxKtEwxhwQasp81GJzkoqsl4MyOLpiEguMiHT
UuRy/WGDxmSCNog7rWg7sqIHuHzp2v7E/ecCMzH14yPHohrbSd614zUtB0P7kMWERorfHjEwKH2l
JbpzvRisgbQDvWrm4p8Yeh4I/DGuCkz3QabjOHIfd9Us4dNghCbsdPu5jG6/j3m/w7uAB5bamCg9
ur96DGq9ydlsBaLm7FiDFbs7IeYgx3qZpVogi3bU6ajnFTN1l1R6riYplawgqewdXhc2XLxSGJWW
u6JmX9XxFunyCh3ZyI9aG67yENfgMG9Lu09zC9jIecBjCq01f3xznp5RDX+oREIeox/vfvkbCwZW
quId+R4PkYZrfp38Z84lS+Z4sm35IQrP8Z+NEMMwXHM3EtAvzcccxxfgbA1F0fSMrzJpgn5/aMJz
7mi6K4SbIr26bN7YbATTD1BSpmbF594zPa68iCzrU8MXVYm+v+4A4jyIFwWr+F05Dmv57Oyh6OUe
nDTzldUTPCXp25j5gBSi227RslKiY5MuJ6vsT2JLlgcf+AaqSZHzCljNFM0Wik8H2PPB+57dAJaj
rSmRtHyQ10qbG/o9dIz4xAmg5wwF756lBFD7kmQmzNBDEfTf4tQAtCzMrUMrGFteX0UlZbvo51cr
u3LHVGnKGMZCBaIZvKo9gGHM+dFuopc897Wze1YIRxPOM6hImco7jUEZm4n5xJkIS1+e+fjmV2LO
usQM14svMGR2YHlqF43Bnc/9SkgnummElR9LdP5ZErOop9VBvNyPKpNNdnUFQqxXgNbbAs4c86Ou
tMMoHoawARHIAKPdPgeMzRlrsbs3b5OAvORsX7ZqcH++tgYEFVmyWUgMERv6GfpOIpqw9am2Vndx
vSXHPThOmPfJoJZVEKWn/ok2KLzGx3hhLx8zMEJ6l+HWEh4zsC0LfOOzA7DmuWiSACUgXti5FPxe
RY3QIOrveLN9LE/rG0aZx0yY+a+K1NSVNzRwTMdY10d/fP40UDxOh0f4D+Ek8wh6ORwTuwyeXgGE
um9wTUa9sBPJxcyA7ME8K+3iCKG4ADeLlfc8YkonKJSJm/Fb7BBnPlIzlcK2ijgMFaXgdoCNUCgU
1SIARzA3dsQpZ6H+ugn8CXqlXxlRKOOgqU0IylLs/5ZcGZFfjh7CN3/D/lJ6oI88i5ZG0E46Se3l
9c9hDtWf+SiwxkxVe4PPW4U/zB4vXCfvKBf1t7RxQY4ewAXVi1O7bwvZ7dlots9YZWw7a0TUHar9
1ZtOiPEe4/WzcC70/iR9I22hVEKPnvCTnysBF6xPGW0fZkwpIhS8xRPs6/1CGZ1/VjWvSe2aHrDW
6Ff2YY7vlVKOfU7bHQAhm+M5UBpHdOeY60bI5R5ozwywtSNxG344HR/+p4syefv8bh4NqMySsnV+
Wjcv3N5D/VL2F3sa+ULXZXEhvrGzitfdSub9sdlrwEVQ6DsII1rk8T0ZSV1h+r3HSnx/ixZk3YTt
J9Xao04b9dGcRyyn2p+JYzzSceVf/hIfE9kDmgsndnluVIVWuilWAEv5dOS9w5pbqn8RPmb4QT/N
uXuf7Fn7O/SZ/8uy1IKhJVq+YW4OxLeVzr+MvsVXEOdZR2l1RcPj1H4V8jG5n5TTQ50cjJYHz4Z5
Ga+TRAbd8Xj2aLAO4Mjit1lp3xph7uZVAA5mDeFyltohI6A6GiJBolKdnS+6+SH56X5OpKJExfon
XmfwWzOgLGX0uBhvbo8tEKqWxXvopZAZc4g4xcK+JDxLy+QoWMCaCdUpAcZ9/eGyfTgUCR5Pp1pC
9wyWuU7mSkSY1YfTNdM7uoeyhXMbKIyAewzUqzIQtHsVOLVgX6FYZk6PIk+kGGdh1H4PxDM/7lCb
+FSs9jppEXEbJgOzw0sH75EC+EvihG0l0aSaKi8F1jO1qZRfc4RpsK7/tWU4RAh1qV11H3RVODZA
t+kzZwakGj/+JCY3ESEuJw6XloY9/MdVZweUXAvV5nY41ejd8pt5vAW2qCOGnC3EPXI+akbPFuCP
6xG4eYXhxCSIRHqgeGHWRFsmmBSHk8SLWSrTzdQyelOYhc3l8xRPCkvC8sDH4UbGtUv3l/7/3YX4
lHr9L/h6TvSnex+lM94v7PJPdp5juxD1XQjYuZJ0zAk2bORnyH3a33vxvMZQILaJGdnHKy1EL4MU
PeIByogSbWfGj5yDd4zhYpO3frG4izJ0YdE8Hh5JTQbuNEmffSgB/jH1OIQ7cgj/N4KLLNdb8svU
SPL2mbgWdVUFXpWFvA8vBcTUYI2Xka5JCz+aP6bwB4upJIw0z87/tdXs/+H+E6BXVKTTyV0FBAxG
g3GuojQsbjQyW/6ZoxI/GpHuaE3qGppn21GK3+N91lSOipCZpwr3CtUDXiwGjlRuCqLV3ZKTsBq1
4skPLf10r5ycWiHNQ5WitZdBYHTeBbIkDcidTCvFYz/zaxR6DMHZxb0+GUBmjdLjoTt53o7IZzQ1
+NeXkqyDLFHZvpI7eTezSxnZOC8wQXmfB+ja8tITb1cgAyqpgd5vPKeLS8R/PRtqo3v619hFUh5r
txHI+XQeRxtbq3AB2VTD2zQ/tM23DF1O79O8vQBHkkJJxDonJDjRp7yRoMonbmLkf9xZIidcCITO
8wN/pWfUohwnnPNFz9bx9QMGXZNV55j3i4wcHSplRBu/PsoLzrQ6Zo/TB0n9+taX7UPfx+m1PsYZ
N3qro8U3giYm7jwl+hREIO5LfS/ZEhbtA1UQ+IawKsGnLTYnEuvzMQVNAFJP+8x2NZ8k62WKkiIG
tUpc7vPZ3r3qqNPMkjz0hqBYD1wzmsVBgIX4P/AOWaa7B6TXMjXHRnjXCOZbyOzh3IOPszB8NZAa
4buUMEIFAMUYot1iy79ywGZbNexp8jLSCwTaguWnwtQPlPMtsM5ohiuWGv1k7wOJNoOXVOjVexyB
x2DeT+DajOgR6gLUeSKG+4b7//uWoORvmvZUaCE6MVYyDcZZecKXRyGRJmIgalIkjMCMOwgMkQbg
NXmVEHmhGC4XJiW5sZWcfWgUyHYbtqv05EZPXloJFMg9Zf8fqf4YxBcw9YQr0aMKdJIcJ/gXS9k9
3eeTf95/gl6A706LlOPm7p8+vucPtEZEY2b6coG8mMK87UcyD7j0q7NcnzUSovfBjoMRuKH9UsML
jnHEBEjKpzR78Gsu3V0/0zrkLFl3/61eV79GGmlFkjCZATKuu+6f5HLmAgnynEv58ZLGrbz135mm
sLYR+/TEKFOF4wH/zEj6U5tYVCiYKoSFBRsNSsqMLjZ3LVuqZh0mFFQph0EO3dBD4+0vAE5vXO/B
LylWgzDOf0OZFIO6BfCmhxuGzvaszqWOr8baqq/Lbz9xXHcg5HRqxwpAj0Bb16jncHYFqJKqgUrm
2MatIQvHVYSUkvTuOCOXv8hLc1XbtPovD5Lxg0aHth4cPqB2CMDm+UZc+yFp5YSnEe8FNgduwjBx
ZtC++3a63Oqa+0p3JvPPTiviSIEpkmdPSi9iIxzQo6F+303f7aHoFFGTL5nwADt8HRl1I6BvAXuq
JvRtrh+H6WOMzZHj7NCSVNFYCDfidw/TmrqdO2+GKX56PN7ZstcqaKu5rDzpKWiND9R1WjVdahRt
60PBLokwH8yJY1XGxbTMSsjSrdum5u04qPdqk643fX+rzGINgZJylU1RQ3nORapUESp/2jkAaaiJ
HIJaqEohL+gbjjUf6ILlKbRoADXLcHom+i4PCFHoG1FOo4pvp0UGl1ecl/S2W7a4WTYbKHBGQwxo
NFztIcp0Kpa0sK3QyBJ80O3K7gtWlZL/nRZKM6VZfVuHoT38EbPXyCd4JvKPkUnpBH0k8Ba2umda
SojRJ13qwoFkjzcMklPToOw7IQH28sNOmNMblQbLd+7qWYIQK0ANlDaYqC/ghbUWB+ZfHamCJ8yT
6SMFGwzkQGMF+aReG9hvoeEx51G2x33XEQDhmy+NwhyfPH4W1IUe7ECMXMYYu6i1+9x4Jpqz1JLr
a5ZMK/bXDjiM20MNe2f9eyqYThRPBsJ0gzuxjoqMCwaz1m/T88JkPeK27IwDrKpWcgvwPUOkogWm
ou8AN9b8wOz1bp3Uo2PpQuibM5sbb1/wCl0vVoEdiFUUxWCOEs/7a/z0Gz/SgGAoQ5BOcYU+g8U8
WavavolyWZaD83TEjGRBwvEDVTuBmHLzrnYFpHxiFpSTmdUUGhxC+VGD5x4umnz+giGuYHTkZAKz
QoKyCe4p69KWcB3wjuBC0yw7dzH4vV7htvC4/1wVxy/GnxGa4ecG2yX93MHx5JDVbLAr13HUHuOq
IeU7n47425NwWT1yq/k+T+2XlMweh+43cUmAprKdLu2fVVFTo7ViylNJB80aQ2y/cDmvmQDJSgiu
cajYtXdkpqcN8shOG8VOKTI8yvq5UKVe7CuNCmaU8WSuFmLd7ZdHe1qPaqyp7YPiClOLfeWz5iEt
nNxV0RH0fBTkf11QOjjyOngx9aCqP9OjMQsJtx3cpKLNJQwgxvEYhGbKqgxpcwrO03XlRYOMcPC+
9kX5s5XxK4++X3PVfjwTiEQbaM2Gp45WLWLIez/cwTDYxwUOonP0uWd2kXUt/B8UjaIOcPFGGcdG
ahOKIQn3YIvGaifjJYvSofpBt+ZoRbu5OCsYfl1jBt8UwN8YPfCqCu46FwgqQ+yWKj+Pkvd/5Tx6
VsOtynwjaa0vzVi3+3ML27axzIQiazb3v7hheQ41aIR5lnyALwghywsxB+zWQdXoJFQaGYQ3U+QQ
Z6AiFkDstCcx2BV5OhU5ARYQdRSWCvxCCeJZwrQ/ex6EEuaF+IQuZs5V44GhI++EdhAXaKZPozcp
esZnR0LkSZp5UMaCRdlbYkDYy7zrwuZqyHiAerDvNUO0ixzljs+GgVnytbQqNbmGLV+RL3jNYpTE
znqn4JU4BOZ5I0S3DpuMLGLcai5Ffvm1HHCEhNA0a2XPtW5ys3Qkhb/JVAdKFRii7blKKQmjQw/T
MAraVmzTv5vCDIqWiyUhDEIu30ppFrJ5mK1K1CszOW1HOZBXfWMq7RbPVxZAgOvhijfh7bWGh4od
GClTqB7DX7NAXlyY1yiEl20Gp/meAjR7NUWpIlRoA7UNNIJA9awGXGt1/uB32CF6YhCXnkSbNov5
b3K5+0bCuKXrt+Vu7Q1lH6Xx3C6Woy2TJRi3taA5ri9fqfQsC7aTgsFBw/lBl9wgOiVVXpjbWskM
6tX77z2slQVEU7mTnLn7HhxK09PdxMYeTy97iJpn5kVx0oqx4XQ/EwlAL8TdGYEMTjuO+l+q31FK
gq6oBvfxRzzqK35fmoQbDkfkDnVW5UA2pzd+fj/TBVhnwAJsNdnUrZbEIPKXqhgLsy8ZGE1fn6sZ
BwZOqfP9zlox0+jVdgMTGKFjLmYqYkiRFcrpmwcnjn62VKXatZIAyhkAVI/7uMx+c/Mzp8mbwdg8
ETZTt7LQOezHlr0ggQFlwfYZRmvRbCZm8RnIzCUmz06r5Onbha/h/ldedrzOW76MlsOqQjtBk7Vd
6HBbZDCrfWXWVmXQJRmpzL7y8Xrki8v8gN85P7s/ZfxXWXDDGhpyUQLEe8QEWj06p1AAyL8IcM3y
x1fWKI86f/lHVX2FMdRMsKuCmFQrGzI11u/MSE9YX6Fildhk9vZQYgIN5kOyT4Kv/brS9njGusZa
i0bXM05llxiLKONxtMPgPLf1dmYr4PSu9odjybaxsqQ9JINOt2z0DDvsFyLkCvu0UYs77RlLPr1E
w/eAdxzM2vMb+zN8AZFfgeH9cGO8SqPScHM95parHQ6z3cLWY5Hc3AXlpuRdDrlU1OXwWs7T5IMa
Hu+Nn5Io+kNejrG9tVedG5/J8ubzs61vDvUEoX7aRoRtpQZW2/VU6dLd/ch7tO1IP7JJy17j/E4N
ZSRjGKVeVcPV4UtlF6Or4+/S7ut8RBy05BmLamq9U1CMxbSavfT3PpDvNKxOS9gAxYgd+L5qWpxO
ay8mXW1JxcjTvyxSWQH1OALa5/fCzOBMtDyhU5iHETuq2e9wCTZ/dqqA3mbGy2H+PradNykOJqAM
QOKtb2Y/2X+HSfKk9fKhYMzSZzxeuM4FQp3GsmetMRBNu38c+0apeF7F/tFHTqE2J8WLn05/biVR
Dl7AMOONFaRbVKHlzCibdPNYpLUvEhOIV1hc8/NWwVAIA+EI5OQTX6HQZkfMy9W0hbp9rutS1jFv
8A+hSj8CfLrI27x0EDGmX525FF1pWcl8HuwGKWab2OprkjxwAa80ir5Cw1MukxeskWu5Ci1j74bY
4X2Q+SPxNLstLnXG4usFQFzkdlExZwSHR/2hw3uL/pMVocBfqwEhVWzfZ0MN8uMbijsi3jeSksEt
Lar7HWVo6ALkGQE1Que36nO4NZR9P9C+IUPN5bope7jc953mv5YYSgh/zgkbzgsMxh+P8jEHWA75
1EqaHrSHgaTHy1Qjdb9yMTf7KX5s8aKAspazEYkI2GLpH8E306OiySd7UpzzZuncyf/gKW7cs+sp
T4ZIDcBA8O2WRQkXJic68Xc0swIbhE+KCxHXxgXEpAwqoppgysM8NMobI0dL3pga/xz5b2IwdMDt
y00hpX0iTsFtEFVLgC2Xj2O1WEdTzh7yJ12FQs645qYXv50/u+6JrsUti4oCB5MF8BfFRR9IvL1h
cSA5klIsChZWxFMxhrsYgd9pMXCQda140MA/C43puTiiF2BlFV9eC/UNqTavaVDp52qZhc1mjXFN
6Ryy3BX1ZvYMPBtss7nh88xFnUH7SA2hQYJ9X7NNcJ9R0LU/CM2kgXquthIsbFn68Kle/5HtE0+C
JcFSd184wYZtWLhLGMI9yehI2KDja25YhAPSoQjN2Pkz++utSgGnvV7rj2fASVdiB6q56DVxDJU2
VwNd5qWszBJmiLP2TfFtd2SKaOKbw3mT6srA7y0hDYld0XdIXyJfhuyO8hAgnKHTTSLpuC9vMFrV
AJv4LLZYPpoABPvqFIr54+LqyeqzGz7Tm5zQ83FLe+5tMuTmFdJ+n1fPmYMXCzGN8Z2uBLshUb4g
ihBiP+67932OvyGBM5saYk14alecJ0ROGQvwvpY2FYEemNPOymjA7dww8vaem3JIr2iaRbYx3yVo
VOglozr/ZITr3uj1uaPOMPbeE9b/4KXRlQRNCNP/XbjLz5g0ohU2oByLphtmik5X5XL65E2uemM8
EBVQcEVsolMUryLq8ams32fvf6irSBEn7nZlyWSHRMFZjFkEDM1a9NdF0Jz54fOv8Apihw0kwktc
XwGyezVNlU3Aw1EVtKpezn/+apxtmXTPnsbNcok7twMWfyw/qxhmTCexPbXI6FJi4sw24PwFAdUK
wkdZJgriHED4OQuY7Grnl+IF0SK1zpw0MbwWIJglmeROxQ1gMcl43tYwFic0469cMGzohlOIZZRz
UT8oGvXGsm35U9uqiD2SKYO4DWfWRMcAXHH+uKHNmpMxKflplYS/G943ZpgUaaaMd1IjlCH3dh85
dCORglUykVzYf3tUwIpenmMME4++Kp6TzmKWd4HNrrBlklSFhcC+VGQw3LiXZ/Xd0+OHza/z/NP3
wZBzilSKHi43gJbW6xYNyW6it9U8jFLnb2o0vNZLep/JT6t+rE7SyTJaMSXgXCyw+d8bEyiOlhWV
PGaORYm0Zu+Zk/cRTcOmPw8Y+ERMJhYGOe+OJpZgT77xnhBQCKvF4qWsN0U6klxbKzwwL20vLbns
eIo7M3+KxiNU1W6I7+Jvq0Qa03wG/IwnsjfRo50QY2dhIOn0MB1V/TdWvbwdQmY+0pARE4+j3K1K
b/ffi2tO5uzMyI/pY8Rsi4c0XJ1iSOyt2Bx382hA2S+C8Ff7hBteTM7TtCmeWeO2rWbfoeD908o6
wR5l9Kzs2g8PbjhN1TcWRfHWzEJ0QAht2Pqai2QcN6Te1wkdq/6vcDfXsPxDz0LWKXg/SicrMKUt
032t8dIRG/3NiF2uvyOBIm3F5DJhx+plEXPZeNZ+e1Yw/wBJXu4uiPUk0gWz7Z6WtNK8yXYaOSwh
oOQ/atDJoK4TS/TlBPbHhjOiKBF7NQ+1eeO1ayi8IgDu/qJNe4XpPR3f7drxGXXxwlthsQCr0f6X
DPycIlD7erdkh4V5znRxIvuK21zVYO57tIrjfFDe57gRUL6SR5++EELJ/SiCskVK4dp9UvmQ88Sl
5JyS0mpHhr+qviBLPoBkxapnCz7coGV80Eoni5YCvuhWrbghxV2P2u8ovlnnfSgMG0FNPodQx4BH
6kJgKrrCSIIPLLu0x+B9GM+Eu918MIZHQIjzyFMqyeSQuGZkktWIhPRg3UK6WekR2yNm8VKuCP/k
7gHKNzoljAM8KrXfQlZIXjsgCesjuUgGdVVBsbaSxKL37bGmjLXfbno6sVAjWi/BCzh12FgKZeSr
+YCcfd7+6Jdq5N1nWdAWU9cYM26fd3rcR6DX0buyXaQHUTLCaSLMAn9sjH/bwRzT8vFZkHbVPQRF
k5hbOG+Pu8QsWUbR5fSvh+1h5EAZIcvMIU6oPWTdSjjNlFGrs3gdC3y6xSw+lhFd7RpH/I8z6n0e
2zbnSePb10RO6ZjVPRqln6XGMIVhfSWtzBGCnnfCp6KfynUJiBqPdYEEs1UiAR7u1A+uTn052sOK
gqnHzh4NpRwEfBYIxo41TUjcVlT9A+cRPK9GQWIOJ1r5dfYFhyhnAG/jCpHnHiWy0IkyicQRl2+R
Th91+RBooHf4NJ2SLnDatjBCkw6xrGhuslWMIOsPZFxJyYQ0iFVXvcD0VreuHtHG9hRz8wzxvF4A
cPeLtL55snX/pFVuLWJmwljJvMc8tLbfy3p/3xXSWdPUwraT0YozgQxdXjuTXBHeAILRAVrNLfux
e9XH3noXYW0ygYEWUemEF0wbHGPMGdUzCGJowAavBB2l5HhM+5vXe/Lf4V01HVH9Ima0gm5V96Gz
YUbVbhp5nI1bXzwZ6grGJ2Xj8WTDe/DRKlye9v4b89ElNxs8OpX/9hzCTVtYDnudftXAt42sTDBm
8NbpT3dEqQXlMUc6Ehkt9fp6cqonEqLbfWanBAb4kctR8GDKrru7GDzJfC+1gn/EcjyTSZ/OhYZI
1JmcZ+7YMrW1dQWluZLEOMdaT6wPu3mqzcy4IaQwOLqt/pWtwYyrqxt6T5xM3HMZYkm8/Xrtibxx
FHCuaK6+0SNM/TYhZyGDNwTMS5vVuF2bxyf15nv460plhRd/PuKF7s0CeV6N1IFvtxTQwsBIfGci
Rb2LE7MZkkt4ooJvJtElajo9mb8S+NQeQZ1Xb14H7vF2Dm5LkOyLNdm6gX83jsU+LPmZFttYRlAo
8/5AetPOl4+A991NbC6CAq/Mu66ZztqYdAQfoWEIlv8ScOKa5zeJF7GqdR4gTheuf3p3phQlpNjJ
dMnb3DCTW8f+1rRKYMrIXqO3e91/fnkn2lroV2NvotqFuUkpn7geUkexEdhML74gNrdiL8/5PsIS
zpZ2hzaSw0xhJJ9W8XRlqOHAuFmIS71bWb7hrd6PycqlqHMpGKeJYXxCvJlU4FVga6RjvRjHCA9n
rMRzL/0X5zDBkl0kCxK8s/4tQ4lCo8EFDRqGJ87Xo0pmUMI7T+yeyb53Wq/86SpxMycN+hhaUPLs
0aUNUSO/aYcrVPGkYOY+QbBFWcUP139OY5JQGBvwMC8ksJYjM3Ku5joDmUqE8FJn5CZzT8fPTbrq
Qhaazg5qv/QeH1j9uIO5+TFVQSSypgcxafa6kGA63Bl+BGbNfc0iFhxphr4VvD1BBqUY/imCYcVk
8bwE2S3ZoD3Qh93k84sasqhFxaXXD8IgZMywMFfy0dpu1nNJQXMaP8FbD2VaCg2Va2LhchAwO2LP
iqtwnF9H4optpWfT3c3eCzMrVPjSk0Rp3cvdg69mlu3IppaQ9h++4OLr4NAe9RbYUr7HD5IatVT9
z1iXsLE8kK+7gCkpcoMK/kET5o6KzQWLEYEWS55FG+Kn3FiNXVH5x3hsLwA47udpPlO2BIaygKMn
lhqjqQvsESQyNbZFNE9dk3bky/EoVecRjoex8rnH52dGYmidTiuLR0kBL1tygFd68e2EtOm62xE5
lFFLcwgZxRmMCxlOa3z0XacPfZMzk4/KrlMXIYvLjqxnXCrSXPBh1AgoRLaAkLx2vo57JHKflrOC
cGjez/SH6UkCmiTNsmvR39I4RbTb9swO3InlIhpsaXPeWkkKpxKgz/lxWR5AeLwyyCETxTbO4rUU
/exTig3YDr0aGr+pdG4DVEZ4yqE3uzesl2I+F32RUyIIGGBgV1gzXmN8NKLpGk1C/zfqF2O+iitz
fZjoFNknHs9a1PuWOp6Bpwoaspo9Xp0IhsOxr4FwHjHAqLI3cwzGBOczYOZnVhzD11B+yWlYglsN
Zh4eJbB2UEs+O/yFrG944clagdhW8Dnkdd1sSWGrSKpsTta1xdG8xpPqF1b0MjVVgq3F8J2jltjC
MVSbDKw+z8U1pwr1ByUZSFskjy3zDvQw8MWVwFDmPPG1Fo1y67HoczdC58dKkCuW6uNiXVesPiTU
iNfwV/VzY9p0Sikds83Mn7h4L4dPaoqLIld/i4g4kMY4muztcQmEp8BY5wUpdQzeT5VTEYSlSTkA
wBC0bPYPkUJxfSP3m6OSiBjfbvB6445pEU72BJk0l87lfQxeQkDwBxp7uMU4va1kOs0/NiSEvlku
sgJeU3fvKHVrqFuqALvseNDTxynC+MIAJcdNBbC/SjUH46pegpPg7bqzVNc+Npn//kcbCR9LsXDj
HgrEdkxNB6xi5sdObc3ff8k/z/nbHU6USmygtjz+g/bXj7hprsMNqMEbY6YCfrCpFWBCl9HxlYJo
5KxMeL9bhCrhhy5+reJ4g7w1WGFa782kDC/VMO0JEed2WpukU5ixnPu6kbK9iflgZKjNgZPxsecf
rv4W+/7Y7Sg9tnDcewRsRszwOyxl5R0c3dASY+SYcc5GlDZZpezPsMd7A0WOQk1R8e0KUQqdxv/U
mSwLsrraSWiNQn37pqjUIg8+iwmh6XHwJWX/h3z/wriKjQUADrG2qEP916GeixwWOJTdf2FI0ckn
CWJgidjMgYcaCVQeW99wxj/+R1oSXCUTGd3zH2FX6AN2n08V0gtol2VH9d9w7XmkDvl0Ezfr87dK
5r8dm3PtN5LE31zNwwCwsqBgmBb/eLrkukjpg8sZ6SZ4bT63BtbNC0BA/hPxUd4l128/hV1QeG5E
qzFhygT0205s9TrektPDcdQOhcOYF9M6T43soCJLdjjZmO2yJq7UZ3tKBwDrI9Qf5S0+b6BT07wY
Kxn6Nlays7jw0hloqcluakwWPw4mKS0CHk3BRd+fEWD/jxrRIELFhrjrebv8/EmRdtH0A1QqZTn9
xL6UWU078CYilbm0MQN5GWDqdZL7Nsm+9ACubamS3rv+4YcBWdj6wT2o3SQzOWjLyiUETp4rb0BY
knBe17ykBQHCd4StG/MhUGF8j5ZmMl8/xom0dbHCV41b4ZHjerifdQ6B5HTqE0Tw9AXbndfp75xz
WMXhQXjYGGw4yGFKsZ75a14Fknkide0k7yKaI487UXIQh9e3hUfnqD9xHaweO291Qe9Luc9L/MGV
zCgY0enY+ZmVcQLl5fBLk4MC+gFBY1yq92Sm1ExEC/eVIWze/T3z/i53Fefx0t9gTzm63X/H7VZm
eQknX9HPNyqsINIoTZCaNHNVF2ZXFH5CLK90ZynhLxTkI1vfpiwFYoQtwXy/5dt6OP80hdaUJgjz
FZS8siuM59IjFlTtzb9QDUg/JxVYpaSEl4qXHwOKSKzwTU4hmWpHLBNi7ax9YCfrBd7Ww4UMFEvY
3zmu3hhqD34FrDSHDjtcvfSi8dTfd82RetY6RUrpu7GLtgb3DvVeTmdRf3impu98WERl1IV6P1UM
EBNBf2WlgIUv9iFXpCyhaX4Z0T9ZTASsuAFFFTU7SZaElOgWdTZmK8eDlkrGqGwBE1xWNNQdbrrl
qYPwW05QbL82NoeECwVZGEbmgGsF2Jx4xWA5UiBq98ABi4PD6g/Z3QfWxbPoJWoT34DDggWBbuZU
U59iIeR/uENSbTidMexzTGwa2oAWv/vhzLur0I0rtF75jwaLdEay24u1mtdOOuF2JpR4PeVpTfSD
HjaujkDNkX91zYb9tXgzzpODtg1vEy5FIckiTs8PK565X4/GbF633a3T0wMBjbCjmD6CkA6EkVCg
qFtF5WeQKm8g+NqI6ddx+zz8IzEHROz7x/DiISxL47XDPDy7l6652b+ZabL46um2daEdVTr9vWkr
k9kV3Wvl3XZFC5lXyeyKmD4PuJZ7BzQ5YzueGO+Cf7rq1COPPQizWtufGBO2KJlzy+vLioCR7b4N
16hZlXbDjD0rQZRaGnzGNeA+IaC89w4JjY9+Bbb/AC8L4d+MEpZhoTgc1Lu7XO+ehlkiRh2pa50n
UUjH7Og8q39XpIyW3KtXahjpSuUXwI20G+OZQb7G9PffkcnodmiOOGuwml27jTLyZqGMYV8XeQtF
sDuskKCs3S9axTUuj/8+YhRJeNILRHxqL2jjgN/L0VhI+o47o493jDQphp+BYuD4ztFS7Cmxj05K
QlBOP2bH7DrANUQouIuSQp34GiCima2ZXon/5G5fy8bL6JZ0rcC4FdbCj8EWEbNXKfM7hq2M/iFD
4YKfc1gVxTQL33L34S7E8BsMbt2ytpuV9hjt5tL/UVQxKtZob708qWka4gpq4MUOBBolPHnKyh1o
qrEfG8bYhyhXIAtGKmemPn/qM2q9U3dAqVkTsZUnpaopFvR+wZUZyeS9D/byCkkADALcdRHjU+Ah
5LxmcCvxWr9URDPwU4q68XZrDdwky0KMUivRKPGqp5hA4pfn9a5PRxfGHQ7rBI6P4qo/lrd0rx41
esiqkBG1fbExUPk9mwpa92Pbi5f0mxvymRupLeMTWJIXK4leA+j9C29mHh1ZCR0WwyfBeBZgykjX
UQAOUU9EhaB3KBgy+hvhBH2jk21M1M+/4VMgi/HB3QC1Pw6lrDtQN1/lp0Usa9I0J29Ax5Nl2voz
v4uZNsBwJrA9ylzCOosVQYTTZJ/PtjYnb9FixJQrirCq/HUqHAG1A9H/8doRYON1vuGNUYHA52pq
38KbSi3wZ5GG6ZAQTp0OQJVacxXNC8USGll6Dstv9YIwOg6IcyranqGmmUiyYRbhNPct+vpux2OV
Dgp+Pndg8j25WPNNyJByrSH35My1cvJLQfEaM0vsOBV5IDV4vBbgRqT7KZd7E8Zpp3O36D9MEfR+
lBm0rmWuoyo10YquheDHAbe3NuFGh9qj2ZhYkEWLu/jmCxzW/arGEEPFa/I1rasPv4BO+/IEnEl4
2tlfD3epiHGuNIHxpXqcIDcVSIaTevEHFlqkTg5fZ4HTgUPjyDEYJfkUwP6eGm/Ip44HEfuvyvWr
SQXcXhJ1qrcsAZpawMxI9MP38qhdCb7K7dnx1v8CZ8NNv47ujkTIEP9NQIp2EJFLookjs+2SWt60
xjjJhCcB1kdjXihKTUAdghJjYP2bVPojlDAQLQMNx2yLaKqzgeP90ilSisW7yCKWiFZwEGrylj9k
RoojbRUbAoTVOZkCFyFRl2TA8OZV+On1z+o9H78KEL8RTnXPICfTFk/5tUrwROCvqSoldo9y7JPJ
+RPguoDVz1WvkdXV04WWZSyZPc4/iucsypTlk3ONaFSBekZRny6jWrZujX1wMQQyglmnXHVNxBE1
9KwFW8UkBsd0UrrpTpfZVpK9nBDMn7GD3onS0LeBqevNvJxMWhWzQBD5P9Zm/aCGZo6K5f9kkGc6
KALXQrWfnRquEsFgltw1bSBP2Xc0d8+3xcR2qQrzIwd1C5g/OH638IoZPkv90fCv6Cd2IgQd8uZm
Wwa3ZsX4CzlqUbHU0899hqnqVkjEuWd3G6SkZJhbLKtpm0hWvTONutzKpOv7diu7wNGDVUWjpyiR
d4W2zDor3JoTLwLTHnCsAbZsACBNUOC+iLlsoxa7lkU1GaUjc7kVjPJN3fDdMDg+cGcDEG5erQzp
rciQkT2WO4t16ZI4ogUjqL9PKsYwI0sPeqg0QWeJ4oBvfbJnsOb3CAhoIE05h8TTiPyZzcdh8Lgs
p2ZTBwI9nd4NrigT2g6cqP33gY3qX91nadozk3e/lm30AepUlth0W5HjRFeV2V1goh6PU99tZK5X
cWrCckC4f46a0vD/Mp/QLrhlif1ei8PXH6vXWi+3YKz4BzGSUW3/XZYok5/sb/HKIfixlyAs9/IL
pesVYp8f6pVh9S0WKTW4m1rYwltx0PiwhCeEqwDlsmLIzEha34y6pVD28I9ZY6AgmvR312eElaGX
KT5p8x8llPKS0cXdHsB5xLsadGyNHLwCBeov+11FVNas2qEipMQd0Nk93TZFzShROMVmEgYKcvsy
aYFO982QVPvFJMfnblXw218C880IdeZl/Nbub66PIqajqF99LT/V6gOMRcV0K49/900ziL/exUJA
R/whEdEQ/Z3KKmrklxku8xzL6SogMowkXutdq+jD94MxINJr/YiErJ8gyoNdXLbIqBjT+9ICr8Gk
nWGgpuZrRX+760ul1lGDzjZtLNw3/qe6xywxf3CA9V/jJLDIji9HEOBdoBBFCOusyRM/GpAeMQO6
AzR4ky5nbxKsa+LSvjqTMZZxRhZJ913aJbV1fvAt1Ly/lc50DceDEE7+8rYoQExzQhKsqm+e+piq
FXLyGdpynK+bfpLcJ1F6J2ioxwT2B+uVYVYGwC3yWpgDnubODWJZCkIQujX1ongiMy0SqIBDz2c7
o3Z+cuIIR1XbgyiDEYUPgYSrMOwO2cLgXSNJHXOCXkUL3n+WzI53hOzqBC7JnahpFZra7XRl9B/H
XuPf5ZDmLnrhwgCz8A1kSt650VoLechj0z3Q3FKCfYvLeI0JjDRUWf5rH3j+gbGokQu4AQ78s1cn
6XuwH2PHO7EbSyFrYljSrp+CmxZDUlfkJZvIgA0zXK92fjut2KA0yAiz/cFC6SMJEaFfWiFayb2D
KEFImxabRzFQ8Gk8nNS1MMGkwSVV41itT/FfsuwynCaq1k1dLw0O64FjQW8wuBJsJAIl65ExRoUN
8VpVGoPvNd12aDOvop50OfUlOUSDq+Vd1nQbpxdjLeSPUALJU1Z7vs+XtKaRpGvS/aBKi/AlFBNP
dt7ZMXhdT1hoO37odb4bj+mXHVwob+m3NeYaOFe8wjhCWgUSi1M8IH28B2D2vPmogQBvat+q0WwB
RxJPyY6NoOw9jOZXesN6lWGK91KulJH5RbGowlaA9XgCJ/E/it2bPrP+wxzHy9Uw993o9fwnaMAx
2v1hsYA0sO5TZDVSV08BoLYwe0OQaSXVkkI1/Myf6c/Cy6L5gKncHCXXaXcl+Cg6hd85UsPCymxB
Bv8/+WqUZnQI0P/YdKC2mTIB4sUYhsrYssNHJtY8YeeQYCjB3BHl1nhuk95PKwJi2onxpJIYWWAC
XXbhWHFNwVfuOetYfLnD1WVXhsWkGk1nnnCGPTUIQMjL+FMM2Q6NcWOKTyXvNZZaZOXK026omwly
YkVx+Y8qMm4vX+WXKdOY743wLCr3kvCPhF9tsGaYdhP4jpXOuuJ3XBVUq4ZwUII+cK0Q3vQVHefI
vQX2vbi9SjSCp+3M7Zrcnvd5j/oDUtnxe9XwKYgZuoHG9JirToccIHRAiqicpgapdImknGf4RkJh
Q5a4qSj45J5z1Fh+ojOAjiJN5bMoM+kUN1mrpfbmEFCRBvKelQjieB2Q7DebYcjgFgTIJfQHMFkJ
OH++GMtkmdGyo01mqDKBeXZjNadwTMnyc3FQFfq5+GLBWugACGE9pGWDdtCAURHesl3Gq5xRjDg9
GFjLuhHyS9Bv9RVmCr7SxMg7C56UVdpDzSaVyK+D9emBBf7sFcQGzWnT2niUdhpF42G6OqO1fPkr
S5kkc6bHIph85j+u9k4p+JRu+C3v9ME1I1kcXGDK8GsB6TUFgk3surhMRecgyBx0CkdJJNHQKMI3
bOfoiRjIBiYE7VzBQl2EglQr9SIFJFGsr9mQGJcOpwXXNZ/bqVu1F6O6Nc8VzgKAB5pvwljtGw07
L/fkmWvB3YYVI3UdXSaFEXukRiCo7EByqdbZIWUJIzmsRv0SHKh9blV1mFOZqjX+j2x603NP7ub4
HDWonSH87Tha9++V2hyIkmWSXhENQ5GedGlL3xgoreuV2rl6vVWgCAVd4J+gR/Cz/Vgtjjca3Rdq
odNcpd2Kqr4CogKv+Vm0RoVnkyyDi1tzAUmlLR0NSOfA5R4kHHilsAxn1Z7xYqmgxylj/TmYEVtk
p91guzojy4svvfbIq/pwTkD1v41LC6DZISFfFebaSeBnJtmsIJKZG5p5TVIhJGzzl6eeLjvecATE
VjhLmwYOtmkeoe8fGfkEbdU91QJMM8IaPtF5jU6gm+VPteXzZ6BBXzOhXZrTwdw52dmX5XuEuhwu
e7CMmyPRgmHIaaILTEEkPf8zGRIEMhiyBm02o5YuM3RGZLupuTPZMLXBcYIkGFxO003A7o1y2FWW
nSmqZ7kSpU0WdVqn11+bQpdn8U8EejrzEsMD0u167jm2o7+Wq8a8NvOtzJUvlXd6ZpHLjooGNWdK
8h0pTDDInyAcifZGvL+BSHJN/cs8UR6i8+nFsJe3y8eKx1zAfkIQCyvuWHDSqw40qF2LdAU66HaU
/4gmrdK+qyygOcOBUnInVUzb9pCkW6Ho3BFKdcqYs9WX5uWHKBLjdckz/ZaMFBu5euwvuMPfXOfv
6Gnu5IQg/wLDBnfxHJD98wock805MkJqcvmBJU885zIRniGlbqmF+r7tesnt98U8M1vhyXenn+P0
kjQBMqDLl7p3OSQmG0/FW+zRCRTNjeSHnzfv4SOszx9k4+yOL3+48QYUcwE+bexgNSzBbylurbIN
H5OKQY1KCLqnIxozxHRiTtHy3ClAelyhqZM22xpJnVGVoWKgx3jA+XjxCIx7y3AIabHlq86HQn5n
5+3xD+/KvnRRpB1NUpR1ZfwVqmROtSXk9IDa6857Zbs0IVBrHZZGzlJFfcsSdkq44GiRbalBo/sY
HXjH9BD6SYG4eO5Ty84KLqFUgiSMhyoaLrPWASib2VM/KPFF+DcMUHCLlxHx3leKfkhr7lthPmKX
r/yEVDIzg9nfWzjzGudig2TFNfGNsn0hqIaUrWKaYpW4EzfHDioXdPhKPXHKwz2+831l5HqcPTM9
OcfAfXXxoz0asmJVMDUk+S0L8nXySVgwaX+jpTkKAhtvYOU+HuzrhpY7SN4SbIloQvPTsQvgiaOk
WMkTKjIGZfL29IaWbxIZUKxJGOQ6WpBF8a55NI2k1/nASVT1C2UvBe0x08uk3/vi4CvOC8f10jVY
8xewtiKxzyfhwo3Na26/b1rSZFQQOIYiV8vWXoROd6L+ODxHUJQeTMJu6A+V10OWgKSn83t8eFw3
qZ5ybeY2A+Mvr1rr59Vc5acpOQDiN9YnhNjNWozfDX6bXl+VNtMScTkPpz2a+hWtZfO9Ev3OJN4B
MXTB7h738C1gzAfWdG62ouaVRVixn9pzRs5aqAgbBgvuOd2Xro0T+ev3VGZwMlVZqpBKu4SEVs9g
pgEPhhxivM7kC2Zo51MzEYBmd4wQmwLQkFhQlEF7GT3beR9E0UsXl1L8sLh4ax6CCwznyVcC/DiT
zuHYdm9g2XXY2+7X1MAAX4r8KDpasCbX9aabj3gpUDFsuQ1pTX305fn1zqrdeWT0dIkr5AsZtFFS
grNS+ZBesTUAbw5uU/mYGgjZb1Neqj5DAtGK9npTyIM/PQg5vkKxzpe+08KI8K7FbBiEM5mXmE3q
ntDDQmY+inE+XUmCLak4zUz3x8NdpFF7EwQpKszjdsyTIp1z03HGKh2KD80UyFgZpDUJPEdSV5ME
LU3VtnXBR42T8uiFO0s/Mbzc81fYnFeuxbebaBn/KSHBT9w5mT/B+AlXeF9jDl1VqOY7UQ5EUdpl
YxBGVWtwCbxpIo0ptd0ow07j5U32oJar5kZ6peGKRS2x82j6Pho+MFSfN1+cDRIdvnGjdgYMl6Zh
DW+4fWKPF6X6LsRSzwNPU5/6QrzmoF1uBjy6xp/kzi7h5h2aEhQpO7GKnaRBZQ1NXK04B2EbUjn4
m0xTeUhQ9rMortGJjm/A+GiEn32Wu5W86/VLZgDmoxiKFPMTdavtG7ZCrOL+6BrP9OmRMGt202Cw
Kp8RxWbu6xwK3pyiZy/+V0Zq98tx2wmr3tqV0NV/Xgl1eAWEbUDULrqS7odnlRoD9tOR8Mop2hB9
Xl1t+p/ygAWKTYOUVDRSdS+L48Dp7OZYJbw64xbR6by3QGVdWVEZsZWKf+w0cfdghWIZvNUT0naM
c9cSN4DCSsyhbLqL8z9z46kpGb7IxwaGq5yVkHb7Xh8jID6JJIxPEObcTcRnUhGUG6QaM2xMlGwk
iQjHtgZRHPcKo4wTW4C810bYKXCJrlIrf49RUWgZf4cv8YHV6fXEcB3g6yitdGKXurBNC3aT2HuR
wUfTA2Id5CGRr9jFFpqbjL/g0Cdf70rWYYVQ0gdsfTax6H5LGjp+/W9cvZ+qDAeVkd3iqObturEV
+3SCdoGNZfQP7+4QOtqegL+BMJYyzQAxabfN1XprPXR+75MSWliQwWhO6s8ygaOgoIacCfgCMe7C
QwNs0svKZN+dM9nlYr3MDFLxkdpiupURa1SdqcT5fZ1G0Ph6abLUfMGyDkIvnimcs3xvMilKlb6J
02YGZThSJcVYd5G9keFD7i/f/EmyHEYQpLRdt3Sb2WsZBobQE3RiuJJ4BCmpON/JyaoeHb6cwWAJ
aGbaLoNUHJ1NQ3U/Nu/6E+UBopDsny6Z07/i6aCFom8je0omWODrd7ZkFz1+w1JyyV5S9ikflbUS
gO3yCML1r8mE6Le5vWduNsgHIwJVaKeycdIwUK9lSa3275Idtqf+kRp3v8VwAO32pG3GmyDFXoPx
Ah6Jt2AyNsvEqJJokcL8+xd7yq789S2D6oVlrFs16gSTQxmtBfTEfQwHvDA9N9OAi2BKtz8MhvU3
aPgJUHqJSxwH3eWxluZ9+1OtM5cTfRBHtOtnkZh2oP1BEmdyMYo0z9hwxcn581str5t7km7/CEXF
e8lJSlGsvfFav05gJLK4DI9ao9tUiOIwxgIRnYxVxV5caLXPBK80pqbxptwyQAacUa9Q0LOnZ1N9
IIEb1dOtU07Qjlyk07JLDyB8nVXJK9sXDXfr+kJ4m+27IYjUoy7FAJvQ5IjopX+ySz1X7jh1GVSR
kX6qlZ38VVByKxn0qw1mQdTRJRgMRM/P5xakmZN/oBDEUBF3nJoYLEB8HNHt3d+f5Pixvn96jNeK
SdodTpew1gneQb1gcCGHLhoG5niDiYSmWp3QIa75jFnOHLKFVDD/A540OcNbf6y0txO/RyVqd/Bd
NtErE/jQ+09WKa3ynNn8M9RvEZvw+1KwSeXpl/2i3Opxcuolm+U8OWy0WL99kyNbO6sUIsBPzN79
rK93Jh9wgYhnTgmXv2hvfh+8vfoGkn+S9L+Mbq/zSxXTUYm1g4PJG/PfN+2m9yRMF54XXf3M8K+i
koNP5C+M9w4UxGKEfKQghlJsc2as9oHv2q2RrmuNij+2KGv04YBhkTpNrXXzzoVHKUCmAGGtHbUG
Ypxe+UfmrZ6rCSInrIEH8A6xtL3fqkN2a4zCRluh7kj1HTpu+UrfxI/81Pwcda0IpQ0njXSySUpK
eA8/DFB2QNzPe0uD4D+glbRV9tcv6eDBwh9Lno/uE6oV9y1KfMYKOFLKwEYYqA45aiqxJxnsLzLm
UXZ2bGvXSff6QoZTphHnYyEZo2BuvOKIaszHXof++5+4D2+KJWqbcqCUgkDdSWWbHZAjX98lNzXy
7lp7P+Zgz+J4glfDxSqWrLFsuuYFKU3kuRKBVbdFhfPbxX+BSZxrAPOMoZGbhizzX8p8bYEvMoAi
wEAqx0he9wWitUjfyOkp9IjSwdPu2sNmZ6cvOVN5Vz42MnpGpGgP9pFnoOowkhvNvXc2sY4JdP0z
rNF1GaaCjp6Hg0DD1xXDJVOp2K1Ds5YpyOIcozl5ozYIWv2ZR7E/AJp2A8p2iVIQxcGf/6dzh1Qn
MkV0IyZepYHX+vZlW6XhSPsC4p78EJQW/dgwlJZJl4X9+hs7RxBsl/MXevZoSPdWcNjgnOcvd1rU
px4HGgSA07FCHWpYpFdQWqwBV2Uc81Oz1UGt6PHBOLLvREf2xzQbLT348s0BuQbSHhzkqWgMDLGe
48sMK7VJoP0a7meMuWvDinwTYwAVttE13XQ1a3RMFaNs58OXU14o3aIuXweNIbilusB6vd6Z8/ue
kBgJunjs9CEBifR3vVHibLNsnIx16jNawnIkI0fpDEWvO6Tc1M8Qjr7aSiO1grmNsMLYXjObF431
5UScvtkHagoFBOiX9Tv2aAmWe+2jFSHQ+vSk+ZKOv7H3DnlnFW1wM8lpAcOyFUkiPU01gGcMEOFq
pn9oEzKax3ziNGMKIYHwzkQjyMuOsVa7TTAMk/ZKgoOb+oV1YLdwTYB8Xr5dqi5Z2Unw67t4nhKz
mYaMVYv36nFVlYK+VOP+q/yMP7mLjMrAun9CuoSQsqzulFTfBLOI78WUAqtwIzNzyel/akzzXQoC
idRZRIyGzQiZQGDRIZvgGzqmuTqfXjCV5zq4Ta801ijgxrtV8CMJFtlyZd77gUj0ilBduhJBSeTp
4CcSGeafjGEfhEkxkcfDwPdgzMNFyhX8n4ES0VCr4QIcmP/aWGgTB3Zz2vNMbqWm62jxIPWkCA58
jGzqcqxUb0X3kABnNnye2uWW+KCWh0Kb39/DoSb8a+PWski4HL6xMVdtD754y57KeLOHU0gjOuE2
EQfsOJ+7yrAN3/AiMzNZfgifqDWQNOsDbOWOTzIPbXzvfjP55qI2nnpE9PxjLP7rOgm8Zu25zIoY
k5FCDWACQv1DStRfn2qs4Ic3yFlIk0/lIx8as28m5cZTdGe9k4kYEzEuEmtiFa2ixIvcVwwvwpUZ
BnkA8kW7gF6bYuXevNFCVb+N4LvUe4VTVsxIw62XJY5WwICi9GFkJe68ujMzZMHtcjhK6iu41OXi
t4mYJsjRs/UK4rSKAVssBtspz1CN+wAei9ia3XzFsaeCX4bLUDWrdRxFTODqMDszmoABTYHVCR0c
+Ju1fzul2e5tKDW308HNXxSQ5j4qF06yk/rWRkH9fkR3DYq4/JKcad/5hIhW31YztPPwBBYvaLzY
rD//01OFKO7qVP4AcXFIaoozp5e9Cw8qRxc6k9iaaaAPKik+r4OlJoUY6Ycn+Gumf2U9U/rq89+r
ywO8mKYPX2np1AXKjEpq9qd6Z+IRFMo/iz0T4e0M0NEzcbp59K3XyhtZWytvQLw2/ZzxDU9Ik1LI
d9E7D1VZREu443iK00PDE80zPiY878snrth0582KN6G9Hwwt6GlCFjKWzmd5a5uKm+QaID+RB2ne
DBaGagVxBEk0xeEIo2kMEToZ2FhEqWyTqUICD0mAM+ALejsJh4/qpeegdQkcdrD/d367GJgS8l70
2aChfTp711HeM9qc53WngBV3RpEPKRNsQ8fWPKtnpqLzImL6X/5ri6Ta8AqOr9K12gbli7gTKv4j
efTvsdN6AX+Xc8Rv+Chf7EVul82SJH1Gbxr19ZUluEtBkSyW48hP7p6XkmxFEFTFOjE185X380Ie
qpzDKMOxNtPi0XAvpcLOyOLB1BdDbdinqoFVmvzPCxrj1sEawv1Z3PAf8zhUJTbYzel5wN2ZhrwR
9WI7enJ827rVaUKvSh+ZzkpT19MeC1lAMgdyXqLXkya/YkmVU/3np4RRjY50PEyKdps1Bw7S7xnA
TossWDMebChzkqryO8h50PMEP9OUDGDhF4racK+Ph98kVb8m3rSWwS2Yh82Xqj4Pi4IeKDW8OFk1
XVAX27Q3WU2W8G9WlJtunwFzLTBfBKBI+neGFbNfyzz24x6z9squuYCn9UaEMyt3wVqGP1HaWJX8
0xu6XmwqHuSXso312eHJ2mwCTWUiACpZnob00GGtwG0PzTbidprqOORCCCSc6mBFzyVqF4oBe2lY
Y7LydXZbEdFtCjWl1nNXZYUupfbxqedEmqVHFbaxNYCReDPurTVGuHxqSEeT0Uh6AwmHKHlz2l94
93so7NZHIRkziDE+lSFWVigyf+NRCMpxWtZU/w/f9lDs+U4czwVAEmSaPXMt+7Oqe8h5tUIIVgA4
9WQ5h2XRbLJu74PAj/Am7DBxNxFaynaeQeK42tFj1wmRwmZNKVG+EeXVmRQCNdFW/K6qJYgQRFQE
g6SVD8nQ8KxNUfyVBHhiExk8kx8uPHoNd+YzxZdThlVmR+E/z+QknOtXJ/JsWT+nCPtmiUN4Mkk6
B0YfbIOSNlXSfj3xLhF480DgfZwbgD+PfogDW1779uJIdc2GfpVhVvdom7sIvsZbXeGPV0xP7x8J
vN5Y3A3S0A06oR1H66b8efktjnpE+luYc77ozHp+zNUVt+3CgELngud0YoL2XQ1Bar9yU5Yr/CIw
KUWYOCaI3nF+h3TOas4GjpvnHdHzdP7RS/AL5K/SYuZiGqNBT2TETSshOiCeIicMyvKrCeeBiqXz
gMysPy/iInpgmOKPemYEqfIWLH/QCD1jKJozOMBlm4l5rLMoMZ3Jo7/r4se5CpPZosYLjT4T8yfK
RX3dmoDjBtIAuqGViPW/+I6L8tKlSJ44Y7wLWpw3N+O/k7sorjn583AEjZjN+uXPlje91WadvOzh
hfwT3JWL1418n8aS4bTF46TknLz7Y8xFyUyTeriT+DnJCf5Q9sNjxDGnL02TwPSUjAMTFMhlPNFh
loJnzyhmCJjHS2HttzhMkJ5f1o2c//ntkv9jgJPMDlw5KczxQ5xW6rSo/Fve4NmGfgt80ow2gTFb
qS3nPm7mGg1k5gJeuK1MKYqzYMLokoyYcZUiTn9pBHFid1R5iK6EIX1JOtbpJOKsd5bWFyw1XXcG
awUgOJSnCxRviRHOjiDmGYF45jWiTX0EccFtBBVFqAv1dkK27NLCxjpzLYla5anTBnR/UR3NIehP
S2dIz74Xkw2Ae/sGG6XCffLjygP3WNrBMJ8AEJIShKJyB+O5Wh3EoVTx8LlXQ9nE0iMJTTwKC8aB
AUXl7YLSeSDzuv/X6wRZoe9MzzwvNFep6Z8JCga41F8ab/W7KuH+23QPxBDideuGI3QV/neqMGW6
zdJlf/J5RLYAiWILjbe0lOS/331H4Ao3jspcIdBc9BHvT8Bdre6u8iTTxsmzMy298ex6AYEqyrk6
N4su0dvXixGaxpJjsaWxlQJcsUuVR9zWeZdTTY2W2ahgDemxGi8LFbgCsomyG9ErXCvcbmwY2b9L
s4yfBNmo2qK18U7HZ41syW7uSdEXz3KCRlMeTJq6Vq1kCiNOssDRiByTaP0BMAD++DDPZ1s2U5QS
vknODJdHuhjatvi+NzHeVfKyVo/qj4pl95/Tgg1GxZqkt4tLuOtWtNm+WVCKoc3+iZp4oOCtUe3X
lPtdK05N2QkhPN0Tq9689kIlX4WKTK6+XARZrQAaiyNVHzp0FMG2XRLH6+psFRDdnmMEppvL5dBp
Kb37jH9T7dCxTjO065HLlImRfm2KZLdhOCsiUSVgmH2Pfbcd9CHE96AufhY7QhYm6iJI4nQhWaAo
UvpQsT5G1HVlyzYacGvt+vSJaT/rU8IJHWBNz7bT4F8P6+vHzm/eHlNtVlKM8wisAYbFI3QI2nqA
V6b5tNa7BQ/4nA7oQbHXQyuO1vz26tOqqKDXOC57wQRijvOi4eT0/tJGxUSCE6XBxU62HThP1RDu
YqrZihT0uUlLOIczkKOSNx1yNAfzGiPI3kHwi36jkDC/hh33ozBrhhHqTIMi5WjlEE8RYI7gmlmK
xu2fwGunS8mpXh6KpqSBGdFYHhHPcjfwWw/JRQ2+fsTVDx8K1fkhU1s26ArbD/SoBsO5NqQ6c6lo
zj7R1ZvAbTSbfZS6dA3CTOg3tifgW2zHeLcj0PKXccLaQnXFgNfF1ZzTWysdBIKVCBPKxCGIGZhR
j4knb531zvCEVmjVvAZ0OJMVMGMnk943EcVjMkHX+/PTgy3WfD7KbKMQ+XkuaHyz3xxRvgOShamE
ShAcdllzvypllpaa7yo/4+mY430zauj0h33FxPXWHm6yy4MbBmN2VTfD5Ox9fsomDZBJVfpSZDIH
tLo0/ev7rcUClMYVkyRqa9y6qAp/nhrcO4YjtyD2+FbdPufs9GPyDWv0TsIMHYdG6tTuAkHq3jcV
eNN2yLSXN0lj3PA9QyBePI2NEwAyYA8v2VIKaiLVml0lu92Es4tVCimM4caD5pjN3rEWZr+mwMF+
EB5PDy/wFp9bHIsAj2ap5S6kvDnbnksFPvbvUBtpu3lpDgSrG/RnnFCE3CckVRZFtYAQWDgR9axw
acranrYZY2XVjT7pNhdhrxydW8yzJy1Q+lIXzufFA8n8w5CwqCUdRr2YW9ViGRhtMRT14BmNOh/k
hM4rNw5sc67uMBOcL4T2djtQ8SpLSNOT0t1DqaCi/xbn1keymzVswctp1MACiNRkobh2+nZDeBAE
UCWietQVvHS29fAbkxXweyAU0OW5oXWknCSZFnZu0BDQQ7DVjrS0Hci/29BbFKEpLiXrzJcl/Xa2
9L4t5UzWOWC2xmiFp80UViELu00+r+HBMNuPoPT4IBuNBhB3DoZ/siE/T5uJCxXIa2YoTz7JCl5C
cp6Yva8m8EZEjM6CckgBmfmjIOI3d6IkO3FYGyu+DKmPrGPQDMpBYiijHowW2Il3lSBNfM6VcumA
cpiCjzl89H0lmA3uEthFt2mrpqiBmg2tP514icaVNnxFInoMcSyIr4A7YjX5VkRIiRG0pxWuRwyb
WletHQPej4knyuiwVgIrYpyd8ggslmRUETD2qGLIR0+zZj1PZyuk2+Gc3sOICFGiHdwJeVz8O0Iz
WVR6qPNMnktlmoCAP9duk55cmX3iO/1Bf6qZxKGI3aeAsCyDr6ypmiZO3Fk9rjYr1xF3fDiBBUy1
H6ZIAfbPvR+9gLnLpsWlSCCCplDlDrZ/xhLNngpGbMEXoxa45RrGlD0MpT0xFE/TT+DD4esNfYwW
Y1mwNj0SY67pbGxkthd3tYfnorC6SV8pVUjUSD1V8sl+ijSlivVxozJL6aDNzqp7i+U4aN9ojNjG
DAwgN1R3xExWoAaV7emPwVuLmn51sDDDybpDQXLg2bKJxkWdfkyjQ4gXNgVEWo70n8Swn1vy5oJ4
ZoFxvOicn0oYTCjoDUwzvHOdK3a9EjDxqnfTy0uvpad1fuXqkUW418+UVtdIttf3/55DcD02ReQ7
FbABhTjI648+BTNWd01H5xqnFg6ZKW5Lpc+wx/caRUku/xGYz/LkpDcL3uiHZWyiFH6NUZZCd3Mu
ApUenTk9lW0EOijubf6xU8zLOLTlPyjXY76IDWuKdht9zFldVlU34ko75bZkFcXgDTLI8vB+pe8b
CifNYEbG8WgBVnw6ROghlKDAZEcF/k1112HTYHXGmlSe/Zz/0r3kqLwN9SS7foObhJy+ckpowjVB
idrqnwuZ2J9HAg1X/6Gm9srRExaQsnKmcMgKLRErtIV9srXVrGGcD54Y0pItQT6K6H210yO9pEhY
Kw3a/P/AS06auv/lbb4Zc5skj1fXrEnMHmP3LOk/utv249qU/+z5uGnLLWvNTCdfc9lUB6slMG8G
H4nziy+G/GGNxGUYdGKGslneC9wZWrAVfiWsBWt+xCxifKdgS9scuOHfvF3y3Vb/SRB7MX0FtU8C
oVAt5mVBclhxxZjuNiPYjTZYHAPXZMaTWsd9z1wEDL/p5qLuX3qsT8m/7VIypYtGbubgpCOcpcQi
tsk3u7lLUSl172BZHrd+Qi3Fet31xNCsYqQAbo8Kg6sIrS+rmlRr49qov6oJwHiOF8lTRZbAHLsP
5DLW97J50FtPvQYahnWxdZ1XkYG3k9uutP3Vj11rMo2NjEy+yatJE0PLNyDi0N1RAK4UGXBjMlj4
JIIIGBssHkddtQaY+u+b/Cd123rwtufuEVoNg2u3V83Tge39kSyCKbApqrfCfgBNPRYubHMbjuzF
eLiOWaDq0tI0lRXS6lVwPenQDmQavCPW3Z8fuCAoz4Fg6ssYNwKE1My9GOE2Q3SHjT99hzyCmMkw
Ntmp0JG3tz0kX/n/2Qxvi1x8RXSeUIDWm1bYXw9f508I+FSM9JeBcMGLBelHrU/bVoZCzNi6bULd
0j+nFpXwSgznF0mFIDCK8ZMu2AEkQE8+/bxIxqcYvB7yqPIZmEEKoLKzIOM4QxIX+tPVjMV1BFmN
Nz5J8A/W7envuuH1H5/8vS5VWAOzQulA45sIFqva5ZEgYMcAFeaU8trwHhaiyOWIs4mJdinCvk1C
4pHjf8sXOMryGqeGhggJMimXKtl37ZyMBwZmMyZ8gxqkCnyr8B2L/9wsBM5G2UBnOe+X+lVJO7Ry
3QoNuOb5i7hqbtU3H3BaPVmItkW5hdRJLFaNWkkm/h5EHQSHEiL09ZskNFBBfjF/3sMEapOd0LHZ
kvv7D+Qvk6QzqUv3AySYPHmrsiGPlwus3CDWnzrFiqedqoBZDQZM2/oo68PSjOiPTyP/JTXcEk44
sSH/Wu6n6+njEwmV3DVyqtvRtA8f902eGBaU9y86KbcuGTU/XvdcoWkmF+GJsvEY8KJ5ZTmfMmNd
OHwB6LQhzGRvJIYjOkbEnc6JbgkKgTsz0awytoSzI5BQCn31jC4xgCjHEzjquZhOfVvbJf0UHEdh
6up9vcWmjn5whpJsW0qUgpAMEm1OjoLMGOXt9OU6nMTZZnTBFS4N4ImRpC5mCpPZ6Szt8UA3WuKg
wMI6ltJ6wA1Q5aQBxoPxneBUCBAfnSaiKFCmfrKrl8qaqfWCfrFOwMKHf0dCXZx6kPXkHLkWZn6g
foFe9Zlrunf+TOTUpdDWSL8xLMx0pC3u2/ddCH8mdZs8eJnEUPZlFAZ7Q/oU+dow4ffU1lKk/dbP
nyso85m4kDmtdxpo4a0PV4tspr0js/aA21BT/ff/UMkmEVnY3CxRVEE0XOU6bO+TWmuD5CK6ySdW
pdcjBY8G8CVALN/MnnOfg/xZx+X7N919JNpWAW/sP1sFCJFNulcrpgfeIR95P9SLFpPFBmUmPVqd
A2b/1FEHvu0rxAITCD6R4Iu/BnKnc/trnEmHrdDfVsp0Je7mgavngCfMZrnlh2gtCyY6rmh7Tt2k
GjYs8es57U/dxSTAWKfjRel9AqRywK9YjCif53YnLalbgGkiBVKvBEaQxmEKxtw1z/Vqmq5aCyQz
AQvB6Ttay62yfhacb6y3eJqQJybrOyjnbVT3qSWv3KOLxmlZqMs/XZ1mpd9CoYf8grEfQULcuc+O
f7whd2nkUgGd2sS+kuz0OWsO6rPE2VR4H6rrErHmdcztSKZNNckIR49yZd2AtP6ZK57HLr+xKF7X
0GT/jy2q2wyc+XT+Ahey/ioPg2zFOqlS16ZOcETnctIUKIAJbCm2WkznLHW7TxpReTah/CFaSbmg
yDK3pJpF6H3pfTiFeKwhDCzPOq0LmOUsBLqjmKbqlPQjANw/eJOE2X22bsG9WereI2L/A0POnx/K
8O/ra59h6fhGdVCpfS2E1m3FAr/lIRD47wtzNAILOlk2rRrnxg5oGDI4QcPbMGqN51s/g0y1ozoz
oUk1ztNszdvJIgWYLggIBFqtAWHMuRoHM9+mbQVdYICpO9s/RhDnhQNQ+V7/JAFI4Gt94OcQVbdi
yWuitaN/x5tkX5uTQBReRhgQBBHCDRmF6AvCjn5NnS93PtoP4TsZ2AtfpvwZne56KJBGKPyDYb9k
KuwKkTNALG4VYvyyTjoQT11cIkMLLCwI+HQrlUhkUrb4NNgMtr/GwK88aP67Yj69elE5JmBKSTu9
o1lKoSnWL8F1hxTy/8BbzohUPGGjZGF38JBKAvRy+AkjQEMxCfeSflQGeeGvwdNiUUGpdoz40X/F
lJvfXPqqwbgDKRSqLwVz0RZchlyQaBDmpBg+D48w/HeVsJkOBPxUom0PzWOVMawhibr2tstinDU7
4eiLai+MTHmIWrl5fyeTq3AYD5IDSubLStXLwIw7qV2M8EIsr1Jg7JWP+rEMQkXzouR9jNTtOXWs
Wfsszx7/zCYqCmvZ3AmM3fFMNuJxM0ROQ2PD8HloAWUJVHaFhO1QdCUNF5vDt5qqy/BwsOd0ft9P
ykbwEasVPLdqh4U9/oKqmk+nHSTcvOiZB2V4p8ZuH4SRexgH/zeIztSoGK3VIESQjRZ2Ow4i2eU9
NPeFpixaoSOr2yQ+BNiuQayN4hdi0O7PwRno+ZXaV+vEtBbc6LDyNV91iRBIv2nxV3gt05ts2AdA
lATQad8Dkuo1no1NBENnmQyXCPUSQmA0PTBWVMS72toh+dZJl5l0c4I3JUDoC6rIV40GYPSZef12
7smWjEnLLQiwHWYHhenUJujUMs5Wjf2nAvdERJ/4QyisdDgJeDtZeTGbccm9d9I5Mod4gAeIahTj
ZkqT4YKy+sO1MGIfvt0FQn1Gkx7a8O8TpGjH//FRaKIOHoXMrMpRe4VB3/pwavS0MPXru22TLa23
aN9o6BcvAmuchmuqN4HhJ7DhPhS93FUS8S6jlt2/+CJG5o/fPDmzvNQzoTVmIlJ3Xahk/pnJsaRn
/Z8ygI+s8TjNQqQuYjcmmGLIDmdFVXRzwu9/TOEyr8IaSABXnCJ2gnTmFHiMRd6W+iqsqnggg0op
SLtiSQrtXRpSP5gXTGryXyIMuX6/tkSfCJ6OOlXaZ1z4vGAEpXU3MDh/WheuMfOVA3P+GDsiGBxN
cFJ1LpVig3qHSlpSXPcbT2TNEHmMpi5tbNL4APwYuc+niw3ySeWlv2linEJ6844jIC3wKgMGO/g/
9dw1jlSosyWTNNcyq4tcJ3GDNBFO9OxDdmtgsuQbjQ3aHHDMHtkaulhMW9dAmz3voGO5iXIdUUAJ
w7dnQ7SBFo15F8OSMSk1Sa5pSvNUlj9+HHDj9TYA2P6gPC3twpmxnBBmUavms2IISzGRVtRjteb7
BMvav18RN4TeF7rrergWw6BbyI2P4M5OS+b0ylniPgF8KgMKhUf4hh0GMGjoLaLI72PF6bj+t0ic
W0rzNRg2IGgokeyDsGcokfQUxbuRjuuBAGqr8/QoRoIDMaURJ81PksZHzv8W+Thf6B8u+r9axuXE
qiy/kAMil1ZabP5mMdOjLTdSrZQ2Z5Cy37Ps+5Xwwach6GcrhXHVHj1KbZzpi/6c61JKEjNbj2Rj
PBK7Pu6KKCQm3BoEv8DpHe6W0WGTjxOXJVYhHGFqvoM0eASmnNnE0lgQp3g5RJ2TfcpXfkZcZn/J
vuEIDS1xkBuo+n5FiYUFvLFXtDQsHz2yw5UvixMVpG6MTE39tVE5O5KhKVIHT7RUD4dh7xYeGNuU
fYgdSJvZEq7MZrwTdl6cH75sMjW6AfpMUb3GFiV/wdxEvVlUm7QQGGSV38f/2BI/rUogUoaKDoTm
/MXbNHpaQeNWA/MuWYu3J7S+1NNF8leQ0E8V+8KJBnXNB/Rm26d/khyEs/ohSVPs4uSYtdVxg+nu
e/Ez1FoXGu2GzGXYy+uTbwQI/RL9Pzz9zXgNAyF9KprZJ7ZxxuwKho9I9yDPRopmk5JcAhkhSCHJ
Ep5hEEhq3uCnoTda2ZDMYDV8To61aPu16k39cNhk19mDAAO9sF865ONSF5aldGFM9HfyQj7PHwil
gjjQOwXalSMk4rc3rSIzeDYi0kpTi2CP1KEay4GumIdjK8+Ewc9M/UQjnBei5Znd9ICZYShAkivh
Qjqxe8rGCDOrYBePTJZe1gYlsHuRd97Outq0+SQQ0tVqmD8mdiiJYxgTDJsfauJNN51Lw3hmPiZl
7vyS7zr3w2FzaSzrDTtydy0sBB+YK9VbcahQrHbqRVbSA6zf1kit4Id91mPsdh6lyBjtICEugziF
HWe+mb6OWH/elQcZWvl8Ip0oJYNY6pkzN6M6gVqtR+XIg10pFGIr9bOFViU1Xgh3WdtPZ0//plTJ
Q4/aIMbaCjoELua1h+DihNH21E0mVXkbAulCQzU2eANkwhRz3qjshiAk+frTaHvn1JNJRDUoyhJ2
za7Gf3tiWnSL/o9GuK9xdQ4TehqHKawzTBWh5iLF5snVAjeHkXyfZKKF8eqcxIFXqIY+yKbHz86o
I/K2zcS2nzFdcLJBou+0MP1kBHS6y/YWJ2pBjryx41biXl6xKGMUCIaMb/e3987SNJ1Zgam4dCLb
cE5ixZjzOCWexBr7551L7iHo9WNw++SreeLYQvPAgJqpiE1rVd9I2Zi1vg5BHEq82D0XMfe3lPcp
V30faGp9P6LHh2C4ay4qVcV1Ix3+LM5jLz6Yu/wJ62wYQqxNGxgAU0y1p8Na2aCB9pT+rgMK0rYV
9vlpNg0KzplJ54vN0gKvfES39VPfp/SS+RteQ46VMgFXZJmx8ncaiNBJBkdp5agLMSHN64BhuU2b
tNp9LBr+TAhVAQsFpwfvlN23WN6lBZdUqQGszjcFNY4YjIMFMM58XaS/sbuFpesXrTgqhXl3Ruom
11IqMezHPngHzb/blioNt+Wr8dhBx/XLPulK5LzRM5RWy9DnOx1dAu1mMGCnh3T/35jVcaEVRyPF
VI6677fmb59+MQ+ch/ibU87YtIf08IVKGYqbuQC3tVFBBXw8gHCUxjh41HTiioJD3HJDVyc1/Xse
JlUC3hUYPoLx7ILRjHdOxI1m9wiS8rl9UkUhOQouP9ZyEMHpu4Ndu6Kz0wxWAbfLclYPhHKdOXoX
sLUym5g9fJsoYiGPM2Bamy3ILh8uP4+HqRlVJwA2wX7d5tmXWPdYieCgQ6IHwedl0rpTsz9oRsKE
LIn1iCDHoLmEWq/UXyTGC5he84sIeQu/a5lWtImtBK8tOdWRivbUm42ewpQXmYFLsyKY5vMKmtDP
DsZI6+vsBIxIxaUjCiiV4rWA8OHRAcNQilUbugo2N/+2mXRWXbun3gETgv5tPJIWZgiHkFkGaHLC
X5+89hnH5hTgUEj0ERKAL4Bdp693U9FpZ3hqkMpihPzM9JjsVGaNOsiRjYmczYyDNbOvWUAVKsj/
u2fRo8zFahj1wVl1PMfhz0My8h5gKRvD8YjfU6/ofJMagpftUqSspyCeSjqvWD8jaXPqqeBAhkOx
/D3zMGtysWoAHOB0nHcML/U8xpJwLcRIqGYQFT9tp6BDf76DjFnCu54vFMceBY40AJWsPrgFCmPl
fcDQjsWiMLMfc83l+w20GAPtRmt/kj039W8i/IKxjLGY2uhQ4Vo6wHIOn2hIw2Nuj1cjfVHamX6q
t0PD83NIPdSs5955kk9MA2FTJDyMn24jhjg8oU+OQ/VcbVPQlAVP0b53cE5J87knE1R5n+MNielu
xloQFE2BEJZ2mC5aBmnO1SlSOz8Sq5CD3yq1+5U1LmGOw+I+yCmpxPXtxDm2MlCL2FYRSrx+GhsC
M7LUNS26nRhJJMxMwitOuuZM25pjbPE5YU8Lx6qw+zCRMtBv9ks+++HZJwWRJ8zbmLTIL/Bim+8W
mg3ucEZr2UHeD3yUuWyFUUUju33Aq3fD/cCO0CZVs4tGWo0YIHdElNbp8Ve4azA4MBTizmT7loQ6
IyRpahykpIxrJJxXE15A/YmNfo6LPKQVMpqzoX881pXguI8r46qHRSbA/Jm8G8SIa/1ccFkrlJRa
pEpEnqXFlv2F+aXeJnPxVkz4Dh//h40H9Ohb36U91cfxOKUsi/vLwvXVDarGazHuEugOGa0n+qFV
voPMGDLo32KxHmYUn4Ov/95udVc88bgqBAuUgF+uuxGuYpxZl/kNu/rAF29wRXuLGiz5+Qd5GL3+
u8f2RG9I8t1Lsi+wbNU1KWGoOwY4JH08gmsFB0kUu2U6QZSy0fTqcfZEv5v6boXyY5B84+Dbx8QY
/7LirvjKe5IQqAjH/2+IbugR06Y0b00atGMZAJNaKnotQmesdRo/mrb74m6jh2k3TnQ20s/BqcIN
NQglc2NXB5DOcrCrCBux2EWUZGWBwVUznFU6/ZKr5CSZjzkTdxe/+heptB3YHMkWZ89J7hMIcCsn
NsXxE9fF5tanCey7HpZUyqYvm4n4Hpjw8tuVxHh8IApxU9otPbsM3vinnk/dOUbuP1DoFTXeqp9X
hUHMDVmkb/pDNUYc1hUHKE1fVGzMSSxzNk7q92svlR5PW2nGU1k9Ynn6Yd+O9AOVk7wlWKwqTv96
Xa/ArxtgeCsFIbmaeaTvJBJMcbN9p5wJqz/Wb+nuuzGyPl3DnuBBl820BKfa1E9jASU9G8739Eq1
LRPIXOLg/qeV+wbn8JPBzye4grBpfP9G/YAi7ahgQQZX1d4wBbIpX8tMRC6jXwKohzj3ccTPb9sU
Y+JLMxG8Q4oTfOvoxFSNw43C3Rn5Kys6Gi7sZIuBY0I+9DntqFILEa37sSQYvK+SiU9it3l5cg4W
v1qm+teEi0ZPzNcwkGWad5rwSX/Hslk6dfEnQtAPH692IEJzlNfDBUsiDj77KIkvAV63el0YKwX3
3D5ibtcIdMwlVDke2N/EMfVOXN3zEIikTDDx7zQXroR4prV2BM1il5jR3aNCo5GkoQOIa5XGK71x
4DWJPPN5VawAYJMvDnLh4x1fFqxoUVvrVzFON2unNB8g8MJPSlr9g1huaiwYPrLmEr4m2IuVcxCx
7w79NsaVI9a6i5RUogUV3qJztjQTA85nyNYOBcq+695hYzDVdIW/VWMfOvymEpNzldTK7iDdzaZ1
1TwiTJ46QEoHpGoDAORUcTIQCVmGqqSiIpd1MvBVEwtWNfnqFpFsFwYdg1Ru3FC+EaGpfrtFkmNY
1Cdd0YDCj3XEcC4xLK0Su94VZ4sg9e7ECG7e81uh4aVhBR/MuzWJzUkefswlmUjceKBpw+aj/6KB
mTm5mzCJ57/0e5GQD4IbH2ikxlHm0ngEGqObxT8SBIORIdyubOijH9N76DGi0NJQyGWGK6PqrC67
Gmnf4Af0yEvTMrenO7XdqouEYkjprsAQ9FWHXD6KCzOIY/EA3HZ3U0tJyNzfpzqboBTwltnMiXXM
U8Do1k/MgD49f9OxnigaTomiKQij2ly29apLQUwfyKksaqwfCiA79zbpyyaB0I9Ho2wrrGSA7FXJ
T2gFw0ZajFQt2lIRWxaC9BfVpEzeqft3Jl33IBYdtd6ciF5HRZLQ4ye3LDWxebbNuiAmIEUtA19s
rmJh95Nqav4yg4IMOqVsquuqP3Ecjrtc7KA8MTDVxx6+JqP+EVs0I4kdDPsF9tFi+H78mxCY3K5p
hpYOV+4MxMp7IV8RvFQdOgDoHeo461DMu6+BmcXvrGEAZyr/MLB2zrc+JIF7I4nKmIJW4t6vXaSg
WLUCtmCkWm4t/smfIdBaZq1qiawFSNae6/5uRU6RrZUKyrjqM7GeqLQlZy6gHiQBF7DsUmWaOKAt
3KKPxcNjz/IGW+Trwyt/TEWNouK+hmqSFGWumVwP4oCi79akFb9MRYhw04iLLoj8/4nYh+FCbF4i
NFe2egSBY/qtzxfrdqJcaa8WAeKKnzSIWdise/D9uD2BLbKflGuWjv1Bj1bhYDm/Nf+AhAhyt3WA
XWSNbHO6Oz24F4O1RQUoI88GA4Bsc1dapJM91vLOhbYv4A60yBTrM7KIKDBREkxvkYHvLoF2A/c/
XXPyGOIyslLKzSEPZOsEVZ9zXlxQ5ayyqSnELCxCMK2itJh1azaiy2TQXi8ebRS2ISbGHMVtvF3l
qo8xttNNiM3zwJlql04+uLhcNaDKY+tRlAlk2B2bbD9CtIqgor/SLda+nHNKX6CjoDOZhYp91JVR
0PyujKymkxvDV28aygFw9axlArCOpr0bYQMLdlnrmOddSe0jq2fSeUdt6IiWNWdOCD8mQaEwTAMq
SHzt10EGGZ8OV98hKRe832nUSWMxDQ12fSABj1/a5c0Ata0a2qV1UmeAJuWjHsUkhENaUZGfcYuY
Slszkukwh5bTFjX0JkyqUNPUTTqOFmys35wsTIQgSJt3sN7RoUN48B3+15NjZP+UQOgU43ctvP1F
3Gta+RZAlxfLuiZZrvgP0mPeuqzmvIIPiATh18eZXAznwHbiMR7Yo8T7vlAXtxAF00btp5wa6TFI
kJiXsBEpW+nWd8D57TakCt/Gf6EUzhmlMCtfD1CbOBzf/BJcqyAON2mw1TlEIUFXHuQWVGKUh2vn
WbbN8Suol9n8jGVxVimK6oNSHfQN9aGRp5ke4e+viyHIqHj/gfD1jBVxU6lX19HuGbTEXxtj6plu
Em1JA7MayYz0L3Kf5QpZ7ZA7UK12zS1wTDbHP7RgqJb62WMUk7TJoMQBXpITSfZ11IeEsLchl2v1
W87jiBZruOSuF5LZCkqZt5tA7wwrX3+TRrEV0qqhkFaf+oyv13+ZcXocjH7A+K8wKqBgQBE4fjDe
d4J3/ed1aDdUNnIOheR9OW9lkHtoN7BX622emPGdZHDmdMBL7zikEa665453Sy3tFFvk6v1/uz/+
mqZ78X2zUEpBoL/oVNINqNTzV5Le0QH/dyRS81a1jHQJJiWnrXwdXSqX3SRYfy+yOEHakACJ31uQ
7JDxOmAVR/1HcNg2r0BTmyavTfbFzJMh/2uRScvZHzCFPv0Ede9+RWrVgt+7IkBTsS9cB9kMaG1S
2bkEuMEE9AnnMRomwsugzXAkKEKFZEXNx932r71ZUhIe38gbrGBJKOyMXp8yBnHpas8ZqDzF00tu
IwWxpZGztxG/tYQUR4YDNC2bPfyUqe6FzC+URuyuX8luNdTWxwv5fZA+I9hOhb/83Midxki1fBsR
jmEcpM2wi6+bisgVu5+yi1kdwqL573pUUu0S3KjezOa/8LwoajBSUZ4Rcliki1CuHcQhn1DkS8K3
iPTKJFrgwDmvthdHCGMiFve9Dq8JqWX1BbOl9STc//BmDLrirdaOp2qCpKzuziXwaSrsN75w1f+K
8dLX2S5cMOKPeb5HbGM1YjhFV1ce9abzRsojgyh1LHG/HwuBwhjRCcU/Dyg5uGwLmevlX+v/lDUc
/HdW8Mhx+f8jcbVXeS50GLXK/Euu0Kvv4VPErTp+DXfugfK1nEwuAfAbgpgMrsF0obfF+pZtgmQE
UEeC9/taXI9T1gJdKTBFEfIOWOfo4wpdVqHgLpxTbyE6r5LgkGkIu5rp1d0FmH+eesUPtr6KBRU/
t5gmHbNAHVTCVlb+rZs2g5BeVqndg3TXWtDqs9bt+5090HmA6dprpgVERZR1q5zKChis5vdLBvxv
giym+a9z28HtuEAUaAamaOh6pCCk3zToqv4iq47Kofe5WtkXW5iYrxSs/sxQjFQUt+0zO9gwROj0
TcqmHf6qT2BQ4o8zkIqH03oh8b9BGW0okgpuLUnVgLpjKlauHasSZll3qy9iKtw6TDf1EfVXK57J
QM9HPKgFcucRSdGzmsm+lOu6BgpRR9lV3QoEcOrWc0GSXgOamcLLE6Lek2TrMH72/cKhXPAJgs7T
pGK/XZWcergMXgr0QJuH+GYLqorYUKmxq1Yj4OIWXlwhBlxlkW4OhjClrX7yrHy3DbJw8qkMYteS
YOXw8WmnWt/Qg+PUnmuc4uv82r0HpNrrG/n6Jh9+98FRMApRvNyX4uy2meQ9iBYK9ZDqODNZpNq7
vvvzuEdZZxCHfiP4u8NgHzWF+ldn50IfdCzLmdYhZ9pPloHnwhNjQrP/eACt5tVGpo8NMBF7Efzz
4zO3k5kKXTIRGFqfznXw4iGBDgSdQ9bZ7erYwGr1oos3bUqpPzXgbXkX0OoQXLdQEXMjOBcSlxrH
d/jYQVJ17KoaAUUXAcX2QUCWkFwrlbTR/8iNqvTjdOGJZhqpU+S4FwKpIzI5oYI1iXvUytlgDcX7
vAFwHr1wPcWxBDuOM2SRfdI6CO+s2A4Cne9Sx2wqfWSnjkLirE3sDlzuVv6Z/RZLrE5mEKJe1iEc
7YtSxyRrzBrp4IuFrbRt+kYzI0hP+mTMnCTgYcJhYVROOWX3/Jbuycog3y5qKnLtZ/HybNv5Bjht
VcoiZocC0rJEXFWaxP8QYrwSusSA+xIpBazM8qp/mlwHbwSheXmqezTc7+SBCKym3Cg+A1ocUDu9
IKZzmMb6sOIeb+TFlHy/4CRqp9Jk042vLXNczeZIlUMpOGgGfJUQY/G5t1W9MEoL6SNg8N/NwWtE
RPAGgofP1r2Q8b2pPVO1JelQ3B/UFLP+Dg1trh9Tt+tteD2qGgKbJmWZ5xDls2dQKvhPYiSibFVC
Y5o9migzoN+vizpmNMpHOwgehfX+h1Or2mflllNAI+uGZDdAkNwXxUBZn5mnJTbapkPxzYSkzD4X
nZptXuyKNiMSdFfPNwzaj9JIUVNkzo8nCWGutbqgTFMX9XpXl3Za6lizury0plZy7Lia3zmWNkmP
PMr8wW2efBlPfzAsK3zMchSwPjWDa82b8a4AzwCTIQi8cBlbzafcF0FRMsgL/cHggLUMTxVejHGA
YyrqkZXacQbFVlez56rZXGjiF4xYmZE0JlkYIEMvmEGqE172JE2JSpduO7wn16rzyX6Jp77Bsatt
/ujmhqQKiMr3oBJ93oWF0kkx1seEj8yvi39V1mybxQfg6QyjSHMXCwR8GHVd/t2UAgpUtpm4byOW
6siviSVjsSxPmi68ILKW2zwJ7P0RZ9smbVVfXbm/jrYOjmzoeBxxSMCbX8dEdhy7KCQpoUQO6J53
y6X6ieP1swqoQHzuLXAJU1M378iazuw+alT/kti6qL7yFOcpq5jd2LBcBTUqDnqPIwc7LKmCpfyu
PvK3p51pJjO4ancPs4wrbEJC5TKJg+QJxILTqhuferyLFAlco2qqnbgMIdnBDr0giMJWgK5Li3Mj
nTqHACwkPlPa0+2KPINy6YNGZLIPKZT/BSh+wnTjd/lv5SbQxuikw3sxmaBJmAruZ8uWw/xfU4Pu
rRcgw7kv/5hFt0PXgJgqKbxYYDY9u16khEqHkKjIKr9FUoLLp3JxO0geoecCcdsyCwvuNlWHGlCv
uZcnpxqEM7V93ETm2W8a1eddM43Qq2dxy8afxRqJiVLjf/ZA1rTxd3VeHiYJQdulccwfyafkJbk7
rVqE373IWJYYDP1N/sT+dcEdg47BKENceRMWaSz8/dy5++7OM8paXUtwaHnIGatqEK3tTThxuDqI
A5QD8qLYN2g2X9Tp9cIrdqKHK/35ThZC2Y+e1yk/SYr43//4DG2F1JZn/cTYbQU1jcyPJlsxTRpD
ZzDZwl9sQ08VTh6LgS3MOecPaFeXFnPKMOhtV+4aEpjmKPQSXQvnNwsCTGpFDEeKIhLjR+GqMbCO
pTdiZ0Ww9bh1fvRsb8KFiXxLfNQZT4cTHqbYPmD/SQS4hJwzLAvbFMMFe3XdgmIfnd4QFbD+n67K
VLSvVvU5BfbtVabLD1RKk8LVZZBvDBZWUiXFEGEkJJbMuaT2wgkX0FNHIRXNDJgK7obLOFLf1Rw1
dzTfUoSb/AYyH/tkP17s2hfMz5PiGEkD1FqT7f3k0/E5UcEkqantrkKjLIyOjUlP7SdBzUJ0wKax
CgQ+rfKMZtMSpFV+/7SK0Gd6CRtaAhlW1CECVDcOqzvXj/XYQ/NumGkK6iyZ0E99qraeD7k8Y4XA
NduBJTCOWcfCsYVcrXcRXWbuGkxMFgeQ4Jxiu4HpXry64DZDc/4PI8qQT4fQI9WUufjwfODilKgQ
P28FSKOic49kUeF+BsT+iYVA4NMQlrwNJ9udZqg4oQNDJxiqq33c6g33dSqvTgJa0d3zUw0+4Xwk
MSSMlc44NArlhGsy63u8hHeu06r3SzHsct6IxAEbLdftRlHDF7yal9QSL7j+MGTgDlirdgQn7WH5
OdpcqQz9GM95j1AvdYrMH6qt1u1LJLD1nGMeStN72UeruU6ME35JWzL+QMWLid72mGSbgTiGBvTA
n5hYKOopfRDex8hIEH+KAVuy8n+Drcan/T1TWQ7Pn0QGmFb2ANUFMHcMF8Owj3lDa5NgWg8Dmdgu
VK1cxFxbU2ltNFmWAc15eGJnhKOr2PxijcmwIbMff+db4Lx3tfBXxKgc//OOKSFpJgcw6zbqU6rd
cuOvg4GIhUzegjm8UOjwJoK8bzkuFVjoSuTTpdso1FUZJ1409IBzAeXl4n6eDJJba63NEnl3APji
6bXM9mw9Xgaj8Eqxq2EWE3nnyLP+zj71Xa11OtzUPBu9MJrNnzIh0iH2oTqeSmgMTd34y0xevEzA
uNV0RusRr9Z27dHiw1h8N3FrHQhRPTvZVCrj0vYrujBw6yQpzD9Od5FkellRdfIClpn+fesehpO4
XScJ7wJJVcMKWuik9SBjPnUZtZLDFRVVLghU76TpLLah0xCJLgi7Me4KNsoFO+syDoZWatSxiY/v
gz3PIioy7iunB91a1XXZgDfuVqWPvirSqD3tHH0ZA2JP3h16MCBhMkW836Aq86SJiEKcggd1wutB
Zfp/5f8HOvCsCwX/Us0RjZUGeIDtPOqFrzWn2hXkZxf/Fu2yvP/Ljhv7UkUF6B4MyUb0KTRxy9eT
e9v0m8FMDHNHpgdaAJhbta+e8l9tXVdMuC2xfFGTtTezWP/aibTTCp3ijUkC/a39JkLXzWRCSpJ7
34RG/RC+sbUOHgupY2nxsjRzdeEVYpZm/x6b9lmiGrwvPcluGJr6x+rjbiFX/6an+zK3NDwTeTu0
CLgRQCkbyS49uRbTt6q99XSmwQERrsezapklYht5hG8b1n3Hh3BHnaENtZW5C5COVdLP0mxZi/us
FxbGUDqN016AoFXb/2bJjqTfbW1BB7P4aPByW8aeX0Ryua34m3HHzCewUcEX1v6cqCV5y0m/W/Az
AhTxfpm18prVeUNgv/k/dQ20A5M2sxsmUWHM9Cl5TdzoUbm4yQ4NFIZdD6CU1aimX0eNPB0kMZet
BZgztgNPkgzNv6/qsWoTs504Y1Y5Jk0QumeXdxz7MRe0ucX3DGV+6XSvwGhJPx/Gtsmi7e17We9w
y/qZ3l8tWHlLiEQUnRWA9Xr+Qsb95iNOz7yFv/ItHsKzQ0cAvGzsTHv7/cbari3VTFYsjTWU81rH
4S7NNcnBGjcoBAzMQZ7P6qH2ik7LSHqZvZ5sLZrdzWUMvm4wnp+GIZMF9K375OotXq+ALyJolBvE
eVbd1xoCvBIFEmQQHDTXZHfLv9m3UiSTnr11hBf8+il2Regsh30AHb7heKU+o9Mf5p/wd5CDJwtd
SQ4W05p3VjNE4J7ZiBaHDyVsdK9zAk1O3inxafley7Ne7D7JPlf0jrQGdgde6amOfcj5L3OEJpjH
5MQz/ZjmeM616SBuZzCA7ePPwm8Iz0nUQDTMThr7BaobZVgfkq5TZ/egZpxuZrm1CRX8TqJQwCAK
XA+przwSzDSKd5hkdqPEdMFA+hZMA7MpkMBsAbLXRkK7HrC1dEb2x8CyKvhps8+FLQCo2V3SWRgc
vUL8HDKAGdwCOJtPXhf8JWNQIirdg6XHG7LK/ZZbt1gUynV0dWf+mzpwFscltbCttLrRGNlDjQSx
JgWPCtl8dCJcgmyFs1Jk6ezr0kWzHHISloF7ElFyn/nZ4RAsN/Jv+ogcxZiVFY3qK+4LDpSWTlJa
3aJtw0YrK9tUcKVpefAGmsGCvgMzk3XHSpvwyXwh7zAmvvf4LaseYiJ0ag//4L0dWVbCFZFoA1+o
MEXr7QNiv+w82fSUhKgVYJR9cmtZZfbbz4v/KH5tH+urvYEHgqCuGJwLWkWF6tEfEazHsyHlgrqg
GccbCXCAVyDxYgemnodL14qGkQBRMP8MyOJid/NVHFWpNMQy2KwIhsSKSoMalnlOG4TAo7mS3kFE
Y6j5ozq12hElEDC/98K0D5AS/Laqm+/KHAm93ge0Pm3rnUfJJKRq725qXaBxGRuDv4C9e1jzHKbk
I+IqBcbHFWJFttZRLPp7SbOtGRaZutHS4TlVOcV/4Fy2j3eRNJWF/mgbuCzBOQ7dSqn8JznA+0o3
Z1x/iCqLiwhoD3z9Nz26Xd37RNSyV47rRX9a6u0xhEcRvUSX8TWbupvHmev/91hFVed/wmmQdWqX
FGXOwYE/BBp52uyESFRjyUr4l2obDxespO7Q/aU6DB3rDsjWmathHZg/NiKwWpv8aX1tVyWgzSHh
xS2sOLcwRrq+6T2QnC9gpMqIVAHCYakwjkuT2ODINuv+yFPr3AizbNlvvZ8Hdyc9HyH06vDKjoBw
SgA0hMVjwfhQoRJRtYECjWEuQfjRbL6v3OAn61EfHNENFb2St8j5ut9MWUOSszR8OmE2pFYSFGrq
pqXZUeXphLMST5aMd0fwMwutF5xEJf3V+HP28D8JqRlQc+SKVui34JA+jRXhDqUn42akc6Qn/xat
sVAtlz4xpJaPv1JzGS9p2MmCi5X097u3io1MadGo9Uu44iux4zy/PO0dnyDgJ0snmhbhYDDtMr3X
AENrV0ct/OQ85h4q2e2pl37Tabhp2yPRjmGlv3K2AxzeBNLWLEtt5sanmXRWY4QYZHiZJ2s2qB6b
A1d3DQzx82112V0M82g9fouh6CwM6xy0BDs7/XoCArKEbixbs/4pyjvJvTWAnBy6szd4YTgyeRKQ
iB5A5oswJn3kMcULfjIcVu9zWYyRX8xCixVyGZ15Pm0IGgqGLINxmKJPDqdUyjLJz3aBTNyq4heL
vYad7oOsdj/76Cz4zTB2xVa5dxjzJS0fQnVjkt09L4HvAtc/GsRBpvYyJBIN/ylhJUBO0+cxPXwc
M7RwYJCtkdUJm1L46ie/4us+Za/JmjjXqp1V6YKE1DJgWA8Wn9Ke2xze/V7e2lmnfDj+mkGv0Mx5
yz+VzCPokcbPvF+TkJl9QxDojXAqJdSsBB6nWYrrStwME3lT0bmmuPfBCla8Gqst952B6PL2JxRk
/aNW0dQA90BtxyuBbACffnxvk2IwxrLbOGV04mYaUlXClMSwsNyhEHyYDkMX8IFSNtafTds/wUxe
kCYpb8hnhFRLY8emqMYyhRGiqQ8FsEhadDV52G2l/hR5knyRhDllxr/joNerckYFQMQwfiT86N6R
frfoE7qbByWYss04ln9yM7+QEbzx3GcsY1C21/hwLXLuwZ1V6bxzsPiyybQ7s4w8KzALJ5KyQPBW
K97ook1oF4kzQI7C+vuOo/XUAFRweoAdOg7G6FmFcZq0GGZel85ZoYpGJbX2wb5KBt15ryiTkqgj
h848Nm7d8te0FtYsZ90OKj9svmvWhuCR1cuVgbtfkfue6Q7Yc+j/ui841NtA7CmJokPYmdNrVJzX
liAxlbL5KQ9rCi44LZBIAc01ntkrp/kWDUKOEfUNZSCIM3UWpK0b0z1POXB0P5MhnfwgXNrVkxiP
ISc+2gKD7jTshMqj9wfBwZ7/ayLc+NTSX9wzsr1J/DA4fLhKap6kpHUghxtCOtWKCTwTbHywDIVa
XIFbMM4632pnJciY8U0pjEKSCw3Fv3qV1bnq3RdmUeaHaK7mNjpe4EgEtx2xYkNI/TlIZRp5q3Xt
X+yK5E1ISwV3oKQQjiHAKW6znLwmt47ZKZcI0sKZRV5y80Z+cAS2QfrnkV7pUMaTFc9C9Chlbkcb
rFtbovrEBN2/xvf1QDFqf24QO/a7et4BbXSNsjbx/WXL16E1x+tYyOnSWn4QlsGzjqv0vB3BzyTY
yajInnAEqtF4bFKxAqbNeaW5zba63w3dSx3IbbB9snz2Sxtivox/NSGXQooVQiOLzZY0Aghv6qeM
BsARd7jTRnSV0OlPvQ+RGqt+RdaoboD3fbOrYntlIuPYPqWbOI8GaVuyzFJJuunDFTtONUOY1p4D
qp7QrRnG7IcoqnUtwOoieGTfXagO7taQ+XnLVrwXCkDoeG2is1HBU7hKfvS3Khc4NL+MHUew7jkf
QYvg3pmHTmYWbp2Irp28k9tszNAfgd6fh3qa4HkFll7pACsk9+TRWYC/fgWguqligac0w4Oi/bAV
bC1tVscWPXh87h7liyjbU0fFpw7JfwZNW6WyAS17NB5c73Izm9fry8+PR9NmAcGJ+eSATYpIZJcP
LDu3XPYcQb93RpJU92fKR02OGoNUFkYtThK3bHWV2IMf5A5L2J5jhR9B9OB3JntlETp1Gmy1vhch
g+jypip1j70JxUZZ0rV1n0y6A+rJCT2SMA693CxWYTiCQler7HG8NGHi8TVsoPzlXRw4HU8gnAOr
JClq9VBvri4LxyrvpabGVpYs35X/KmN/DCTB5iOWPq5QlG0X1u6gm5n/hcAVFT0Ld/P7BUz4VL4A
4R5Q+leWzeoAwS7bYIrqNgEl3rRvZTuh7Y4t2gprxZgZixF9nInvgMNjOnExSUBacfrD3mWck/xE
31a0o/ut1T1Lgl/EOaEoF8O0sFNM2M11nPvrXcyeY/wGCyUmO3Wm/Fx+wthBpkkVFB36bjxkMShJ
NoKikzeLInEE+Z5qSyhLkT81gd/AS8mMSwVcJ39/BLo/ClJnwGAggUKlGL+C/w3bpdsUOg1SXYbl
tv6PYowil/0vB+kfRo4MvKV8JT/dXVkutUjTav1HCvqTyAbhxbLbP8lY0wk960BBbxs8KVqoawQ9
aYbbOcshrYc/Ix1UNe9oUSAdcXqjYQBkZNpcOA8DgWNB2aK1G/38vcZhquL1bKrC46MMlsqnhX+h
WvkIX2/3QCUTqslpQPdG0+apEQCJRci1N7pAYTlkXohUQLxte8OoaQ/XfUipBDrk67EHtRE/27fh
onPnpkxL12M+zXjR7omflNilgrzkdGDin+m5/3fLLBc3o8HcrPmgWEkzDdAfccKanaqHRtxg9hf2
P+CMJ34B8iqPcfQhVM266B1sMRq++/VDA8qB5KNhdt1TLI5bRqqV02TTTjZ6zosZzazNRQxMzxA3
9VUaYm6xtat+UTx5rK/zKk6ovHYCbBLo5oDoDKuR88CqgnP91zUbqehUWhsbQwVOJUb+oBbFHcJ9
FYGodgAKUjEQvsmkZM2Me0/lnu99Dkm2SWyWkKtifu5jzXaxiKOP/ZlX7ME41rs0cgFTK6UZ/nQm
eAqGTsKW3UCn+wgQ2oWnC28tHvj/KqqzydByYEu4558f3M6yxNHGZIf3DbUELGdksfoyuh+gvgR1
gNjICz5pguVU90ZbhCkXItxTSHalyQDJ43pqNuDMvI3Ah174pfyc/Fu3zQwoRgkt6nDdY1ZJ31sG
GKTheETXCihqh5fQoBw/CQUt9+9VFrQBbLvOHUAMgUk2L4DLZ0AvVSbZ6Rj1Pzzyyb/BM+jbRGXD
cWvEn4yqMZ9rHKwKdOiOD4YSMC5tbk9JMrBDYXBWLj7G/ZrA8dQeuvdY2tOSYwPJN9WbAU6tMjoy
gii7G0Qg1zjLtbzRlo6Hk9NOieKZ+NRqHjZGxiDiqek8OdBhVZ7Z4AsfOzGjkkfVvyV1+hteBN3w
FQT7nmBdcyfMu7YbNsuAZmreJl8tXMPhP94cugG9+PdlbAyByeFP7TnTv2qt/le9fmPX4RojLxgR
cSLpwAz9L8Gc/kHYPDZgNQZHomyjVjGMakWlppCE1mwky6WRUUWHKy2vlMzN1sKfkDIbPn+gk3jI
CWQUWVBs2cdgHhdkQFO9AaxPu1h5ZhHPR6RAfyEkmCLDlCDKYkBAeNMM3vLfqu6m/U9vVmMKMFbW
aS51wDbqfJZli5Kbk7pAQAFGhmpRkBy1KIztmrODE3hlnsQc22tJYUPDBN/Blf7V5yQM4GGExrwc
p0zCEdrXAwNTvxnR2u/HUMK/q45vcEimxa6PIz4boqeKYVCvEzbrYgjxFOfubJ2U4jnkGJbSn6Yi
tPHDHN7iY+Q1qoBCQzpQD+oXvNejgY9uo4H+T3PYbItyAVX9DFAb3u83GR0oQQoSLilCDpCIHE0H
azubyjO6ifTX+8CRGrAeSRUt20ScukBTKyz3CRVHc9nsmyo1EYVqrIkqm111y8rIV6mhe24uHd6N
fSsmeyACEv1b7/u182+9u/omdqTFdppYgJhQUf9+hGRwiNQrRPxmMQ+nr3dsZ5Y8awyUZ44IQILQ
a1ITbz5vMqbJrf6yoH6N1lyIYmmXJ+YTMkA8pV8qf52zLqv4CQqJvrpjS/2+pXjIPGTxccOc9+/y
DdJuXwjXkUHfGUul9z8/AMxFPruL+sKQ6yYlRsv3K5w2lZVkuzRfCfDZVPYaPCbX41IVrUHkls+W
RPPwYyEgOZjH9nVDdefr/8Y0o5rlXJLxJKJUWbBQTwX6CxgKmuI0yT8O/HGNpKPlvtGpPFA8suJ7
Qq7wOZWuNWzY3o2WcpK/lNZVKFQCZHqaCRkaZLsbgnjfRtdNkSr1rAfauF28qTZ8ZmOczn4nBahV
bKBpVSvtUv6z9l7yizCD8b27dxaJ+bb12g7GaLhAPAx0vonVRkRxlb+iJM02htFfF/YlcScZVFpr
B5oVUCDy3YGkvUv+HkDY/+FEvM/eL5D78mo2I4jthzuq+1BTWCdS68ye/8pCWx+ThzkUmsQoTfBC
MjvpML6ZfdFAbnQYpmiogYR6MegPEi/j7QSCkNzYt0otCJKB5BdzgNnJATBODD4AK1DTEtKlZNLj
8CVi366BQHbd0wnzqZXyRExhC1AQS/w4E810cPU+tPkRnCsKun1PDpcerqLT5W6LWMJmqW4lNs3B
2wqveSpJLRsVqNFJNmqMkFLZ0JA94yun7v+X9f+5uj9S7qzVydavpItBKiIl+Y3jsqR0JvBNoc9e
tB5N5RbftyongAHjhMERAH05NMoYPuVpToULopmpOZw1VpTLmLPJptTgV8oTNAuECCWHgImNaCA7
97m+KXKKbvN2P/K0sj2dCw8EOWuuQXX2TU9skRjSO1S6dFCffktljYOOC+ZYEtAt2YZBsD2kTK10
Uy7w7olBXhZWsExPXXJ7OuxOs8vyM/PJknqEVkJjAkq3vANQA8a3VwxliYtAf/X5tzOrB69OmOyF
UMgdUQel//Yd7syM4Z3zV4jFSqArpd2IAMD1HwPEobsXH6ZHlYZdktVLwtnycjajWX48hmI4BznK
cD68ufunT+HTJNfUoDS2kVO4kUuQuuQS848Pllj4GnFIoj+DXNj4u3jhKhOE8+lmIX/lf9PPlmwl
vX9KUpfIyneetiyF2sxaClQVEX60tHrVYmQJtUnK8ZuZMSjdGgrGBu9/cIaW9Bgsx/p03/UX09/z
YX5USrhydt7BAXAcKsurPm77lqhE24wd8/INBYsrhf20XSSCjSuATpBWREuCoZxcp2vqrAXF29hi
ulIXRVoR60N1JE5J/HL1eE1ztZZrDX+fuK9GcOLiLUMWHyxke8NH78e1caNbrksYaWfK5qTu9Z0w
YD/9RshlcUhADZbjs5MHORFAmYH1z3awIWaN0sdAnFYOkkJgVl7Qs7NwqDZUEu3cr8gRlESzosvz
/aRIibGPUDEEdebo0MbygmbyLpJ80vwO2M94wBRFJmdHZ658LCffVG2qQks2NYqSvgtxR0/W7TEg
Vwd4624Dad2kPLFLpgaBt4tUckdSe/a7+Lhn7WPGTMPnofqJiHFygF5P1YQPlxBwA/iOPdRyk9+r
q7baXzuFFQF0gS1DbICUvQDcnEuN4TYw1dfF3tQ9a4CzXuJzszJfGquXczftgy+fSfk45GjvDLAO
5XeGocosr5RmmPf25zO8/M85geLqdLetTAPx0Ie94BfbZnBRbrcENua4/AkkLUsYQrVrK2ccHlRk
6O4po22+5OfJZBAcuCaz42QFKLwQysVlbf0npZCdabtqCPIoecTdrsJEKrQZWIX4r8H1fePKxHky
JYZtbXY43fbt8F3Npt5eFYOXmvTgoxNHdl7O38phImoBnBPrYDNeIk99kxyTriW/1Si9OzWpub8C
ywjg2m3M/bR/tgeRyGchZXA0SzXzfSpIo1h+inUxvb7V10zMSQxcZ1PXqONidNWxCbTfIbr584Ax
2Mdbt2jHXTPtQd6isNkE8EQH0GqMet4Ux6kvZFymLYCkb5kV6THuUlk2IuhsuAWzwmyBZW3dzm4s
55t5ePvF4Sjh0nboLdHctvk6DlMJAPtS5EPlots7JCY33VCHC/q9SkOkAAJhV3NienGjWQVJvHTI
xXonljKMs7YQ9GLxEGNPQqkAC9+PJ2KWETKh9NtnPO+OyOXXC4kLErDgZ0aoKQhScbyQYrU7MjVW
HzHCapBxkWRmlPV5IEd4N2uIBGJK8V/nYn3LwSe0cEUFSNmvlnOEnFfeaL6fgcPi7sE5OYiA3tye
pWrR0fz16zwoCwsx/2pK62aQBDmjfReq9D25cdkRhDwvRWwscy7UoTdWedD71MbC0fhuiL3Wqfcw
XHe6ohWfUpd0IMTggfbHIRcTs5o66WdbGsjJdM9GV9yH/AU0V+Pl/iduAwZ1aFrL9kTLW0HHsbnp
yTtAWFuf7/DsZln3TlWeUrPU+FhwSaZ3DKoJDJ0PWlmYpASOgfdCOJIrv1Xs1jdLtuR69yTr8guq
F3KTVhEPc4CqP3tr9vMC5ABbD32M3Zsc39bpfagWCcPTpfsrFI+1oStngspnq45x229NntyJg42m
VFZtSwewrSzclL0Mp7xpZP5yeYtwFo8hiat4xnwtz4sls4+fwWjvETbq6Ym8aTLtHgj0T0W/Wp83
qv3SBQiG4C44QO5adV66IFxjitMdb2W+XABfXFd34eTMwMQRo0HZFQ2eNO8oSgnx5n1XJ3ODgftI
xbRud5wXZXxWoe9IqDAFqV8EoI3SRK1qt/MwpEnDpvXo3BhPHwUi/0QrWCPNmWHFKLPJsVP+YVg1
2M+ixUimnrMF8ZZCdfPo+U0Sea+PEtzRA2327U3wIFzAbUl/3tlknXE2WqTL632xAze8Ix0zZa1u
vePMaBJs1Dt0W2MplKeBTNLHutOR8snNTfCFiLW64JkLvQmIt/phcWlS1tEz1zZj95YbwChQgGS6
7tyOfLjvMsGksN7gL7jrB+jR/8FB7f588Uo6mzpn8UfNNeB2Z7ubq4aimN1kQNERjoTTOBzlXcH4
knP3H0yty7C0A7V9A5VJhEgBLkd5NdwSNtvaXeJZ8PyTUJ0e3Gbic410YlcAMmxW8xAk4GwlvxA/
L4NFsbHTqPi5PDOyVpKihQvakxZ58XwK1LbwwnZvn7faH0ZHIfbfOXCsT8ArMHyCLqQ0djuDp17q
+M49jtxbAXhzleDv5DBh0W9RPvaRYR6AAjU8PMIQ2sgiwP2f1ZlG10czBnQQgsr8QzsHxwxcozTY
n9A8qwcYwpK2f0Y0x3jgMb20gpisKsEThrt+Cf+qd4mdGA7DRho0VpPixXvKkf+H6AD2OGHVjCsI
GnuZyyR3eWkp5gGrmGmevdS6EdUU0Pr/UWfFpe8WUfkRray2fGv2/h66iwmxoluIDw8fLFPryI8I
1f9AxZ0sAuIfHiIWl9PrXjtjeBFuZGlf0T+3RLfxbrjlFF4Qmh4F2jOIlPRnRlBWhCZzsIV0giOm
zi4q+a/7vU/yubaBiuXc1ch7fqLMBah+L8asbqk9HzXPYQotbuXiRWzpfMg3W6E7gyxmkevopZvd
uUPhXizjfW9tb2zP0zsMr+8n1zNOxY+KHpP0snHNkPk01wOn+6KQV8ofHcxMNi/KL2uXPamUV5MQ
M9KOm5aeSKug7pupGjSuRR0GpjEDH8LIfoiVh3at74r3rkmix51vFFBB0wX31m9fGFlDn4iZ/OFO
CYgjfwjrVXIF36BzRiI4j3wvYeEZZIj67ntf+zjbqXCNVMXhWaVH70n3oOAsP3Y7GXPPrPHkcFTT
sfOQ9c84ZvGRw/plFG8sBYrtbZVUv2+a7FypFeQdNx6F8DPMtP/QU07ehhdfpl6wSKDGoefDkt9U
c72Kh6EknVg1wl8sDCKmXzOPMQD49VSFqh85epkH3RjPbNpCHqFCvqzKPVRxHSMpIknkWFEauZdl
n60/cwYuv6JCw004w7FPBvWdqLjvbDac/sElJuaRoQXh5QW0cGJ8rfWHgvrEpTFRC0DeUkWU5Qi6
YKJ+F39IPZz8bYp0mAYV7W6WY4Hl8dwdQP88tRPSpKDDkIemNFCRifqAQIrkLzfKYjW5eqGzaE/N
W9FJbiLsI8QzWfIZUkt9tXO114r2YMt2j/bXJq6mkJDfAi3BBIP8eHvsIgykSMa9tBZNLwVNIrO9
oAyrOhvoF9xAe7NKe0V1T1gMwCKvfATlK6C8gpKMN3r1jdAc2xfdZwO61/Q5v9KlSCT4L4M1HMpw
jIgvv1eH2My6q5hnmCWf1ajaFFSfnJ9T8pEb4+UaK51Wtvz8AsBzAKmxc0Kua7ql8q00rp3Fv6bv
7faUXSXlNH0tKmkjCAXC1DP2vqi0JoHUzYBpoVJV39Yivc8rbQf/NisIFI/DQevYzvtQmagot8Xs
DFoAdUYfaqCPFuoqHH65IZQXN7iwYoEgBJkr44RSPrbScPcjxUKPd38hpTyS1iIUDVnv6jvP7XDG
30ukhgObWAq6qbnXtd0dqxOIEYzf+CBy0MJ/FE7xn6p/a3iP3lgXrEI4JxHCEV01t3vmXSfIEp4Z
NxOM2k2qXL+cgPfyG7hxknKk94C9TmkcFShF1sZAWbJL0vURqfjzGO/0K4Pm3ymEckSv+wavRZde
CuIwT5fpjJrhXKmvjXtZv1Z4dSZlehKpiBeba6AW4nMi6oueSmo5OueoQyvdiKPKat7s2Cb/5lxk
3xyiJwaV9K/MywD4d0CzAej+gskcg4t+3JL8oEKKS2OrvhdPGh5bqm7oWe4pDSlq19x6Y9g/lE/e
Wln5m6Ti7H0RHT1S73g/quuMW1NY2oF4lnW9T/J9GkrBuIS+o5RIY9i7rpXQngCdMtTX5s7G9a7p
LMhu1DcJgWnyGBvz5BPrLObgjx2CW38RY+ov1qTD9fqGzzgI/Hj0HZEKdkXz46gDbaSc5m5DoAUz
wFzF/O2NAxNVc9rdN0q6K5a/MDUacy364yiZgB1p9NhNiQ+gXX4fT/D+XhiE3M3+bI31vacqcb1U
PLIH7qHHsHHvbLR4eV1WZuMrwu+vsv1qcQe6XqEr5jF3jWc5KI1uhIKS5Ua8fVSRVk1DZZiMUR9s
NpgBPp+uqajN6hmTt3esFXp9XDj9WJCUbvsN9Tkl2Q1H++uokag7mMZOBaaHG2zAJ8guG6jLP9PG
AkiUa9MBE3mwmZEeocWs/VQXOXYIhUpj/LrWklmlxpIIa5IRA1kTvx7yY3ymv3Xt8YrEfXT+lZHH
08R59hl7nRoLX/cvkywHDTlnwVj9mTCmj+9wTpSyp5FsIeyqb/fdXS5b/JGcU18FYrTyOpU9aESr
LzInb6sZ9TTYcrU1w9D+ojUiHOiv5Vld9ScNHy+cf3hX1G8X/8PMcJVqGlmmVLTm10FzSFEF09Hj
IfcnnxJHCsRN0AUFI4ldqjz690ISB50EJZTUdRFCCGeh4QtfnO+sRBHQfUGVXkDAh/SX7QIg3K2H
AQobr8QNp2nGaDONhFXPZ5wstPgExeXckSXZfXrbwXNbKnHiU6sxN72BDPlnWnOMwPgyDgAAQePl
VuvNsXXVvWU3pnDxlT1XdtPl0oIJ9EfPmUvLQxfUn3da83o24iNdEyx8OamqHN/sfJ/YHIN+VyO5
Ok6DC5A6bU9De9eP+4hIH5gunm+BM0/qBFvDNPezlMIUbz/iCwQTlUCDRqwufAGGlHI1RtdElvf0
8N00qzESZu1GHZWuHQv/KniYzAi+wzyKkDCovzT2PeKw5ZVu7ZrBv6pWOW7dC5XCTKG0YVWGn2P/
bjQvgI2DXye2bZAPKj/y10x2+OJtztGig+uuz58MVdbqJalV6GmEzhkSbu3EynetD/IRpVsEI9CN
Njz8d595hKYfxMHpCRpccINj+73eaU6/GrU9g4eXcSqNo3RpazDwMI3HwhlM0Aq7G+ROW6KJdEw1
0Evn4SDguRwKur9oIj+7M+08R5Ws/i6red+dRz5Pzo90pTaTiF4mxzQR4QpcbaLMO7iF2xgS4mFt
LxmGi4y1LjZaEMvAbKu+K8YDoLEZOLwYJMI1R0BHxR3jP80rqY19kV2mTx57vWjHsqhN6xbyOGYu
oFglL07w1o7hrOhhdnAboIbXC5uDRwVoVT5v2VmwEWMSdX1QNYpE/SfWOBTu4n01kqO9mYCc+wnD
HxRtCASL01VWKMCNj8oYdZh0GN6mYLguajSkgN9pBx9ClyyNzcxQ9cNv57L+y+NHq3lV9G7EwMhO
eUJvfXR91jwWbtbPKWZRk/pxu3momLIoTC95ehWQQ0WF/nILPY6Ll642OyXk0gQqVTUoSuYiRaIs
4LUY+2I4w8ug0/c5ZhVf83G0LCmcJxrWy3Go69tmPCqf4tLv1qKVtI5TE4PNX7M72mYyIEQzETZ4
DvrrawtzOIh1U3M09CBblmfIyj+9sgbn36ZD3PmJkjX8go2whJZbRzp42xZNQEm/aOha8aecQi3X
DizvGg23KkW3gjtFjh1b0OcTRnQNbxsij1y7yuvygoRSkhEFWawMCk9wkqZ1YZW025JouoAMCRHH
SH7tzRmFuZpZ0s5iHAGEvFaEWUsTJ52c8+BvnlyPIF10Lu1siz3tP/SOiLEY/0yUGH0HcxGyqvHD
H+MW5JjnaaMmgREjV1gdTn9KvFuYw1UJ1KR6DY1E1h/Tqyb0zecbgHaTuXGL6z1XOSeuOROxb+PN
JiSOuwFq0dP3hP+guYnRruTk7678Uaxr8AtSLb8mJA9aoeDXQe7hBEVhdhS3a4EHaNN9gJsN7Xfm
09p7mTgfLxxxb2aeNLd8UJKst0PfEZIPUpDy1SPWwSf0vmdQ7leyRDOAH+Q8d4Deu3QStfA9gdYU
MYogR0We4hWmFS9dHrR9BpKyRbEDaIHheZgWxv0j2zVh/n6NvnldDWZHha11pI5SkXvVC2WfhCy/
N01WQr0Uz01jNIo0EomtSG3DE58e8Yxzj9UhxkDywXGrSccyDsdDFLR+K58jA6zQtoWFiunDRHmj
ZdtE2nHoZ+iVrxwF+0rkTIQaNroGZ7gDm2y7VLpDxzTVwqXaDc5VHuwb3Q/x/P6AmaDtmuoCTxg8
O6lQxop659wTQJ+VpHEgSjGRmgU5WzbdLGHIE+fGhH9BLBQoiFEvZ46oM2/0kE/hvNK4aXaX7QP+
4psQLC7Rxwlcm0JOnzUnauWlQqDRBwpWETN9yRNIIwiH+UrBjzyT78WYHaMDuHaq6bidJLaOc99s
5GjcPcB7iwdhiZt1RkIHPwt5YHNe2ESdsvnoJc6eJ7pt4Q0VXFoKApd2RIUnZx/SXerkfcIonglK
hlKqdoz5P+Tspr0jNQYxdGNjDgyu1NH7wyr6gSisAPsCkxcjmKPn1v+Yaj5T3fmrKJbzXKiHZSCi
OvWvVoYPXPJBpCT50pc2ET/N6lkI2jmTrNdjJ3TTDtXR7SzFMVsr58FFP9TYf8YSkL5hhmSbdSpw
+wxug8071L+T+kz6lTEuC7XQOqtFKFMI6cWnsPL+jjJLXF+eZqu4Zif8AzGS2ycpC9ft+3+8PXmE
iB9OPa4F7V2RKBr93uHFcnty8yvydo8W/OvVD5mpz+yFEnJo3IbCDZI058+QElmdzZbE/gWgFO8u
EPcl9t+vhIgd6Ftm03q74CpCoUy27qULN/GPiVPFDnq8rNBBIhqaAfoQE80TEXckNq/ix15mMZ/O
XJ4SxpBDZA26+Z6fpUhPXDIl9z4W3tL72X03MsHhVHMmDLFfH0hPacBHutJHrsyALSd36Sw/U9j7
32bI3aoiGkfbxpUTmTqEqdQKqoRaioga7qRuU+vUYkF5fySGn+cFg3glpqDEzit19OKuDJYddVuJ
qI50wpVU9sh1X3t7oVfDnL5hqM+NYSZ+cqg7K2RXdjICgMxRwqAOGJFVghJv91o9UHrCHtxaUhnF
TOjlsQ1N6U7nuVJQZz7jhrQp2ZBIu5XUIFZph3NRKm7UJ/vi9F5EzcoFhi6VCkgjqDTz2A+trEYR
OB2pu14uq8KVnZGx4vHZAzNbp0JcWA4Zii0HhryXCBzvGj14S/qJh6CR9JoOabTMEDW2iy1pR1Bu
57skBs0c3baKXO6+Lf/6W5/BBG9qZUimHErIjK6u+NUgIPcjJd0cDWURaEW+OPFA+3zcNlC7aRii
Ubz0TSxHW0s8K+4cxX4jufD9r7pExLDI9Zgozu7pb0dHWIegwKLasTUi4EjNBdGjLgIFMYQQijO0
hzugqIi3kh2Qt4Sq+i9Pnp07WBLr3Lg+ChUmt9FbojUB8mZLwZFfXZfqkAAHEn1acfdkUz0zZDPG
mdWBKJ0kd+7f0IUJgZGemSVgcakFSD5QLgJvTFn0dwjlMlSmU6ZBhFbiWiiPdX7Y2eyvUSMtBixF
XmL+9/8rTKifXoOMpW7GjkUoVlzgJvwrIWdIlGrs8sNbWpnEBtPNsTniQQP+JDY0rxxnQimEyrLo
VORY1ljif09ubFG7Zzm2SMlyIO0EeYy9hWIw/LHgm3qp2Q7wGhWK7J4wAdt9C1GHbUfhe5R8YonM
bgMOjGkQlEgcinUfr/b86xQYLCvpQf9tG+4rZIsIeqFBrDP6PaJbHipOW5CG1sA/3QkyDAIz0gtE
Spqw1dXhCJckumSsxE6k1xt/yUbY2f0FrUAO/xXYVwZiRWb9QYDu82eTtwTLNLlIIFV+1u13RgQm
sYcafU3XddziZINwVUVyh7fWSLxxLi5GSNPQQGtGzX3LofiAgh4tYcL6ucaIPLP45iKCH6PK0hOu
ZwuwnKocKkOdH3WGACVitA5K4TOAyqP9g60XOw6e3daFiznjFjDPtZSUSiPIyQ0l8TJ2mdKnXur3
3c/Mpm5aEvJrMWZp/4IfSVDrvYvVIQE90UJvwMHF9ukNetfBtFvr/A6OmZ8yxyV33Lns2edvShzG
LHUmz118k5DbcX36scGEHY5MWZvHrDQdh0EbajOD0Y1GatvIo5NBYzfe0IpRvVD+G9Vy5AVDJTQS
ClzYEVUSxOhCjBPMnk5hXZWKD06i/9MxkRaK7mdZWKHSdPxLb+1f5VMmvPtab59vf+xK4k6KbNX7
FV4ygBR64qZ9e6jSP3RUK8kUYcQF327XXOkR32IKrjn8ES6FTNmBh58JJ0BISB0nWtJJPbsrPxAR
M78hTnj0wO8HCopJnpes1hoxrVBF4PEQQoAsF/x1w4/moQ8YVXb+NvA55nU4yJ0bQKx7FkYz9Ztd
4e2a9XbH6nCi0rpS4Og/EQzNT/9MH/vv2jNcw8uMRK9+7syECmwjzVSnH6pvqMMt2hbwjVa4ALeI
vH79pdiLP/Vy9aJRF6/e3AE0tuvqRcP33EFCUFJmkng8vQfcn5Y1Uq6e2UmuzRSbUGWkDl8LL0bS
QcxUVCQnXgYMK6FQTljQMOubAxriIpha76tgcPj6iUM/nV+JOALlGAy8TLcmBVNqF/8eMny4NC8j
sa6Kp3RkTYR5kPkzP1MkENm8VRfdDGujTsLqD83MqIUTKMI6GRSwCo8eiRPn7D257nIUpMF3VH1v
AEj3uT8MwuaIymJ9idHkUz04mRDu47nZQ8Av5ninlDPoNzkwpCusfNUmCHAjhx1JP+2eYVo+fkcN
WOTmiGWLaUoeETQ+DC83jXNcMFuM5I2Yf2qvnZCFl/tV6iJEHKdQm+cO/5wxFxQPmY+IeRjGF44I
FZShoBAbmgIV/HooidNnU4RPqOeRVHNLoKwf3cFf/zHfphhPME14OuO+vDUnohuL3XHllO1DOIhE
r8P9F+/ioKsE6NdVh+JyvwmU6sowlxAMxXoTSfRCwDEdzcVWaS+5oK8+0moMv1QM8OA1aOD0/rnq
fv1GjC1SqpXsh1c/OGXVhMexVJSbHBeyuGuk/PoBmYLe3+W3MA4G+JxpOJHxyU/CU85fvSXOrEbK
GMKLOn64UJ/7sw56SorUin1rSMNS912XVx2ASGC3zHc8hOEMWHl9/59Y3msqHv+KYiwNTWJglDVd
c9wemqeMqG3HH3YP6ocdmBB3AQ5OQfX5eOVjii6EDTvUU97ymBKwBtHNzF6Cup5cjyr7QFNYl8UR
PE522khTFU7Zqv17xesP3fGgqEWb63Bv6tkK3THB5XeHfZxSEQ0u13GkGtG+mSUDAs2km0SyHUKF
HVOlS6/qQ6XsnneGSu/3QfK5GSs/4WGIJiGCk1M6PXPdqjIXlyjwRNXeKyJNo3XDDYDId8uwIJkh
AejHutB7bqPp9z+MEH06m+VJF40WvQMwZqmnmD7JAqFtu4tgMFESKgKDDLELTOgj2yW3fdmptkOQ
oAEG0jrfZ7xhpy0pU9qBu4MhVVeM3P0/UFy2tf1YM92M3KcyW4+XcFR/NENX3jZCywRH+Htt4i9C
Xx1WZEtB04eouG2Xvo8p9hqgC03WM5X32/40cJKDPVrhTREUDp9xkTpEpSIODrhMwR7IHBOmSe+9
Q/TrWkZL9FEiL+7BComn8HAxp8+8IVXeRbDVFN8aX3YuH70ZXDRSHMxfft8MVXFOViBgaq13Nd5Q
p5Z/cTvZSvKP7CI5gvEy5NymHgGU+pXmCKpduQppDacHjPMo/b83e5YSVSvN4/XievXfNV1WzYLv
vPZCll5Igisc91W7K49eTGbCy/RtYcdkT7qfErwvVzyFYmo8gy91PkL/wTRQ3hi4G2RvhCH2D2b4
es6XMi5V0W6YkbzhDixn7qHjQEKJZKLRjs1veBoBRsULOKi0GKFpIcKUbFaXTfoPZuAhBrlnP9/r
3mccjAWRCylDOVeExbZYC0dYxeUHRwkzIZstiKJNbXR/yiCme8naZCo0+MJXO41tQJA6Wd3V7Rrj
zX6/A4v5Fr2J15YlEc8/+QLj9NaXKuz1CXZorr+kROpqTc4P+csKZV0VZSgn+FXYeBDVjMBOD6xt
se0quATpPr/L7Pj3UbHzoWh2tv8ZqieyM+dwBYqiaCVPnFmiGKdgxW4/1Z4a4rk3FEU0UYDFNplO
rqr5vm6h64VN0qJsdIETh4cvS1EON1Bklcp1TU1gKdmCECHboCmaxBAObS+fgN1/QwxRXAU2Ax9y
vuMjTTGbPmbFuA/4L0Jcak6mntCP0L1pjY6GAIaPQ1qChP/94Kc4Xj8JFAwbQ9RcL2aPV8LN1goz
rQxwHLzYf7v2sS60mSlwcNDe5Kid5igPpBLrNfsNfCyL7u9S/d2Hizlj+YVORavjGKjjPsYGfJd4
3Hkb7pLyZMJuS0RMSw1vixEwiIVLcRCviOsB6BB3y0mU28larHy50EACnrXtPVk78RsqKPdnyIEi
pr/PiyRXO5/MDn3PtimSAyCoEcaeOpo4p19OsQE9u6CrOm/IUzQBC6eQBjOZA/Nom8N/ph5FYG2/
rClLqi1Uo9upnbyXTCdkVa5NfNICW0m2stIcnRCRXJcLXt01xj9J5RRXmidyTstDmRllK9iNns2s
1EE3fjDr47fOA+y/aCVG1r/g10aptjENRIwHGOtFT9vs2BvZ2LWJWPMggvqnKDhj03FODCzB9FST
6wl/rjlMzn4HgA6QvbyTqg2+2/D1NiaUuiET2RVLa1GRFgipghtZ5LRNC/oIm7gjKzu/kgWdoa5b
TCK6JHy43H2lhJhITjPSEyJx7iPHa3bSnL+wdgqi58NyRsDNuv8wJZfMVe3DW3yuBWEUvcMtgVbv
QdBErXf8sPycRbOxzDDxUK/WHsRsxwkp8hK0etMznV/bAlcbnrdN7kzIDOGRx93N/+hxTakD+3zA
abLbJNt2WsBiYS/ujDmMjwPcOpylpyYjGRyXFw8EwhTExbmxUSzRnC5VNw50pwy90hwalL2gBcfx
6MZ4VArGzqLli0DJqNKwpXh+1zVBJhb6nUwb+BJrAmwP5W0YLfTI1tkPK7Loc3QwLBYKWPGHHmnY
mFlEtLONPdgXUo2FgkiTFTyk5obFAdOFenFh0bBUMGWEBJlcVYMq6H924dIUqEW6tZFRHvwZU5Xf
ZiLuXm9xhQHQYtV3+KN0DfnDS/t+8Zt7WYyIqwkwAmdG7Pqq9Bly9SrOxSQFIftARn87kcA5lzWn
KfVvOMVHJZZp3GRNmkCd0Wo/7IjLBoEkStXXAZ8kmvl+43ouw1iF5UsFyAGUAy5Bc/3MzY1ON8tW
+hsCJWwOAuDyHvzo02GU4GxZvZiT/cPZyHsj/p5UunUGvnSNq69Q0fjL9F09tkySqjsWpTrGdh1v
9zcWQcG6Ls90CkNKzFbkVZUNpiJ2NHCrf7pjBmshTTxVlCLobShM+upZapzmMRNfyi1DkqIJu9Ki
wqrOlGQbokn91Gg5Nbeh9V3nIuK6LJseUR11aoxZsJvMebY9ETyIrHlkvrimSw+q4wkhxekXOsM0
X2PYVkNErSC/MIvQvcArZEGifWEHgZZjhiUS5QHdXWcl84KUIXk84sB1Ae0RKZ+sC/hDSgazpp67
6Yhhb84K0Cw6nI022Oe03tDku4rs2Z45dgJiNdW+GmFH/245ltao+30AOeensJPR4M2E//9EEolx
YX0NPM7iqFGMbYJgn27+PCEzEwyPXdm6UZ+zWFnwQ04u6gSpUtfcJaB17khwX9C2Pb7VLfp56Df+
mn0tf6CqLFKXnnS+vZ/CGImI83ypZpsR19vPjuG/KDumnkzkcUFmOctcKCQqusAJa83WbZcl3lbh
aLCgvYkvSGFKf/WQbBJUJyJE3MfHcDu6RHDj9EbCV/LjcAqwQM213JdpR+hNlwtl8hXzdhT3nJfl
9iWzOG+Qgi9M+Rp8Qrcsa5yu2e7qR4prb7QOvpSYT0YGD+1/3qmsMOpR6dQVx35uKut3X8nz4RSW
+PacR2q/O3TIGQ5YyHb+V180Fl09+xFvriWsGSzyGtGjF99frmxzEXKdZ0w+0FEDIH3Fqi10V4V8
dRNvl+BBQ6oenYQ1cZGMzfGmHEEHg3jrds8XG0wpPdgWGADjKvwh87+mG6DHzUy1hee6QY92QYoI
3buJXkBVNGihkMRbqZPINjrqFIk2i63BNItALsdCDT1rP7Uo5vRBDTe4d6PKf56mSSda93aiRSTK
+5RBqo4YVoPy3fo9LqpaBcF5v29ToSmTXnjCxcwjhaAYDkKCcA/N5hpH5kq6uKj4kPTV/mgp2VZ5
ePSvp3epsEB5JHdN0BXHCy6xc1NVONNsXuL3zbuDE6XceaKTcIRJqDfrfudZSLLF/Km9fSkC78mu
ejcHs79MX2uk7bWMT53yPHdrQAyoOMYIkUzaTNMhrGBvnxmvwjUW5OPvpYGIwru76O83xXCjekoI
7KIi38NLKpuV53fwojiJLPT7YhNeQW9heZUHv0CgBJQthzdQumgYNaVF+a4NCqR02CahsCqB/HyG
4JQ+P+hTL9Qv8uF/YbjPIoFmxe8QmrBvx+2bLhnxSnCBx/SXVstEi8Q5Efz0MmtmDdfbVpyUBosf
mVtCe7aDiJs0j02uztMG3Q0OG8/XJoSFKfTNDKEhva7ccc/P1fwMTNMKgYMn+vLtJwqsVrNaC/Z9
vEkU9rvkZB6d3A6L69uCFOJMiFgDHupnX3/K50O8bsKtHNm3feM8xYaSuGzVn3fonIvTtMjFErtx
Twpq4EnoOFCTZKztQPMyqx8VfpzOyHXEKsqOlhBycsiftDZQ6vjrIfT2AHh3yISUJHFLEh8vnlu0
x7WYKXbWXnvgSP4NJzn3zNgQYbPHWM+PLtuDzEN2K06jLZq5ZrfA7Vy6yDZ/cX7ED00uVpKBOEp6
4sGMXHbLm1pSz1B9DVY/6W6dA78tWvju/0P4Lw6NFmtkHgLae2qSQwZrvWOXzF+mB7NPPuTkiNIm
LE8xGVfQi2yJMWZOAE8WTMTDwAjNAZGedZK5dom8Bfwe9X95CeOpAEnzdBTbaRa+ZCNURoY4R/Au
tASxzNGD69F9j7UMy4qqJ/KVBPzMbjXdEcRYwaKhcdZKVq2YqFuQkzhCACiKCBTt6MTa8NA6wQMV
xcY5Am1evskRm5EpYpoby3l7Ola+rFaPB9NV2mNFnh+YTL3HEeHEH1uiMe+jmb/9av34f+eL3d0e
pxH7LbfuBsSR5fkbdiB45755QZC7ZXdwy7vZDcJNcX3Oxpw7UNwDfrztVusJeOPM/KDzpyRHELcn
X33FaRyWTPO1QkdnSVhyRUUa8Hcl6RJ9bSJHhZN6+aF1IRElhrHfD0JBK2XErwPQpSry4RXnQ6t7
4pNGaeQw9Y3iRrf+0ih2MN/hUH1yw2bQNCf0Xqn6xsT78NKSqKz1GYho7L36Pwv/z3+3N/qIa999
txXKG3nOPyOkRIJaBctZH2RdYMQRkUfXqudCjFexODhp0yG6NDAWF4raZl6D6VYkrlHzC1R4gna5
E3Zu0vVkgX+5+AEVH8uDtBbR8dY7ISrATHGRvdfJh8vftpOrK3EUKD3XchjXlQt0ARTUqUjy9v1f
87/utjIRp+RpvHCcrdql/XQRi/bRAJBFQyM15+5WvlxZiV/tkAlU8S06L+aX7CQQA6MoSWW/y4FY
i/7fCNBuhmV+cha135rpupG3ua4wMI1p9EhPZOL1hB3yJwNhMYLLOXWkPzBynEWIaA/Mw56o+QTL
82DSsRly/J5bVaFio4mrf3WL5HFS1DslzkuIzfU/ZzucqLCU7+Zjdq0ycFXOgooMS8iFFi55zzva
Ru8T0yM8hU4IduaXRwW9o2J9YN3C+vWIBQ6TkRCiPuVe39qihDVNDmgueneyBmAbWjMQqrVrHTJM
1My6X63PKJQWb6ckWv+kYtSmm5ZY/QQu/FLxYuvPFPd+1nx8IUhYBgBSQTQAoe8GGDf5HvBSDjZP
UWYw4RviOaezn+eeYuvy2wDxyx08bRY1/JC9zF4pw42BorBGO1/HdD8AOJAdNUf8hXuspi5yb3SG
wDj/TTF8axH8rVGJ3UmBvy7X8KDlwT5V7HphGTCvDqePx6ZLa70h8RoLxXZYKDhcWMOunlFjH2UX
RGHoWkCsCrV/nqkdoS1ZcWVT9+zcNqit4fiK4IzqL9ntro/OJeNHB1N80LUsMLENGXzm+XKeHoiA
59M6MdK594Ik2chk99BP5Fb0C34lGG+ux1n2vaYNNqiUgufZC97I+Wlrb6vTT/jkTjHqHMbXRhaG
w9r76ecj571z22+XBjIwfK1sOUaK+GEF6KI0MhBgrq/Zbtl9I5BPvtVvAMSzZy2DVOCbZgBPNhQt
stUwTATaqvIgBfTelRS2p8ivCp1TiK094YHw5Zluyq59F473Qmk474Bfy6hmukZ0oVD4CWRScXU0
VyBmrELcLCR0FZjb6rXcv6OVjz2Dt5Xh+60umF4xDEfPNEuCxiNt5piy6nPjVUDIGWrv/iwF6gKw
NAZ0MMvjbn9774/2D/Dnq0lkdLzId+2/wItHzl+ADVF4pfHsEl/ECrKyQRBVbLXeX7aY1Y9rKIHS
ikMfysT6jzBsmaXwNteXNLg/lU7ug101s0hlcLg2kCe1/7Tq6y88nzUkDgHASdoEhhvJw1/or6lF
9t+5MgyiYg7jZN0eBx5TriW3rT1La+TAxCkUO23YZQq0+Hh927y61X2tGyLeM4oTxvUQkLwRUirF
kZppIwH3neZnjNjcg9DTssvNoG38v66+jntc38v4+rzPG8W3yNgRMGDEYxyy0sIvyczVBRVTWgJZ
9xpPZrwcnaxB8NOQUtzVHitoz9uD7UJ8n7PGs/fQEa036auzQ9ypZNHkH4TG/yLocdmYFqtZzE/M
ioD6MzH8ZcD1XZQV2vHUG6pskNpV/jQqlNDI/+q8fLMMgQlWckKJlub9c/x52oFApn3rHMY3E/vr
DOUkXT8avVHQWiiJrgZIftifL9jnj7Bsdq0hbRHJXI6kYMIaQ5iCad8gEi7Km1T87DNHwe6282lz
/Qb+j3l0yspDjJ26aohWp0ztuDjcD0drumIqSo+jWqV7xHcfcxqivQm1M/c6pzwOrwTsc8zR9r10
xM93AaIgimRU2MLBR8VVL14lMoh7PMEUtsenGWJyHY1an+LAgUQTEwiY3ji6xOZ84fg/cNZvEsBV
vM3mrL/CAyLOkBgBxlnNUmIaxfNyTWSa1pVVsvuZ7Q+wJIIDfudFFHnZIO/k8duy/3HPk9wa8UPP
Tg5wvOimd+t01gP1Y7RrrqUAfgwhchx5nXpynOReWLqoVca0qvnR4um/IGISkN4eInrLxg21NoZG
2qpnHvTrlkSPbXuI3f6tnNPdQKOQbd/AiRdhBGS0umlv47MctJumVmD8wF1EaFZ6iIGqpq6BG5Y7
HzqpPLNJDI/rmFRmspPGWcUnzkUNSGNuFQ3xbRDODQ3WCwU+OHMmp4gaFuMR6YipSXPa8FJUiPy2
OPJf4JF3V/3WyABHO4BHSmCMuib0YMFaD43Q/B4Fm/hsTj3JXPBaWHZ1/Ee3AatEmxJjyFcNH+4q
bGg5Kpn61ht8wNxfO0KkKfW5KPaf+R7JtTNkpp1dSKaJA3+QCh6ps/BTgRt8oD0OinXSBuznJb7u
U5akSUblYj0lPZsyBowuNZu3T5rHURX8H+dG8CSK1qpcoA57vaUDhG8ZBbeJtSgeKjB1T22njr+e
GNAyERciY+ucZn+5zXfZMKX2Aw4TQNGUBfDsQTm/Ek0WW2UOmSZwAOS7920wmyP821x5hgoa4mN3
XiX1VJwl8t0H1xYOZ+ofCUDrUb/LmIlXmJA3VDUW7a58QpqKUHV7FMzTmA8/gT8Q6avTVJjWHztZ
iD9188Di4vvbVvKttLxT7lJeyNVoOWJ52hc4apNWrjSikGiKSWIHXpDOgl0FWlWwiQxSJwKLK9CZ
KvyfVdbtRxFNk4WSjqn/Qi/lRq8GUr3trfdqN7GlwapP0EvMHJG8W6V6NepU5kDe1UMStBfFjmzb
xrs2KjL4mz3QMEvW6qr1FOWu2Cp2Cyv/j+eQYzL9T7fa2jdRGt73Fb2aAzqQ0OW7CmOMar4Gh6qs
G6CbNHiq0KfgQ4Q81YkehqTBMykKDoDqeZ8UZF1frTpoKqajAro2s2Lo7NilKTNeUAwggIZFcq44
XhJg+kzufgWCkc8YD7btv808E83BEhB4tqbOOyj0/4fZ7rZ4opbMjSPwPvw9fzTIx42VwCEz4iWv
JsM9JNrIjJEIMNrjoEJCoBDHFeZBeRsiWKSKRzxYLsk12xQ+6d9m2Fl+z2ZrdEh9VKYPU4MrBgFj
nRCujvD+AcDRH6rbVTWG2oiIxxMu0+Y91EY4wVuqfdSYgV1KU2qCnZPOUQFIZis0cV+bL/jnZ8fe
PAHej3xQU8MLpRPli3l2KaKceKvfI1n+pYKTb48RNiCiI5GN17J7CNQEcs3M+VNBqcpi/n+zmN4m
pljIzWFsyXYpXPpCo05gEJ0nOaZK4DKPD8LwrjRlAQ8v+sOQyJd/FvSjKK+GAcTlmMRj3LRr/yGS
OX+PFF1XpayOGt9OsfX1DQfbXzmVqLU1zFYJAqK8jxjx//AQooWb1t3eVZ0KqLvG/pf6oMRffU2I
C0M3xPU5osvZ17l2YRoz8wu3Nyp3QXoAtTZTPrCEpZVs1wD5kzdcSXenfToGXuhejTRhTL3FikfV
NVpvShD2Wl7edTbGOm9UV4A12BAhluMgNh0cqQWxMaVEjKdbxPr4PrCH7TpoyeSbtYI6aXK0cVmm
vSKLTtXe1DJd5f6Y+w0RQXxSr8gSdOkM26FA0DKmRS0OQC+q5knaHMyn9rNQRT6ftOR9xY+XZ6Ku
KQIhhcTcQHHRPGHG1rVMnQfySmDXdZJxdZL3MSee5ZE877nllgV4gFIsHqp/cYDCFVYWQHO348Ae
FJfXn0zxF4qfIzCQ/dNEfU8dZ13GcnhwAIJtEwP8yCcJQFqpV98Pf4fojm6oBC/jV8hkN59Nx7L3
tIUtgOX+8mzjdlOu04wtzdkZNCQcY+E/Nmt5GcLsvO29y3sHARNpxIfF0JR3666hMNMtbfHGejYv
R1ZrqmRXikYQ9MK0ZP/9k3BaUngwZqvnAaImZbtzvwCkFzJbUs8TY7/iAuCHvvOji6AfOAnQlb3O
3u1ZcVc8Q3455dL/yLAnGWDh1cnJ1vofa8+sBOD1yMcIFDRI6+GyQcl/eh2NX/rzlCFapPqYEJUL
42K70CJ/gctmuTV50AJIhR5tQz+D8c6zYpp9YhiBMnlBAASTjrDl3W09TOOcxpYqngcMs/VJauHi
3PrKG8Q9icz7wMpy/DFdZnYydWUQwYT/uPmoqKPUCX2RVdtYYOyyHwWz5riS0+pHj3/mDHnF+0yN
ZF4QcOqWTcSZS3oyTtxC/Yq5bNo7BcfWe+ggEdOqOidJ17DgZWs28D3HnZxXICXP+JpR4xeEhfbT
PBKpLhgsxIRD3mkbdwEdktKihBDqg55iQSFE3TLlZ/AFl0RrM9z2zcF/1KjLwo/MIYMJyjA1qvt0
Ka1Aiw0ykO9/YOa+PBWd/BMWoBn/jH4Q4r5HeLljqiyA7LZyBdcr/Ez16M+5BpFvCHrMEtKR7DQe
LLqhgS9pnaQenLofsC4b8HVzBwthiyPhi6PIDzRTRcQ1ElRuppNq+A7Yxs93cysGITS9+7TnG3mC
5ygx3351gVGLMfNlSLsBaLzIsvYft3lkzVE2pPw7f24M0lNrvRGtiqx3Z0m93wA0g30UhL/KcNo2
gvwfcVCFuRquKN62jw/8j9CRPYaKZd2MstDaZlyANEr6uV6U1PjXvjFHNZflIUn1l+Smouff3ltU
+g9PLcT4RhDEroi2GYwgF4poVFNbakeXP/2UR4WrbEGQhwgdOhMZ5VwVwHV10oEm8ZNwj3zk3bIn
PqgC/SELP89QulfHcnjlUixuOIYm5jTt7O27f1qk26/7RugvHBEi74CvlLyIGGTlDzlQFkMEhZHY
/Lu01Sk/tObKjetZemYCOMvyQKR/tJXOdXnOd8yJv2lLLrJCDpbrZso02HZUfj/xTNkfFigsUOXM
yJLlsvwOaxflr5ZzcTmgdWE9dwQ/5DMfRhr5b3ctnDaxXECiNFrmy0shVBaJabPb12UO5l9wTei8
1B8GbA7lP+LYlsHuV3WwR9zaqdy1+bUr7b44CfGB7jK0U/KAdqcNt6ZKSzuiBDMBsEyf1yf7zgTR
jR1bqKkGmCN9b/viDaZyK33gm4O/aBcwoDY8Nm9CNcfZ3P9xNjUXdZFVqRkNSh3mj4sGdqb5dUiU
qsQ01kA8Q+MuJBr8LOaM7qX6itsT/4KGhobHnJXdL59WGvV3m1Ev8sGp+N6YvvqKQJ95Zu8NTI03
YN05gmU3AFCNLlMbomdfhznmM5aovdrBozXys1GWAiSogSTfLGrIekygliWpUCzXCzdA4ijmVdYC
ahCs6DZgCo+PvSIWnX3HPUD0rQJRJHQr/rJp+tBOl0sGxeVns9SJCcsMffKqmVPJ2W2GFwZrTui0
dViEs/vp+1ieEGJBHP20nhwPo8lwlrCD8IZQuXUGjJ2QI90Nu5BSE/WPa2rwgxdfQSIx0TqiZTyl
hgx/G639CeT0X8hvNgF3oIDcR7QubX1Nde5pIcKjmSr/sh3897z+Llm0MkPTWYI7T/qV9rtTMrW6
c/3jgz2+igUSio96AeN1ReiuNuYLo9MN1wU9DBIzIQzt5Q7xZAE48lx4NGDvtAw0WDDUsDt9cAxS
Brw/rO76r3dF/XNMmy46ODXr6XR0gLhB33cQGIdcBCDzkB5YX11si+ic7gUDOwLhL9G0IIwEGBIj
Tg5aGPMYJWCDNEB4dGId2faaz11k0cw83FOFeLdhrHWrlxFQ1ZFfvBNzqMa9FQGCPpxPfV/Cy8Gq
oPW6DlZxoSpaWUHHUKVMC+w5cHGpjZPV3zwD3tdgTEQc5J+XW3FFe7HLK2BpkGrvUPWJuYshzLUd
/6KrHFzDMgVaYlvXYf92K6YqG/LQqMMALSUzJ+xeKQazLLV0voaXQ3pBHcsLCw0F2LyHPdVArJI2
FGSOWcIbK4XQGyGc88s5huSD3F6b9HqjXqEkEm7gBtyjS2zyANKfy29NC4h8zCNjYjDdfwRiR5Y1
U2oMSUpW9OT7HCyGrMatSNps5Pnn0UWPSJ9yGUv9emCLwhhpw7vt4qdK+yGgRWr54Y62DBoXzRPS
YoIS9syWzMFjgQYdu/ao/CLCypJQ+zSU7H7bYTk04ksp1txfxRr81B7GGI+886LLo8Sgw+wnk8Xr
Tx7HcM43Nnn/M9wuA/dnHxG75eGzF36ozOOckXjEB+Ie8uRnQY4KYw8gjALUb28LbUZVIKrZc4J2
7hT6fMPQb8VchXDZRe0hONslQY7ZJKTeG4SCpPunlOLI3FXUHmf4gNfHjPWOTVO9ofFGdUjBfoAt
jHwv6VSlPMXWvpLV9bubWq3LJCyy4VDXMnasB37nsToQ2dMT4IUKmF9iKzwA673ibV8a9kj3Deic
tWPc0FEMS9n5/607i2IhhP1phQvwg8mep0Q6ErvobXsTxgrxWQnHYrEotAB6lx0lEeoAnADOZht3
w2nByPYV9zrJY3OjwTj7UVbDmA+UsWkQNHe9SEnXws7LuTIO3aZNkt2wf54x+9WHteSAOOhjTrGo
+8IMsnxspZIlF45T3wolDnYq1ocIuLgszAh+4stbb2QWHKoX/7u+LmzzjfTv+gBqSDDQk627kuKJ
nxhYiPWBSUgcJenl+KdpDi3mhuvAaEF1647IAsWpAdBCCELE2f1x3b3Cj9aw28jpLEpHtR/9T7kk
xhBI9gKyEknM2J5SPNyxqlwBIKxw/g51O73DGkfhXi4LhfKtDI83/wilxH2CO1o+4gX4cArRmYOv
BAZujYLI/hfXWkkpCIm8X/qCLeg0fvZZ5WcIeVlAlyFHIj+0RqxvtLD+ovGMzM8r++DrLjxzlzu9
GeK4jteqfKf9lpeRsTSpPoo+OuhHvYfaHjw2VosGRi8wfNJz+DmhcyaWPEfq2DCtIDHcZEbgfpDO
5V5+gWRPznZqBBmtMEE6kTUeMttV7ql8rbQDBul3DZqpQRwxl7aDTfddWcesfuqxQe7bmoSY9aYF
63T9vwl+gA3r+87tKhJCCsqO/laksxboDTRAtL9N9jvyaDAOYZEYxpaCB6eFDfZNyHQ+26H5YlBZ
tnDeIzxz7xCHXd0sbih9jfu8GqeM3UwNYquGSNiMbD04yIA2glmbuSnUTejW2r76RMT3QNed6OJF
sSQrMvsG9gGCigjXLhySpP4XlKrW4Z+kQxUc86SnIqNrON6UiVqnMZ9Mut8Ws9j6n5acjDwlSBmv
8Q6rbQh7cFKwnzVWJud+b4OhxdZX3fLIc/DTT1jmTWU2NvTNSlkTvhMoqo4HJnngSHTFDmc7kaGF
NB9ILfrtJ5bpr3vnU9rk7qTN3FWpo52p4OGXVy81Vbu0QHH1Ls6uOa9EnYiFCSOre/KJPDzbj8mJ
aC5EcfO+4/peHvanXHrJSDK2g7nY2P5ik+yhFLwe3JWB3dXj8+HItRdyefKLsIIUJ/RQzkUs0UOW
HTJDyzpSiADG1/V30aM1Oq3RSIju7FGZk9GPOCpH0178jM4W04ZHERYyx3/ImfiuoYC6/eWMhz7I
HMHh/MgzeGCZoF/ooBCN8oYhVYmdEOiYzIQUu1i79hfAL/FxeRQWPrLGxOXgILzmetEkkZ3xVOXi
Q8VMoD+dxH5JLV5ITorcPwhaQZpBRC0DcHyEiCu1RHYLD+DuurJkV9SNJD2jPEB/cN25sMP39YAl
DJH/pn5YMx3nO+Ps48noJObhhg+Gjo65Qi05gzePgczCxbJpV0OfWciZkz2VmnUWueQH9yS6rumZ
WBduV4osrk1sC9vCo3aCA1AeuG8I8kND6+BIqD9/hjd7jacCKoMyxQdurwU5XET/4YO/C//0C0EH
gQnDtym7CcD0v1tWCbmXHOiszPWSqlcTFUjkwMMXqXB700uw4SswbRRYdq0JkF0WnT8swnSWXygS
rHmAD2pBp3u4AwEj97HDu1HM1EJx7nyzIr/QpmXnS+Q+HOIlECK9z/BoMtSfcFsSSKdKlEhH6qNl
TWdGOZjQ7lmj5fXNSIrF3J9jMxU+3pxmlqd/X8sb3zW4gISbXc5VZXbgEJjgxfJg58ADWMzqjoLi
qPYZA28MCy376DgmnQkV8t19qMXopiglBDNvUvr7jkaYBg3AvlJXkepY+SvIYNefCGZnvOTbag/O
jgwxR2sXnxfUHZyBerxVMnRO/6vZ8DdlWbbutL1oDYQytxBx83ctw7mbteIAQOv8Oa5hspqgu/0h
Z9vGZt0Y9ohIQGpBUMyMy4W2t/cufWJOdcTbGhmsP/aG2DBz9xuXNVY0StFBW47LC5sQTIwYhTjn
ZtZ0xyJQbIbKsVlvMhIGsT+dgVo9PoOZjOChzgnhPYCHtOr237i8omliWxWU9Y0x5+Sb37x4cz8m
A9ee0dDPyO2+aCk0w6E+Vm8LRuA4wOBbjhb1wXhzKGs599tKq2KGMTcW9fzZt56QdsxA5Uet0S4N
gvamEVaumB5+BuCGSKndxvmrUrlaekhpfRl9SMGsxHY7kVIyQeaG2DXH8je3kywst/3TOOUAkXb9
J2WY3LTGhy/2V4Od7r/PAK8K0GXNz54AfWN0Pc3UTtus7Y4u+pzWYHFkbDv+WG9v3StsbwKWSpFf
zNqvwjA8ishiohwVunzNKKW5EQa6ZqCFkvLV4aEFYszA6oAMc3tSXRLuM3nB1ckd9vYFMKJ3+UOg
kuZoW2KdQuAWIFb4hpKo9U5sf2CcpXdYiNec1knNxOEkYL0zjTmeWmEfUqBQLw/EeW/7yhwJJ54r
pxIbnh1FQEXahJQYs3VjDrphlnjF9cHydAGoEVImnfTkFLxMLTKShua2hByFwJu8rA0zUMC3lzFy
cbkGqcKeqGU7fOVP0tBHt0tQG8KZ/OeBhZrGSYtG0G2InTlXm/vqPLDLiAI82JxR3J8ed0F9mp2R
1ANVE9tgz4kyJX3WI/TLHnX/jPznuEFIgaWPwef3apxbMFCmfy5AQVORnz++YfycXAo+8i9IUB97
DhxKvtEgB5bFui2qZKxJ7RTIhF1aXaJTRHDGWOCk/ybzsuvt8i6QhGv9QZmUCFttpgzpfmYlofgh
BE3SRaLDCDg0gKs3gcb60z/gXzTPuRs2rphTXkePqvmTMlCPgQkn/5SZsklwMyunWctXfpj7Kpcf
FSIO+wDOer8rO7ub0UOf+ecJengCFn2uF25pG8rXu8E+txCYo5qufBy68lv6AsxDj7C8qUYA4uwN
xss+7PPUMP8hdLEtORg5iRy4gujZuNsnlYzNuJ/e6hP859SUaXQJwjfc+yn3RQp5Ca5rW+Mn2xgX
lA7FsuFhpJ3Is9SdKhp7yuE7nMO3WXhNkP9iHzMLuQ5CjsesrCToz3WsYDddXle1Yp/ZGLwE3fCc
xeg2Wvm0Me6E86eQvfj5G62uPNukyTEnzFO/6chPD5IHj03WsVapfK3Ork8+SwuR++S66SRFSzkl
qzp9MEPyFQJfVdB+J80kkFy5Hs6R1grsVMix66qKKn0Wd5H5+oHHn2eXMGbCUAS2vtk4lEj2myTR
YE4eA8GiXj4fZOop/rrOKSqjEDf1WfArareb1lnjsBa6rP1xKFJ/s1427/RPLaWZP0BWzXwojsw7
PSAih51w5xPbDCeoZ7pKAC6bM8fe6eIDTeCZqxFsexGNssIEHJd5HUBXT9ZtnVX6NV7t93lAvOy7
kr065eFf0Lnzw4U7bDzKx6ZKiyxTnyXehL+DkPpbB9yoweHDIgT42ujkeFhYsiOx5hk6X7H7x8us
x904bifRN3DJdcoj1gdcWzmo//MoOXRaNVhWZy6kMnIYcMsfpj4u5Xse9pFptXJmoL6XMH49zlD5
Aymu+gk0g6auoYVb2zy5qEjR0Zi37fClurZBvKA4D1htr+7RmpSVMVrgtGPcCkyJlukNoqvjvXxb
RPYXTiHTFe6K12RxplY44oql4L+5k8Bi53K2wH8qXXQY2ufyx4/CI/4cYXysMQtpLDv+zc8xjVJ1
oC+2WK7drWbraa57OhQE/9/YdWSie8gxUnD+/pzhsrO+32FFy6vcEf6vsofbSQdYksbNxsJOoWdV
U32HE3RpxFYQ+Gzowjdhg6SIFQO0tYm5ekxXV72OnR046YA9hwHH94rxvLequQNM4n5dEDkB5VkH
z8IZv3RhmRIKDBUsZGi8F3xnE4wvK5Z4aRN5GZjz6teR2UXKn8UAuvNws6P9qL9559BTmu1lGGdc
p+31Fj7HCrvqzGIABHQeRd2qyKQIVo28Fr3/PimMU8AGDVS5t5lQusRW4dNgz9uEOdXGHcplfvIR
YMd7D766AVKxbzkNuOMrCwcsTkPX0AmBz6ERtz8Zppy7caCubTsOLtby0nZsKf/GH9zV8GV+xzKv
+2bx6TgrIV2CLtdNMlC8i2ha5xRp4TocDqBInHF99OBD/WtSFL+7FWJyd56Mf8LdDlnX8F3dFVmE
mZVDu6UHQEgiH7e0r0kRnAv5oQ0Dg3Yo95KVZUsFKL9n3J2B2hDT/P/ppjWyy5uml0S2bifmLveo
6/HCTXdT96LvbBujXrbT0NmfcOLNA1pNJSiS9nGQeK37ltaeOncOa5itawRLm1Ly4ksLJtvbs1q8
N/zM+QECrr7z5ZyQz10+hrCz42U8Ub5NXzOPhIbnvLbX1zIuih1x263i/wgn/zwyaEk4Sjv8cCow
lBt1jz7YuK1eYXJIZSNc6CMkgsTzwq/mIn6q0+muoaybmYdCTb/uVrGUq23ndxF66qV6pHFDFaaD
nx6HIuF82hThsLHapPmv/mXQ+JUQRnQYuVa2XrJL1o3npErJWBVJZP8MwsnMGnrpcvXgfHwoGc2c
6MnBtV69fX8GZTnEflSf9dSMfx0tLGQY7PKra8YwMWrJY1Q34TTm86QxL/anspHFuFZ60Lhgz4jh
52IWOSsJ4qWoto331jOLHdczahT4i70rHrxA/uU+jKg6Dd/UUNTq/vx2MEEMFOM5VmuTYNva6uUS
F3CWT1t7ydhD4Jx31ZkqPgDlfxHUPbvCgUWcBU5e2ZFsUzCQugSLTMCQ0Q5+1O9ysLdgpuozQZOa
nLFrZv1gHaCzVyvTBY7UIR/Kgm3QNogEa5KziZ9rWTheNbeQ+sfJdzMwBU4d62gGrL0URa+fYAjx
+o6Fy8YpznCtE8rLkkZ3vzrBLxWX0kR5FQVYN7C81UCKJQ78Y9l26DeTykACdieXVIykUBkwVjMZ
QcVrgkHFs70b9vCdvaLm70iC+IThWnOC2PQKtBIO7Uw2ITzMYiEiHrNtN+i8eOgVNpEPEopsbrmU
/SlyoRjkCfUMMDN1fWKFU0Z/uPLJ80vRhwWdfGJVUhHkTJKUF+hdtAtLQozZ474E7iWSmDmifTaN
Akoj9qmrXqMB4PvR1snl0Q1/Xn2C22f5cJ3Hfpd9U1iLi6bsNETxBcmr86TY40C3iH85M/pyyJdZ
nM0jPBfFgP8nQwCWXziXKYjBJyjGbl4dkVEELTEt91q46XeEai3h8eCIPs20QhB4zf7Pdt7P7Om0
jSl9OdX8PqD+WWnM8GiWnzvO/VzHnR0aFM2V4G4WlpRBEVuffYS0siToui0LwmaNEEtRqWMpl66b
PW6OW6i4nqKAmkQSATarDVDHuaRNRHTY5N8aw0Xf0FJOHzUD7kzScHmVwGztk3tIZ4RBIjUS5p2J
C+MQ/fg6ukFEbbmbx5znF+Yp6xLtOSH4gftaWmQlMhgyTVgfyLyYSMD/O8w+T9YS06vThMc/YIoY
/b35CbE3oTz03nfNeBUDeu1tk+uF0s3I2cAL2EGn+JBk+RiatlFpGw5W7d7z7vkIYSlsRxnmP0lE
PtrOCObO2PAYw165Lq55/wTvjxSCUn4vQl4yiwpDsq1IK8bW58Y3ARTfCuxsZ0yuAslRV+UwLQlD
AswkrSQLDcisu9iphKj3JUEZtrscNhZlPPSxRKrD4EXGXYzxtmk5imKnFk+KCGf359jftDV52Ra0
/ANNTqwvxHHUSn0RCxoBa7EmfMcwdiznsLwWPHhJcDAd+F+QETcAf22MyXjdd+Dbcsktd3yUXsGF
vPrsteTxPSHyWPghcAP1RYcON9sHC0FOQjSQj6H9FuwdWnHID0qtUrueEugp4DPx9ZRUkaOxI+P6
6EXZ8do4V/lH21Beb8GIRsFi7MRZr6CxdmUb6dKZzoMFiRMao7CF5RpBreYuudPWaS2XKlMLMqVg
+Ucgrm/PyLELdZTXHl5AjRbGEddp1R2NfU2JRLd8KQvTgjIrsz7VoBAEnTFiuZcrYeL6RgEXY1Xs
EyES/yCOZ2CigOwPkV+XdHaNBYbmTEzVbWm8Q6Bm85TCHCS48pY9QilQtMwxD5H5gVzp/M/6lz0g
z7+AdOe45E2QgzKCed85SYmWfbs8HhC3uYJMFvncVs5hU6Y/1FN4LjCCPmjGEVuzB7KlnQwMDyvX
fX8YMFbYy3MG3sAKP680JUWz2lUt0UaFmZtWmcPBLnRUg6h4k/O2SXKheT4KUXp0HZvKGB0pJ/BN
rJhO6ukXgzjgi3OzgUQltiKXQgXUdnKUDbbT4tY/lrMaUjarhXww8cP6636Dyv92SueIZx2/1350
WQMqZ1+ltXfZqfch92k50W/pHE+4KyXxSsRrBRvZoDFJwz18441XeSiqJAECiS1KNdATHKuxvqph
2RW1dbEgwfGrSnTDaGx6hlgGeg71Fsk+FTmDH+3YEu6Kd/Jv6ZxPivzCpMZECMF4w3jXJQh7PZvT
N0/neI+fNwU/Px+uFhtpLL7dieIwXPniNufyp8IQlG1DqOOG//udd8QZxTFCekP0BoqVfRCNog9X
2KD9C5TNr4/ztmKZN7PMOHEMtbOMdd7u2m8okUPijn/heCuyL6Wj7s2yhzyBDk6W1RtDTeaj0CIL
6MZGozCysiL36qp3l0jOjjhf3DSetgWdO0gbrMhddJB3wxwXK0udOGIEhPsugDUDBDA9FD+pmpDa
tpSZjTKelNxtIlIC8URpEo8X0e3GVZFKoSDNlCG3XKsxJ34emeUxFjd7ontCv9khRMTa5cx/9khM
gjuKuHDLuuwN6awtzWSaJmZLW8XBw8C0DAzNdwB3/HnWCRW4P+YbDBce8fSfWihDQNIII+VgCUtj
+ds2tnExLyr31i7xysmIh7RHBYQqWysH/fMw6P3iA7Gahpa5pZ1GwpVAM3X9cjf1TVF0D2/hG3vn
b4ODGNyiNbpt+kv4liCcJBCxPVJsrNBKCf6NHOxeqNp8SOX/EcE006aqRb2a5yDTBmzwlVllrIhh
EekMKhIwtmkAIQrc+/WdcEOQAUFdMF5FZB7FCV/F4hI4sRBUrG1bz4tgounmBuipEYg8avnpAWUz
5e3FGn5toOyWqoxmrDc683it5FRnFfWWd8m7vUaStHN5JepqiNeIZ8eZJdYNYrLe8hbG3kfa7BYg
G/jZICJP3emZfNy+AOriu9/fs/nNfxnb/azzgmq0Ja4JWL9uWLgq/oaOgMuYOaNckOrByh3KizOC
U1PCctX/t9MliVU+IQxQK0XDJkD6YUyCbczVuwgBcP1wodcotih9Ab5hyFyDtcIzokL8IjnNVpcx
+6dXVzLw8ejdhpXspDvawhrJBHWIsKcxW+a1Emuz+VMbq8yuei5+xHjT35yOe9JDzy+AeLNRZHjX
L0BmgG7ZQKu/6msRmSdoRY+Wy6fKRrdF7dy538fSWkFRAKgmpJRpEPghyzFbUMTeTR9CJEDqqzxI
MNYRpijuFFAJgUVkZHh0Y0M0sfBGX7FTGYJAHcUhEnYERcJZmnBAxBz97dMAMqt4QVdd5Vw+FFqo
ph6lQuHvpXPD9LS7kpwfVX8q5Ki2InX74qJqIOKZrSv/dUzqeM81KahW67P1SHCr4gbSGqws7PJ+
Af30QK3tmgryHrCvSn6nTs0z0Sy7PDRlluLm6DkeB2e10ypmFimdDCVsIHvVxWsDFg9dG5P4YFro
T/pzGlh2l5aezCzqWFsaQbbwNw7Kd9hxVWyjtVBAIdZFH5rzN/tu+JmnSvepcJSmFiBIiY1pIbte
r3ddwdo6P02uRsOpOn0xfNakPWz6IasyYScGyCq5Ad3DJEGcyRnhdguJuNHYveOxHIKKglRoqrPA
OvjylFNWQsHucP4N1/GjmplWyjEiVak8pIz7PBmymZrQhV2jjmnab0p8ucrZsIn3ObX51ibafm67
FygDnafQOyQwo8MPR5eEYVyoX7T08Qe3LY74lCVI3/IY5jPMdHujGkyrLCVml7KGjYlLtEoFflbc
eX5ol7p3Xl1cvX3hMaUz2KDH3qrM3xm/Ey3hD1fKG8JysFTJacPatHx7+R/ESQGct0kn9LCRpqKR
MTr/rrsYoY5OZHN+2b7qGFcXExjNwwyXS7iCcRCUUe+2LG5v/RLAWTDbk+Zfw9ysXbeRCqDnCx/R
S8FrQqbFy+BGrnR/09y3YHz6ECEBY1kHvWFphJyWOBu4ocysSshIInvsB8LFcK7Yx1sTihfAnn5a
eyNxYfyXBzHK5RJZi5eTgIu2V0eaRvA0vgavWT7ONZHNvXg0L2SV4AqDCYV60SD3d3vv/pFVnm1x
aQ4dopiGsCE1r3Vm9khZsBmcuZ76th6ws2yFBLAxRgUPGoD7lPRzoKP9ygRDoXBmJLHeXxvkQZ77
de8iCcHE0QxjqlqYGwW44kdfaRAIUmhH5R9y4EDXvzQy+gmsBHhPFnzlS2uy19uP3KqeEwnwIRP8
7uJ9fy0F5MP0qQ3UxxEV5h/rK7xfeASYWVtAW3DphcUcool7gxrgyWC3S41DubOXStkJdbLAMibe
brDJ8bYTgPJvVqkd7317YdKiX768RncW+MFT9n+yMf3d5EeTfgmkjqUYXOeh5/iIeUoWIPoh5Kl1
sfpfQwHuryirmRjzsKwNw4CAsShSQ+e1TXYrLeJUzLqe1yjA3gbqsLNPjdtVLAitS9vdd0/NHhAm
NTYM3pp+auRi6SFehe1eOISWZ/9ioTd0Hl10WBRR0iar3sOesJqMi77nE/EOC9XAckvZSxdsGRzy
VxixZJKRaYmwrtHcaLiY5/EAav2hz0hIK6ihbyu5Eom6s1XJ3YBJz8iKTkn+3sY6i9/F1kT5rmLT
iyLeWg5GrjT0OyZPXCx5wXKvIkZh++ETSCj6x1vlWEOWZafjM/bd6VjR5G0A0bOPtVUBMHVOWSWg
tsGQyOJHlxGv4oLyVATFuLPHz3eDan6aUHjy9GkJfGTJzaJhEuCF8xHl0wl+Qvf0zL5XzmG9pn6A
mAfNJOkHOD6leTLXADxZgLQ8FZ3OluF8v4Pqd37VrhOOimDZX7MWmLVJjjzYGiU1qYAo27z0hBje
QYFr7DXNQp+15xzzP9NsqVzkmS2kHcx26Biby8EDTannRrtZ7tHWwYKr8wIyihFB17LPbQ3m4lKo
B6argKfRA+94Ff/2bVpPGRrEcxw3w+kQy/uPqqQ9KMfbHNoixEgdRekt6/IGFuBcplbm4r4aDGJv
NT+LAE4U10f66nOU/36Hr8hH7TTLgIW5lKfbG6mcp9vZ8rFz1sv0Gf9XebGWXcEaDY8SfeZMS5hS
w7pfxi7w5ijLosfLha1PCX7JWBDqFQKWIfzSbgPtf1nptXSLueaDb3//QvXIhJRhGZGXRtkkxWZi
+ktIYEH8iOE8u8Hc7WrFsjeLpZXnn9UwVMLMV2cb6tYNCpYMOHCjoPrTfxZwPZJFueCKe72jqcHF
anU8a9djd23zHjaAfVJxgwF59Mbty3Oh0jBsBw6uBeuNVEDMLwVco1kpZ9khaJ1Gx79HWfMoiShP
vZbw+0ZztBfByXny+bdI2aM/sRUqbcfCMFBlwfGOtl0h0pujKOU1ZNmdysjAqgf/gdF7SSAfZskP
9xXNbQQnGdxJjqeH/5k7eWmcOnb1uO7aIaBvsm+Eha/3JBy6RHepkTIlPhs68i0nM5EuCI8ce4Og
w1Da8G3GULQk4WGVWzhXxyCX4TANlVa2oSRI93JUL71R6v2Rm/bx69BJ3fPfFNdyP8H+46f23Vdf
dwmNT3FYj/+toolvYchmJQjaL2+bAiU7r9SkgleRrinBZkOzJ8xqjBVXSm8u5xrknCt9EurOyRgI
mavxVfED3SMYCBuc5Hf1Y0cEB23ZYnhY9U88dDoQBSz1IsXBj+FnIcKFlsDV+tWofVP5g/SxsQGS
aXyrjockg5xFHoFGN99Os766+H/tJLnSblp3PF1XM3XpCZGtM4JSdJpuyMwIPV3Jlu5s+DtYku/l
gL0Vda0Y8uoLTzxEfM7+Zj5c/A19gs7ahGN1rEwH3DI4M353xDzT60WlpWlBwbJHSqySWXC0OvhV
suZuXFCt8lVNmjPwEcCndfITzH3KCs8thG/SNJs4LY48v+qYDp1RauPLMHnW6U6Ikgmapgq5i/kG
r1kxpqTa6Ga+xw/kQ5rak6/vtH+eTdrHM9f2uCEE7/Y2E0Jvk8wxuJAqP3OZV1iBg1krNj07mim3
8CfqdgsiOP9+ZMDRZBarVG8HoO5PDAMlPqhfNbtPxPjozLkassbTaderknmWp3eLZXw6N5pVSu2O
geOXm9UjzREkFruo48IQf1RD3+GULYlFykYxtGhLPlKXZCWmpCuMX6xot6hVtu+ovB8MBNVfgqog
DZUEiWAidA7hr6qUCHtQZN0it7zhoeAI/zX/DJs9iIC5SmEuO/B8T+TLjL93OQQUzdt8E0qKoFQH
wXoVvtv4S3DbAbRITnu1c7eKERwZgh8iBNc6IXQA4Gd769iSVAfP/m2TvT6By4nVzf8b0nY8LZ1k
B8lxgwNn7Lj9NcleLe+hMMKDXUaBfdApslt9Gzkr5IQlEZIMoBPPA3ii3UEJwv1uTwQbc8lOonMR
TM3J4VbPhIiNRBg8GUB7BXh6fLfbrVaquoJJKP6DvHctjIXxq3c8VolZEg0STTfocdS0I/OQA42Z
sHBXn3KEVHXVYpkFEzcg3cLZUnjE8l/SrhG9Phmat+7VTB1P2s5Tm7yEEZT+z0riwm9Q8x6lram2
v/2jIsC/hNWwkozQJ8V3xx+jg/IJ/7rr09XtnWJ1ythrgNRxmukTtDN78Eam78Qz77NBcUKzFugG
qyUccFcahUx/ZFLKG580RNW/iLLp2T9qDdK+MMnJarMUE6j96lPPT31F5ArnSxbUe70JzB6iapEM
n2Byc5jCGo407Ji/ya10y8G6FgGQ7ZbEXP4LDTlrfpJLFS9NsBf/v7RyJ+06tPaQx3BpTJ+++mQ4
rAyrEVbmujrKKrZ+9PjGoIWNgfZKSuIb9uEYanub4P2qW1HVv9tcOYP+cpHMAjUm9pb23q4yJQ8k
J6q/+rAkpWkg2kdnaqVKe8aQWf+bkYGX0liHlPuD19Rd/2Wst6ld91GC4B8ir+YoWGFafsHcyibU
RjwElegXeeXBu5sC7hJ87W6W57jSI2dqnAZCd5G0eOyHq8BR4EfEXJGCkDMMeXOBvN132eSr6FBk
nd1qVGCyTRd+qCP8pn6H+f1PsL7ypszGirYXJTWh7Lmjme+8RXJNZhNUqLcZy2dix66w1cdzrP9e
6e9M+C+dqWUYyHQoP8oDMfapCxm2ecQTkG71YncjMVesh6KcMMrmXo+d3FrYJ/fDlsqohExjcPol
3uaBudlP4ducHjKQw921wgrI7sGDXwtaZD1xhF5hCPdHkDQM/eZYTsYl7gyQ44lyzx1T5I67m3n4
mooCqrBS9sCIJsVF2RDyWgJNRZi3gLNi1R/YEBZN+dEB82/t+GjAEQkE3KQcwDau0lvVsNkkY3JC
xU69Cis2gbnQ5b/h7ds44i/4o7D7D2HgxS6wF7x1Ts1PrK8jes9keERh1O8UxRL51kjYii2Hwgiq
dMuJaX0PzCsJ9iLn3yfos/Xzc8NUuL1qDWuPz1INe1IciwXquCIP8uLob4qsw93iTCyaHUgnvurx
QO1FcPD2XB4WeYqnrYTkucnp7bm4qo8ORAFOUUZw8T9fAbkM/+LkSBm6utvpsp1G7PBZOPuurMzH
FyF0PJUgXuQPxIiRzvk7q5HV6EBRQ1mPnQWHQiQZfOYahAlZOPQGdwW5f3m4qygOGbNsSKXAikWj
kC+tVGT6zsoxSDsThkk++QOQX9U3X2/wkzbUKDGFvcLhBCBzyDqH+1mDyVGCmFG3fKe6p7jLG62C
ATVqTodPC2szNUTGom9KYNonNb/dSxy7NeVgmbP7kntkOGoab3Ga3e8EeJ115hA0QigIx3LzIQvQ
snAG6E8rBPH3MedHfXnUNJ8xDJsmARf+zRW8FcrtjLAkG13OC/jhSthMNF7gAgZQ4GzB/1Ok/2yW
m9ZDNCFRULsU3iFESE010QBvkyjX1o08/D5janBZQZI1jxxyqn/tOxeLdP9jvohlIttN3w7qv/4u
yUbUqAIRs0+79T6zyKkdgrDjghmqEzS5mkGCLYY3R2PSLHnCByMtGfuRgkAxywQcx0yofVgaxijQ
2yxcE8SOK3bfP3pMm5On0WZenxaXVbKXzJGvaycQD7KFG0udWuV2w62xkgR8TiqatFr69HxcT0M9
rj+0CbLz2o1x/WlP7Ybl4hLZsLBrgq2CVgAezUG23KxUp2t3Yd/rmoVeBdK5eT+EHQcVLM5C+9c6
QWW8pas66VPWcPeq9VsSQJesZLzFzt4NMSzKnbB7Ca+NcfJeZOGOVs6USmmmh29WohxBruopP0bl
MLHduthWC9Vmz4gejUn7pohqqLpf+pW4/dHrwB8uYVv0EHVmmxyrkoVKDG5zHQIAT7X9Mf9C38A/
Q8XtXwWxAEgqmENGHonNwoe/MzqSmOZmkArQIHJXJxhxV9wWzrAHe/g3cDVGSxyJ86y7Tc8ySTte
SUtGKKFVFgoozsC/ldzZu3HMwFLfjE/te1s2bPxOEa8xVmvc5TgkLgs976df0r7DdCzkaV9WznLP
Dr5aFlTUADpE+18ZiGTZHWKB+XCK2DjJPYjNTLQGwyIT1oqu1bkzqjDwZ/vaqjo+auuGlnsjtG64
geXyW/FXJpE76371rWnIAvi23zSyqmkSpfabZNeycvPHMMP+cFpGc4MVqIKWOx/95TVgymHRR7GN
L1bAOoi55dIRiwIn6aLmE1PlZNdx0KCTk3mqcgxEOLYJbhTYVS3ap3vsAUiXKO9u1GNihfNaV5DY
tasfvOV4rmzscZUNSplqelQqu/T+CnLBNmms5pq870WWBdm810mBs42S6pkg4GnHEreKw4KWNDFv
5gZkZCmBpYNXzGh80CjqCOV6wTpBdX5SkVKUOCG0rWdyuQPXAhzjaBJxhGigznrwRdr7uNgBH6fk
MHWkcHvwwAOkrxXrPU8aKGvT/pTMkB3IOgthoh0bok9m9MlBCxjfMm0iWuL9Iejwr24JK7XG0/wq
YLAGcusJlxH80oezTvIPkmrbEkgPEUNgUBv0CIrKuuMB109v32XCfFgKwJZKNKBzzVea712E2zFB
ObVZHPoUOlxxwGJ3KSOTMXRM0p6NZrTBNVDR7U/Xdc3HLiJTWoSNgHHl8fhLsm46a0nQgIZ40TjI
MG8JFS+gDaJFEMyWFabt4Ryry9m/yK/9kONNQQAaeO6F+96i+rcG8uVPOIcoTqbalCiXs8wBpwTY
dZo7uRjcYOM84bMMdJ1ZSQ8hc82jcwho1++Er8cnyZtwffJyDo5/DPyfHhJ8cl62KX31k9AMFjZx
mmsfWc88XPYPEuRgA51Z45bqOj+Hniyu3K3hF6RTrYBPZxvazeMEV+qBmHnFuzmXxAnYpBpJ8SWA
9+vt26NqnvLIMRQq8aEy44Jy1/ceuTd1bKfs+2V0GtIHrQ7U/zasTEts+KF70RnWaZAlxgBd6ASH
aevnMLIQl0SlK8kdpOAzxq9OZOdpQztj/N5kVSx45xPFoJ+WG9VGSyDza626wyi2w6K8lAG3xXNw
EP3c12EEy2RejTRCl4dK9N+uAiUGXOBm7yNnco5zNJ4zuQG0SDv4lbSKzKsOf5UutDAIbeeM7bHW
iSZwyPMaLrMyNOZhWGNdWxtywwkvai2sInNUzl+LxO+QUsDeV+t+JTNCcA3GUlvENVCFS3+l4bGR
RGi+UVTvhR2os1pFvAktGdrWlYs9W/v5Z2k3dT0AKM2VTrgC2zo4XkKRwh3eKWHXaJuDyDY6M5yo
TaUadjea6if5cRcVeUrimmiNMB5rKkSv8tZrezl3WUSkX5DXapdvENEvClOiwVSID8/PyNfMFVis
X0gAmUNcHv4grOFIiJIZc7e6xqVgvX1THS5dcbXjhiEBNhITKfef5qkVAoy+trYrMVJGEE2LLOBd
jQz6pcz1N1Qk83KVe9Dr+LbUXNYihSGWPi9JZ1yVg/mRFShXZIHrVN/Oby2Pveh3yjGZjU0fZh6x
xQCbp97GzY0Ujxd5YlAxyr+rw/uemv/m8GsgD1dZlqziAzb3UC8e6s9nrIgqZ0DBCAYpS1qIjMdM
EeOIzwvTnhiSOt2RYMcIw/Y/fvy6ae6i8tcJP+ZQjNMNq/g38qrbtPThL7aT7RspSacwyxX4mbEA
Slg9ha6MoTSkGOgW30fsVZovbK/FEM2Vz7D2ff+58yoF4ZGMtRUvKqGGWaYIJy7lwbDZqXGru3ZA
wdVq69X3XSnMMYosxLLnfXbmq0tDOB2pq3b2xlwN3Q89O7Xv3F84iOuLYAHDW90xd0M/BTVuO4hP
+ZMuJtM3nUGHeokO+/56sjPrNkkTxN0QU3dqNOc+fKsPYXy7HOvMqBbVWrqYoBygjwwYaiFbZ0Ex
BiskrK6SwdEXKyGWubiPGXQOMDZCBb8JA36I0lyHx6gHs5SJtrcwaClYABTWU+grfdj4YRNFfABU
WLnvojHHA8OBvD+ZzZdn8RB0u4SZ3972aATLuV66AkeDWjv4/woiOZOYhhHBGpkMlOMQo+e3HxJQ
SBPyaqGcAOUEgHTmm3BKTZbzJyw2aITNOzofqloX9xpF97BmkOOtsmPdoRgvZ/yXWEKBjdLgxeBr
ndDODeCDgwsFaASb2EPgXQrnLj1gpilEPtnsuJAH8nF06g3mgeJXU3FYfvm0PNlxm5ujSKwYvoZH
+2h/lZQjD6rfhyDSqgSzXDiaM2k6Wvwmh0tIKRAw4O2D4LXHg1rLBME6Sgj02iMZYv9T6QWTTDdw
Mt73PQdQXewBU/frWPYBd1OMZZgYgSqnK5SBtmOuPTj4LOaQfuAsky6v7FGl+Y2rNaTJDN5triFt
p1rFdnY2IQZ4MzK+EAshsBjQ0wv2J6M7KGUYwhJdqAdmlzNXbGX3Y5kHE+oMBm/0yY1xJ7E9G6We
i6A+6BYJ81koqyC0vle4bHFFFG8tnYQma+AIIHLEFgu5MHbnpjAx3DuvkQmmHMhGhIyNxr2eU0Af
8NFMZbDrG1WFb1EDD9G8r1jc6GimciPhNM1zyLM9c6BYb3KiUcqmW26b1J+SFBULfGAsIddMqjto
txBeSB/U6L1IezcKApd/BJJiRHm3iY41gzt0PRLRroKE+ofZpTulMNQTo+q2Vf3PRDHdmaBMhAWY
hl8cYMK+YAoYC1eEV3/cKfjv5nsWgXLYOqjtyZL6vqdCgaVeDq9xs2KLPgjBOd30V+eACOiBQSst
bNY3quuPf9Tk2qNwTCtdDmaoLKLQghNCpttFA/mpi3/pzvk3hM7AydCYuzINiusHAtTcBrvp1EG/
2C++YEfgZq09rbKWmetXUeytGCTdAC/qtpDMBm9/F9y+aar4I+AgAE7XRxAz3NtfJZLiIpvnpPpL
/ULKWkdwyu3oaOe4u5HJuAUlyd2l44bWtkJYqCYXGfE1hsB2ghjTNLE5sD4Uiag+wkV028pefH2A
db/+afXmrdJtsu9vWfBTieD1JPuPT1bHUtEKWlrD5bkN1JA3IanID+eqnsuhhVKn70eXfdNtQyIB
sD0K1zyBXzgrBMRd4nrN73t6q5HShhx5V7Nk2JMGkzOZ/qg2sdzP/lCF9blfGtFd3iaCJbwylwN1
3Bsp4LTXa/KuND8YVu1mEhx0PsVNBuXp2nniNzDZlgJHA0A6/phHtukEBjQGIeEWBTs8mcJBcSyf
4GToqXDnal+EZyGcNl4dix/lkD7xfXiGXlrCr1qcPyOWvuCrl8EgYGhtIMn6KW8SDv9beJMqMRgF
lEHnoaBZB695rUOlzWqWaF8OdgU45qpPEmIAydEl0OyriBZSg5YOStm6mrAaqV9zXbA8+glN2OO/
Hwe17mNiDLx3FrFd5u6AfqFK5bFs+C7mliKPe04JwcNFYRc8WEAtC/aIV9r6CKFy7utMTvrPnQCv
PC7djoGyW7JlQE1annXzISwOxSlFeDfNouxvcMszscRmdpvq756dp1tePBQ+RoIem9MGrUCUKKHb
A/DRxUDRTebTbrciOZOkM1g8OiO2jxkO73yoeCFETsl4zJ9NqueVJjRoSnI0Ynvxt+LVdK4RB0V2
jov7//PSMfaDa0v0nOOjZEdVNRA0ONvd4EoQ/yv0V/oJAbJQIo6caKjJ+cEk7BuMf3sZWW6g0+ZY
Ddze1hx2SBT+Eh1rgB+DV1zgtbrCKfPm6C76dGUWpGqeZjGb6eYAJm6YZv1woW3emexj2RcG2N9t
E9m01IPAcata/YICMGXLR1xwhnZBHHmVW5pDOiInMND6oAQlGMCOL3boY2g0316qKlpDt6GKqeB8
811TIBEzkklmP00Mo6HNbiGxqqBRDnZGZk9qyAbnkOTb4StVlsVj4vzH0tVoXcXqD4IO2ra389H8
43bswhelFT6JQpNL2WfPdm8jGWZA9SX2BaxLT+dquyJcFNzo4yfnRi8GV0AiwYJe/Q33p/cuBdS0
XGZsJi4Ty8jPF3kE0rHunvrxNHLTUKq4YFGYMAXcBxeZG4NlQyIC7bAkAiHuhL57PCXmt9nXK80P
J5S6X0RKe7uexQ4goVpDTsK7xSz1hwCcY8Gp7v3vKU/OS0bnR9aU+LSPMJupFPUBcBdpq20qdA6C
NGCTr/uxkM24CqAWz/ldkY/XXNQdtefxV6FS9Lv4pWFaBt8zBTqWp6ZHir+Bghd+DF5Zof6z/RCZ
Qq2vhlIR/QlIdPozhQZcu3QNKgKIAJl2Ueh14xbFDNZg1QaInLYy300gebqSmu3ruUwIMkPH9RuS
j/SWzXfA/pUOAAmeGL6klkc2Wla6CKUa7F8NjCf2HyEJWIaoDeWBDElIKGTjylbS9vYtVO5WJcs+
O+lRJ2T5k5IyqCFeWb12+UdEgL5zG0ChO1USe3C9SZzZPBDCn6LatNiG7LIhtgKP3uU6N1IbPf8p
xwrR1mwcwGNqczDXxxTUnO0MTjmioAnGZjWUpSqUe8VB61QFZ4qWs9odIuFov1A1ewPMhkMsZumR
svq19RzYyM8rJ44RLLLOSgk3gNk5cAcgh4Zvm32fT6Yliqd5hoA/zOImZ7TmQ3Ui3Uza8vq4L+/0
eoapE55ckkJoQOJtw/9C3KenCkWyE2538rP3vL6MRZGEeJmIx0ZPemFDlVd1kNKvJJbpEB3p8J9w
oHnI5pKaAx9YiqvUlyTatm42HI3e/Ebw3XyaYh4TKB1nDg/SqrTUBZ/FHIomfnmI2SXDGY7enSO3
M0NlM9AnzMcwP8Kc9zS5DzbiobSV0F5dokssrrFghzwun3nTjtxtL+KqKgqsCEkAcbi3OCei7bGS
Jqb7EJ1i1EaH8VAADDh92LCvAioAxf70BQxxco06Vu/XHXEKbcm6Mo3/znphoH3O2c1N5BS7A27s
/CdBs/F2wnnXQswdWqRZcxUytxWkQ3C9tBP5y5Sd62KGzWduovdWkKaoK4DykCVxkd2pqGeK9FeP
3bhoU8ZatXuR9kEjtmPB7zkXDtTmIw4L33ImYlMYVCpLcckbtyekO6PclTw23UnT+v8NefUQWvzH
Nn8XDuBL+AfQmJG/Caa8ZVOM2JVF5zZo4qTdCUgYDS9PIhG6cMCgSL5wrTYwXiMmdn3KS8cfKwcO
raGPwfJU1xAah+hHDoOqGRELIvA+CXFH8DpFJEyDJtaxVO+5UxX98ZGuz8AL5vLYsTEtIRlm7BVW
3Wb5EyjOIjiFcW33WpXyz6fzNEEqL+I0+IpoaTtei+Tnj9rJjGqDTUyTAmjuB8QkCnO2/Jy6E1zb
nPUNMf2jLOif6a99mdDQZajIzbqVO0b6msIv5I4XA7UcR9OGM1t+ESXJo5Ka44hNEy2bpOKLQ9wM
Mg2dEJ8gc0n+p4uLyjN0ZT1FfMpckH2vujbGZCfSvrduvpRtNCgBXwhGqrw3KxYFOYyDwWe7K2NL
ra1VTEvwAMOYr+YLGzcK780gK6U/nthJKOJyTIknPKas2Q/Tx7Cc/H2xHVv6C2Nn/W7z3CWTySUN
BGVnf1pc9C92S4anWphi0XUajImLjCb4g+GcX1+BPj4r/HkqPkm9+NaRo9hjBFPHXDGkCNKJ/AXj
B2OH33IKMTzuLUN5NWkQBE2JFWp+9PastcMZf14GfycWX3xomhuqt0XA3+MhqZ8z+gpDtqipoqGb
nzhvSdxQ/XMH6GKyjPnAT7SvRiW3MELwE2HYvFgOpWvzsgA4oRM6fYIkkJ1q8jmzqnZE4/8g9CBF
0+gAfUYzrkafpiHLHwL1Hwi4yrOAdNDVn3MG1R+dm2jeSlOvsWJe7prPUiZvUn6PD37AkKUl4/vO
2krvO2uND3AiFsAk1rNo02OEoH68/1Gd5+hTugP2X4g+KgpiGIBbYEl5pRoTkDmlh1LMoXgX6y1t
urmb0JwhqwVsg7+PWSrxgboCTwRR4/xKKhhKQ9X4yp8rN84RZPRomcmmrDNfzgPdvGJxmYla7USO
rMhK1PAk5EywLvRwNpu3LNMf0NtqfAiu6QfBYPFZu1djq91ef8MeZ4pvJ2GKfT12KwYNEn+kq7jZ
7FjDY1AjOaOZEvX3LudSWJEkkRpBKob5U1Qo9jTxB7rC87LVDvemO6B9em7Vh0OqpETpNNWhc2qB
Y1gQbaPuFKytHXRKTSL8s0pWYimbdnRY8hsP/hYF8Vw4pjQhfUEYRJtb9omuwDJXH/lVJy3RbLlL
8u8nlOfYtfAlGVRxaUTmwLYt9DTPqUrG5p3EzV2d8/KmXM0cfr5uGxNz8UqWwpT1gDPaTwj4mo7q
zHlfxlENUPZIXHuK8GR1KwOIA6z3Wmy0C8s+E9t6dYDah5CdSyl7LGuyYyA8/IjetIXpeqOb+tTY
HffMuMjKx7I7PP/9MYAOO48ZPL82CMYosQMD9a7q6yePB20mFwEQjxPi6/sHzcO8ZeaSk75Jxn4U
/kkrcjslACByrhxvAlQfqUu05cKvqwhRFR7NM4xXg8UwAkBiVfPfgVLbDVbUhStTS294yCuMr/YB
3lvvKu7g5z6Niu4tpFbGiKb1xh5c/4YJtpiCB4QafA8JNlgHu28DW7irZQXvHjktQPuZtI/OvG1f
X+X2BAwLNF/znIV+AF6lbadBWqJh1rzy21VgMm5V+NIfABx9AI9tglfMyXznmmlOhVmI3TvmceLV
K7HzoxGesMECvRojGzbniVRMvHfCl6h9L/xKKcfzt3BHv5wloKKTYncAe1AHTLeyObo2oVF1heo/
UatXcbX17sTgRGNYxMZjW+lQPLfT1MFrxYvg6AiglScZDh19miUIELPLaktPEOcV3VazM2OfSDE/
jGZtDuKuh9YW2GvOSPY+f9dsyVxT9ucBP4m8H6QIMLJIJKo7iWjdcmt1MCYB3YM3AIr/L+jzouvA
w/sYc8fwA/RtQf7kFQF0KYeMPxamtaHfvi35KHKdR1NmVpAib51owRqMemP6Z+5hVPleE0VUTAE7
w8JpOUl+qbUxwq2THcUH6eQlrmHyb3AfcZu13d5yHDyb6c4pXYpg0Ccs6WA7c0fDQnTsfbVW1rvQ
HKl4O21NeLJO4jS/2s4vJuLPY/R7O2mvLapr9Q4TEEXpxhd4p7TMKYaiDhfkAXBmajbVPoB+b4+x
uJF5VzIDtnmOA4Q0KmtQw4r6RGqn4WEtLvFsiLXYHLUpVfhsRNnmnGOxCD7iIy6lEGUMIx3Zhpo+
eL11iNS0opWE2zHZacEZ3APJSolnMAbbKp5usdR7/9ahT4WKPRN+Q4VypNXFosehEH65LfrUmViv
zlxg3mh6pTt737jd0vw8K1O66m3d4MU7XW5to4eEiNOjCxea9lqaKNcmgBZF1NM4GBUWz7WEZrAV
MnupDPHCB0AzZN9MhVjVTH8LtVLz8kWu3ppwiRZkae4X3CwApuIG1dlMqaq0xu5ncZuTyomtDb2e
ZOCJWkS6cGjlgJ4HlJvJT7YW9BkTfympH4pF/keOot0xbD7o1691odAtECOk/eEZIdJa68gSz0HL
VtGCg4Lxo7027OXmHt4iJoRk3lDPuX/TQek+bBOQg8ayNoPFTZR0CbU2rYZDahiCE3jixj++HtY5
5IC0WY4xDTl3seaTXVFZYViy28GfY9w3S4GUoVpsIdHJbu052Oo9yuNaCFdGxzBjZGfuw4auiqIY
1Op/zMbGXdtXWVr7mYE5ZEXlan2HMXcy4O6Rv0rA2OuvkFi5sIZWhhywM1TA+l+PqtSFawqLXWK4
nUmJSgPCeDHkKR92s95IoYQ6rhfe6HKr+39HiCDtuRRT8pCjQwRMfCzu9Agbc4PiNkz9Hxy8rTAD
WdkTN4m/9GkFYfipixPf54OCveqbg6AIIbhjBVWFu6WP74J5Wrg5wM+tf3AcciWQa4R7ORralsqw
5jYykVp/ufgtFd/g+EqWVKDR+iIGM0ERg1eEZlSRL9NFj95W99xOz6kfyOYDN2k2wZYsb3d5a2sF
6mW9ZnzhrclP+Vb4SWg23jawDJmYYp39umzl95wHyDIaCJhJ46FHZoHPU7LRrPi5JcyQWfSto1I1
qv/LgCqyAkqPe5F5/PG0uMDKVp5N2sO4Rvd43mQIZDZk/vmlcuB1eE3B4wzrK7tAWoJfzRCS+D/I
MzpJDph/0ZXg6j8ZhbbHiknSnCJC0/X0aesXq7G7KiAOhLxhsHM6JVj9BRNGwIINuMptf9hGFPgz
bEHI527EoKuiXdjP1EaoTnuGFIyofI94I3t+o2mFur1n24wq84pcoK0I9mkPS0qK7bo5OhlENdWG
5YGB3x9edm8tpN63EvA0nBsRifllAHceOF8dOnODXebxcgAK5XkpX3HtYebVb5kk4ClBKC1OTXOL
ApC7B1wbbmgmzPd7gh/JO9es4YJp3hh1YvLrqMbkWfoYDEdkauGWLATR4Szvy4BlDi9ziBKdY4Wx
quhDPyU2BTDb3RJ9N5XMEjxRuelkNV0iRoxkHK2aRZakyjvAH7Ie7T9N/bd/Xv0up/XUyBrrQLZB
DZ/Y56npHyV5+GgJ0hWK4+tKvKzAPC1VpE7bQupT4mhZqh7fpRFEF+rBhvrsZe2pbz4WySbGoZxr
+MN3iy2bMH+ScV2DwAzAeTUU07DQc2LsxOsleBclP6m6gYNWDejEoKJ5JIjLkXHgh7fSS7deJ6m1
F1fHP2XgMGezRdUsFK3Fe2NZdNQO+LoFtIVxbUZlOaBpWHjJu/TsAyBMLGfdtmxuPSP2P3+BcVBd
ZN6dzN8o8JAI5xHgCstIZMwma+zKQ7mibPlpxZhluuHCQ1LY8WYPubjNAGZdvEIG3Xwtj6hXyBwx
kJoVsOfZvUNr/iF5dGPv1YZLuP2bpb4glE8OEVPCt5zGYtox/JdyM+dtSj0BBgDEejMG2oV3nb1X
qRMnoCyD3e/tzBtfKOUwq4v+rjK/8lPinV4pNagFKXRYRJUcYQdzJLBTlIETIEso2UDMGfOXAXE5
6ne4sSHJoUF71fz9kCoLUUtE8ZiKVvwxCFbsgD7SnobkqkapGsfH+7YdCW0JGz/7jFLGfSXJfvmn
LUCQ6DwDcB9jsiX3sDR159oKQqBWav1RcQLCNhBOhNEmSbuEQkGVfYO2BP2LSbT7aLjr/IlFnIgs
sG5cwzrDmmf/4/6nPzEqCd5j0Ayn6+PhqVoyPkZwavYdNKzjn2raAA+Y7AOIGli4bGUbzMuJKkDC
XUVd9ACZXoBhhiD1CQE4jTeEzLbi3V01BY6TpfqPEYLm2IdievUAWqtjwj5PCxxQo+X/Mpynt5zg
Wc/W0zm90jZA/X9rFYkDtbQP6sIOlu/vAASH3ZIg/4L1xcgqjiOVsPcfIYHNoiZTVsfVuQa1avRp
vOHQIbQSQn9PGyEBKE3nmQrAMioKpGyjkpAAABml6hADA14FGy1QIx91aiysyS0uTmvpoEMixHQp
cTOKB43Ag1+PZ5wfxGpxDoqGRFI6gB0t0rKKHG3+4Ymw0W8XSw2vWD5pmZeX93E0L4R+g+8OoXcA
rEyGt42JakcRGzfb4RqwFkB3ONGk0Fl21KeqaKDB6A/ZxB1mO50c/McE6XDV1euxcnHmoUMNuQUB
CENlqOj9r72PzCLChdP6g6nbXD2aZRKL97vtXUZhmY9MFFTBDTiH7vxkfo1UnI2mGKNSzk7YOtAG
bsY/c84IXIUYXTjLKcvWyBSERHzTIWnSNycTJ4pwI9PMHz4yobd7t0UC/j5v4kiQX+01i1dVwcXN
9Ig6Sw9pyqS14yLt2sl9azpIZYI41SS4u9lTnjRZ+AIpE8jcsKzmLKi7THyeRGKzX+iE2BwFvpDq
KW1tvIVhg/P6JHP9CeepZz7tYkQJXJei70q7QC8yPCWqzvtDGCiZxDECG6zu2/eiBxWKs7nh0sXg
xMbUGeyZ/7nSpSjgWtO7NIuqVXs2XJaBeAPKpMtk87EHp+F6Ycbr7W4cEPUJldv4gns0mmQAbmy6
mpTCx7NorDgSixQDqEEm3FjG5HmPbvoO1KVhQoRqr+AICjepGxzBoMh1OptUviknIE9e6mM+WRPL
zkTfUS34W8Y9+S8q7u50RDR1gQLvMXL1IPo+Ue0ff+DGy9/4dNlyl+R52Ky+dLS2IkBKweBLyLIn
7TsZ81smJCFg5/6Mlds0OvLeU2SsHW9RbQ5Tqjo0Ae5o1wgM1arCDf4c72EiBeNeAcCX81NZM+aU
Vit2NhksPQJ3cC+v4UvQ/SsIH5e7D1zAQpR0mxLVi77WgBCtUW27z09uyU24Zbe60yvxojzXS4h0
OCC0+lNVCv+xzxkG6XsDjAX0xIxt5UgIMh4BCSUr8l5Lhrze8EmRMwIWuGkA8X9Hpeiru3qoQ68J
AkIoqwJQZtXaOaY2XU/4ogC0nLKj4mDFOHl+HGg9MWJ5cb4lQDw5+us2MswJQlmbWmRCDaa6NDAZ
YxTZ89q+7nzSvjp9TNKb/17yvpZrLcTlpZsvQFHBYXniokAHN4zJPjUj4Ir9DPNBVTDnEjX5a53c
F9gyYSCRQnyt9gYVrdFFeNUzrV4h2+dzvRaS6AxnxRnDq6doKV5G+TKTw3Z6kp8aQ8JUxniFgw/A
CsrBJEu9zEBsWDMpgocNCt6t5MyO2Rhv9Eq9MZY0jBM+hjuceoIkihScNkm2rFjHJBuB591SvVui
PtSXKEULUHmk4sZnWoLLKsJRMv6xSVE+9EJP8pEmAPVlHhCJ8QtQLBN1rinuES1kczxz9kcnBPax
jtT3qzKK97M9gzmo1pI6UUWvrpGcO3p1bP9h2Y/7r1Q6CPy6shXB5og4O1nznRT3eyIVnEb1XspO
nv3UMrdFB2jeW7n62kvaVHk921buwCBZWjHEBJdUkRBqx+R1/fajDfwCsH8oDyfqgQ89RJxR2vRR
OMgOl5sE/MA9LbrwUtklZs5UAUIZnuun3IZENmjCwSNor/SBHibmm2DgLawVkc+nSCxFJeEI5w1A
gwKr38MnhIIyfi+YyHaTkIt5qbJwKta7YVvLzJPupdKMf6VgQm0lCktFxZSd8KK78oFdqdGa3jEj
+efdpAom6Lrs3iNyFbc65F/sYBIo5JlRlwAqk+pRxO4EJ3RNVAuQbLHcV9QuyeyPcy9HykY8i9m1
CoOienfVFF29eprowlN5BGz/mxAWoEQHmDxX+61sTXPWZbkpKR4JOMEz3HpAZdk3EKv+YBOVJJIE
bYR0lgL0TCbnX4ywVkdBWe2oc9Ja22a/c8lotJiZam/Z/WWoZJzbBO8GOCsHchfNcE3RuK8SfHut
LHRWmRyKJMtTpfT6m6BFgRsgUcuwBHtxpl6EFnyiY2TEGNfBe27Nh1Byt8Te8s4pTdO4Q98yzsW1
g8Zo3sGbEReZyG8wTRfYfD4Nf+or44VeiTiaPdG2kxYOQ5JizRaG6zsBarXHioxAZ0E9LVv12CXx
JPj1sHsPPBvEyeyLrk1zCq8FtQxOu1x9C5MNKm/L69bLMRFyMzefe9xAFCO9jU+zMqEMKsbTjBEn
iODCWorvZGNHESMYMhgYbE0hWUFL/Titm4Rj+m4v7OaxWGrVeiFzRkLvXFuRtDZb5zLABRCvI2iZ
BCOuH9xwwHL4/0Epuy9CbrTUtxlA4nOBYegm2BO9PVsEDP9NHTtClvzzKo1xwvPBOeRq4duQ+N1h
Z2/TprOdJhLwIgbMVSvz0FPxiALSZvgQ5Q9Qnzl28Eep04wIoGYEw0p7098GMzLNUANctvc/hGY5
XbNeb2lvVtOVLTsfjSJwIbxnWMmoqOgIjQPWpNb2cKnaXU9M6w5J5c2aywZCaUKm5gAfre3kd/Ib
A5LNI2i1GAowgeYugdmqnVn/vvq2NBLcIeUw13YnnhotaSwUUKvN0oE9URLgICnl1cSP0s6xTqzl
oUduyIuUt7VNjGEKe9LoMVUk4ToOneplDWGzwGS64Jtz55O/ZX0oFd/kFzuamlLsJMRY4n5oKHS7
6CzydMHB2dsJaqEMOFev/Z7rIk4Sl4NtobFTk295udPPW3If6EWzZBppO/Z1E8H/pQ09u6C7E/B6
Y8ll27doTYIMEWtSvNweyCRSqZle5e1HdAYPe8BK6UZg9yM6PO8ovnr33Oq2pqa7ILPjuphEd+Dt
KHBu3idxZ8opig5Eb3XkwBuwejSPHjhVnFGbxeKscQRjzx7FCaN3CqZgZjGr4LTcHNVuqM1j79A2
AN0dP4NZ8K1sMBGehFeO9FArNKccyUkdzwMMSJ7RLs8ZWgSNDDYhA+KKGXFUd/KNhcUpW5bjwY/o
Cp6PEELsMHa2EGc81RLjCxzi63tH+VWCkKZHVboqqFttvh06vt03jlg/HSxMhdTuOt+ekXMbwcnf
FsStd8zYO9QIln5TGXXAEjR8l18NXSzgmXQUarXh2dcDJfSEDV8DhKj2PO3VVit+DMJogYF3XF3s
rd3qnlybwdOe6dBzxnLsIr5t7mjtsK6gVmkZH0uaTzl71hNI9H0iZfWn0rb+uqgs3gGahFQu0wfp
t1yGoBz8KdZ/dk9ertV77vyFWHfIo7tCsBcZ2TqyqkgvwRpUmtu5GUupTL9i4vmhRoMqVvVxnHDt
qGS91b4s81+nqsGVLTSEU/IH2AFy1ECSG2AzyvGmCTI9Jsje7RfJGu9L+AABi2HWFYykSV7rA4Xw
QMeP9NgV9sF4tFFKw3SVtytHxE8Zumhy1gc2LIcvS4VKjYUJfL9BmrZumFvk1NgSh269INbtbIOT
kr0EWKjyv08lYwn/qc0bneuI7SrSJFvUL2iDVEm4HT5K+zL/Wx51TMRGGWFSarYohRKzrBvkHC7n
9TB6z8AdJxhvmDW4Eyve7FanN1Ha/MA9r01bE4AKMlNaAc11Ua4Ib7N0JapiHdHm6YCj/lk9pY1O
XhMkSNp8eNghGmH3mQRIXaRd7NyvJsYM1TzhYwZ4UiBB2oJFnmjqMP0ecm3RRnJPCppXBLfhRWJ1
JFWQH1iFmtoRQZ0ZCk3Pjb988pn85KgtDlp69FZGWiXxUEebZulGOGIMMbjpK00mWlzUmA8AZrq5
nJbzj6ZNbpGgdD++QahGy4q/STmW+L85eBhxf7Xa1t77T+BP2Wp/Jzna+DqSbY5/Wfb5us4Ims1g
1EJ+Whw0aOL0QInOhS++jr2z1tbiCnl7kq03MKO/e7Y0NjKZ6u+PKyiiM+9R3TvDpbajBkpM/tuE
DJ+S183Mo8INHw6NPxeqPRdviXM8aPvVuFVHiUg7RIrivvu5yEtVdzfR/d635Vzl+sjaME7tTFqV
Pj1sYKX1KSqjFkCuSNbj8V9+M8MhTEfMYDSjWYkkD85dEP++kN9r1W9X1tMDSQCJQWRNYZ+j+KNm
Sq8I8zbNbtR8Dkp/hZ+JXmYm2FBSW9yo+gpA2wzHrDggNcHbLaDJB3TC2ocJ2cTLKv8kFtaeZaXa
j9MmExQ0Sa5S2nzA3MQE+a6niqCyGI7k0FX1wKVCvR5H+NtaAjO6XarsSwksGWHxM5mlC9chj9rM
UG9Qc2iTV/GcZ+4AdqzpwJ6tF+YTwos9LRnrJTdUKT4PIYiGdiObm3JWYCDnlnnD7krkaolWNNRq
tnQb29s/QFlBct/sx8bll+ZMGOXBSKg5bavpcTJi+zRCrrF6W6xVKbvqVOZGqPPwSHPqjAnjB0Bz
QU8+WlxPaqzx0oi1PqF3ooAgEUWia27lKlx7uf/26AUFIOshPgHRA83AxwZG5Ncrfkpa+wsamHkm
2DdFYQA5idrwlA0rD8e/1jgrJcIyfOPp/N9SQ18QcDq9+V7HkNrYovkfUfVhwee2/ZLAdvtk/xB4
QqtsRev2+mnr+wVJBF5KzoxNGER4I6aq58KUEHd1PgFvKhhU7VCsRj9FBDxQHjYDouukAWuFo9xu
pMOHD3SFSrdmtMbYl2myMFfEkghHqdTvW+CBTJu/UsQpHSVii0wkeOa5EMYO+T4Bg5KL2RWrToeC
hT2ahhC1xscFhliI8UzaEMp5isrxM5vPHXNj74RxO9G+qHclMlRgMwSk1Pn7vJgQcjl60Cxh93VU
OtEFqqK57N6ECIXfubvlLsX2LFAFQdk1JMiMMjskfZZPZ57uDilFgLMU706CSSYIeY6AaWtJ8mEe
U9+yCRqqvMNDUCnhv3opAJo9RDK/+m02MlVo/g31KyMUnqPa9PGj/zoe1lB3vzcUtZ37Viknu7v3
Ogfzqn9fAhOqW4V9LDBUhjeOMdmlMFeUORPisKzZ9vE/F5NmWSZOHV9t17PFrLXEJ1aM0caFOJ7g
c9AQlR1s6DQbmldJzpDkHWYLefJJ/xCds07KFhxfWV4ExYEmw7IHoFZurz/Q5TYvOCRYdLtQxNzq
6EgZR/rYeTj741wWnk50NzsNJqGj2cfEpqWmw/PmfmTHoTXu2VjjbIbBkIN6ugCt8BU95LsrNm6K
wpaUR1bRHUaGmvIkS/Z76NyyqDd8JLtcVmNGPDaz87JPKIJt23hBHfyBHdX8jou0EFhNtn1V5+mg
fsFwkIDpevnK8GSGakOPMH4FLGyBd0PsJhM0SWjwOZBtJXvYXx41Y7VlrWwSCAlLiqim2QW2KfPi
+7Yi9clr9jsfJoX6K/OFmD+CmBB6WXIM+zGmKyEv3aL/wCddzArkMcghQ39a3VZyRWvxTlb40KmP
H2FLSmSU77bMHIb9e+RWK/r/TzWb0JAC6lBbKS9E8Ck4NaXU/KiBFrrteB0okfSuEKP2/112tsQZ
7lMM7k85l2ossZToRtOuoNd8RLS9yPLbMPWWVXl3NF2XP7UKUIFaOOHM2swVZ9FjjOimxPzQsiZa
9OOLx8YXIeZnhX8imll3HrBOJs21Kn2edhZs7lU8xRebLla8VeP75jR/am17T91nZIoQBUMy5O4g
pOUNZHDdd7IRmOO0939eeUjDDeVfjpSWgoMafcBblzfK1b5Nc3o2l/rwGEnpMivPhRULYXWztgT9
540oWyj/mi/jISa4E1SnzheIuQ7y+L2zfqUX0bw9H5SyMMvEa/WmHIkmqHr93xeK+OUn9kt1GE2M
9nJ/1xL5NwmFhD2W9IMlDC0Gu8/LAaoVVkNlNTgI4wWRVE+ogmf41w2MgDIqmq/zCOVwWDGiTWSC
Xa8xcZrUJhBVRYoVzGPkN3xrIlxF1gC8JYwKsDrc7LQoG6TGzu81a96WvGORkwiC+vsM858dHAot
aJOSFIY9V5D8WnJvf0/9/1BeD5b6TmYqoPOHbHM0OchsnwFkus+azQhWXTDcW9lAmz4LE5XM3A++
lGCuadumV7D85dkN6Phhf9+it3zeT5gnSxrkQSyhO9+YOE2ffwRFr8mm/9bXtqGd/h+ecE5Fo+Il
QppZcH23DYzi9oRP6QlCDGQNxDc3dxNmL8lK82oD83gncCIxMXTfbkH1rhmanUxnzh2yTyJkvmhs
vyebL4c4FvwSyiIhMSJbVX0HmDrS2x5Dp+idnxz3BemqLd8pVI1hMO3U++ZsSdM5D4vIXJFQUT2m
S5S9+4igzww3AhiSln4bZjW2LpCnCOlFyErJn5CuMPS78N/bqnSzJMsAb+JUeO/e6MGqBM2nsgHl
15zw+hQ93aOZzeV+JUC9TZ40BagNMP1cP76bX33+H21GwcZ+0NYz7dDe7C9Z44zLbcqra3z180yu
fyevFkc1gMNfSgIJKiWP9ShSLWqsCmUOcUGBRdt3mzleN0/I+My2Sw/O4oSkkU9CJfsid4ocGK/X
f2z/B9aQGxkccM00fkHw8kFEpdcqXg/unO4p4R9AFJfRqftNWFbURoUhXbt9fdN5NXI0Dc3wVbud
7VuL+DBPaAJ0hk3S+Ef0Mim7ZfDxMYd1iuc6YbNGgyw/T0yfxUV762qzMBTIZfuquDim1cGdn4IM
12MBPTOLArUrDH7oUk+3HgmTYm/l065496nAXnuMCFE8cXW33v4zL/0jaGEUaWOFiWxaFReNlI6v
L0ZjAxqqZ5lYUH2UVgkQSzEbQJ+EMQG5p+SJEduyaQT50FrWl1Z0wDX3Hd7ig1piPyUNDW9Sj9/y
lTJ5foym8G4H7qBc7LeB3TdFNv/ZTRlhaApNNTXlNuPvMeOXitcy0e2PyhmwXv4wAZqgSL35oWYA
cLBFrAHE2ZG3TrqZOt9NDNKP9TCoB2G2y5FT+pm+b9TQ9u6UthiuEj8kHtQ2wGoGLjC5iioxdnir
75icPywLPyhIZTmjKN9+0/aa4CBhU+D5ESjQL88xMWZA/vh9OoLx2pAOgbjAPj8lr5+kJlM0gURF
40UsSbANcAZxVuXUiCawwjfjjfoFZcm8qUdArNU3UCbRfdl/3eNWBsJUObz/Mmv1G0/SBeBCgEFf
z4l8tX3ue1LhvDUD/YL5LAM7wFCSsm1UlzvndsgU0raBx4e3YLUd7ENpNoD2NZmlqZUtmPKlxhn0
TRjz9d0ctmb06PAfupm+b9temvhTzdH/IfOK03b09tIfqXpanhyHzCmOlzt6l37qT0Evfto3YlNs
qVQ0B8jGT2wTmMHd4tADMHoGTJXFOkREntF3eCcsefsHAzX9sHQNnoEAPdnkvW8THa2EBDbnj7rt
NsPEhVr+7IIO9yLTepPj6/Kcr/TFkBxWkaNiaj1CAuC/cKfNO/pESFLueYnsodB3hMcFnFqNDYaY
pelgEmelPpS0pl9Rv74x9FTmzHSAY2AiRVTZGPQsdFss/2JAZ8POCtOeVoAuAfrJxPXK0O0z/zen
45AzV6tRILRdiDbOYfl6TPGh2lSv6ywegqw3FjAIv7e5UzqWBBBsfQsS2jtrC6H9SCjB9Ou/z71j
epUaDArGhbyBkCcCFLt8fPYMSDOBw2dCPQDyqpsUCdRLsACS6qStm7ETd0stnbfnqE6hREeXf468
RJdHFZ2fqFxpJTGDukVkcSMnu2SPMN+p1U+tQftGmhYFrCX5/uarYsZgt69dVvPYIjqfbWjfRUhf
Pla0pChPLWO/HRywSoVF8Ol6hIwr1o/M4WyoawrRMTRv+FpbLr39aUGA8SwZDv5x4DQb710V6DEQ
y+JdZbLJHbg1C60U0pgy3NiT5D0/PUODlZX0V36tHeYC86qkSp3V2cT6vzYeqb4BWd/aCgFDufOK
Ni9oimRXX/xkkY5FILfmDXh86lrVXGle9TUVd8EGCgE9De4IpOHTAODxSQwgWTbIBdIela79IlBM
fq+N3RfFUA8F5/OEjO81+Rscp03J4zWHkKPnObuXPFzJLAJk3fordFulobalc0brSGGCTY9zn0QX
6sTvqy4UCpbaxV6vymhJ5jDP2OmWcd4mgJcEbkrVWDrjV/HE2yjpi6daEwH87zmPNvmpjLzXw4jR
GYuwKmBiLIUlSzZnP/4z2dryhL+O4jsTAISjTSN31TR8Q6whRjryaKXfgeKVEuhVwuZ0hUsDRhKQ
8rNsrgwD/5X7SQDw+ci93cbnBCxAQbwCjWlC4tfhiZwecd2AZZP1ShtQlCuRJIPeihI8BFVm6dSj
R7B1Fd8a6mm3Xh6DECMIy2UVoyZ2totiMQC12hW7nZzj4Sf297oCrCiS9GPw+V6f+KQlUt8M4xrp
iE4OaYBDcPsUUM4vffNIY4DS0BlcZk55RguV1tezMoo2fNfXB1YHyGMSkrj/CgE4xVKoRA8o2IUX
YIANLPkY28bLepVU0p/5de1YqLmfMZAkGpYGarVzDXMDbBBeKMmVq2qAMMCWmreNOCAAsiPCkxal
bjJ1wx3YdkScXO39zYQDIlR6xh3lP6T3x5TJHOSvC3Smy1/iVB2d1U9KeC0iXN1dxWsna2U7XDd/
+fX2rY9hZVc4dKffolejVLRlkwtpwdJaJU2Lz1bsz3A8g+uG4RdmQr8anD5sPXOYeb6wn+bnLETy
8IzRATdiFkAeW6NsutaLdLBZcNmVkT9m3toA8MB6seCz0Btc2euoY9TP6m0QaXxXlLaBpKBdr0B/
v/YEpQGM15g5i/V5AQG3fNjmvEjP613BfdYOXedWUpzH0QQLkDqjSqD16icPH/SrIQakpoemqXgE
rA+aOLK+7SgkmA9x3t+cH97YbvKm6vhfGfCwWenyFN2/Mr1s1P6BW7bJ+7kjcUNjedMP+I+k88DG
DxxUHMT/RnAaIwRYFObZvTJterdks47KwSsQENFasSX3Rbac/aciKeWxclc+dgE9uOeFp/drZecB
cmXHDkqVYyzAXUWOZ+s5UfmBSSpMKd60tZlKHX6UkrMU1SxB4imX7fDLx5WVia9R7biy2K1TM5Md
hHv5FeFCgMnlBBA0EXnRmpGGGL/E1CzHRpTPmB3IpjuiDFr2UOlT4MIcRJFtrtVSIkOZZkoXfqHw
dGILyKkgm0CamAOs4eerNWqoZZlKUANa3uVnLkv87DSwY1r0h50g/2yGPKpzV/Zsm2tZG1eXd045
mA4rvYLPub9gdF/axImNplveeNQMlaHkE2iKkj9ftHdgDpS1hJ3bdOgEEg2g0/v9NhnorJuPWFu5
Ba+9FOOGpcLhRrpYI7ezVfX3VmP5gly2so7a3oNTenSYwbn1ogaFRV8ANfSugO1fAKlmkV4N2Vzs
ZQOiv1KHwVBZRaZeMu6DrbkKHcCcmURmj5wjCoK23bdW3SEA+ZiKr1WliX9+YeSfVjIih4RKGJ1R
stl2mgyDuFNX4ksO/MULBPduVWm3ATrwr0/sSha9ngHz/XE+p2F6DUrcSzuJSK7UZqPEMpmE8jwk
yaIDxCOzqDRaa2uu8xZNNqoMMDOhD71LcaUtc54tkss2W5L6lO2S3f5hsvFRp3lJHmRcMk4+2k15
/Xywv2S2k3t5m/hmxfL4dFzYs5bCEFooum0+H5IQ1+1nkEpZtrCHF9fgM7PyIMs3Db4HyBvUyrK0
boMPtv153xH0by5PwnRT3AX4RVPNtoFyQLXGADrVRogyMWzoYxOPjkRdmY2YvE7OEsO+FB53GzMB
wWQY0pejVKM/1sIzUn5j/z37RmEhtBoGrMGV2pLBnmQyasdbeVnOD0qGLQdNOkYGVzqrmB/THXnc
VgS6dh+sSGM/DubNoyfEsF+ngzNoU8FElCR6Nmqph6QxB9Wu02PSFS0msXnvYVW6mlTXrUOI16Sn
vybnpXQyu9s8R4dEzJSqS7u8Alut7GY69HSwOae/UQey01yTk0zHfBBLocEFadF6R7F1cxJgCEEg
c+AdePaqbAKA1ABpzxDXA2B54Pky5cPw4jXY3I3W+IbkUGgCeWQB0P8O2VVC815z1qhNsc7WKtrV
s+fhiQtZ4bcoPRDFeJflVvtLWv1YO59TeN7NWHIrPnlF8TSy0miEv7nrAjBECzMEhSRHxRnefEx+
MwSryC+OI2c88dC28J0nvQBLyDbZxrgrpcMDiPCq2HZPLZB4M+O+bEnYklAZQP8WzAL1QgSVYJU5
fpvYn/xqQBxZ0qfoitb9vllspD66XW8wGs3eudwZSTccfoTIgtUGbx/vnwikIHD7UnQBuDzaP+VJ
qZEzrKctcG2XlFYmNI9KGkJz0D9rWYm1zEqwLZnE2kH+OnE6eDmSXn5GVqkVtKQVYl7X3EAR2V1g
n24Q3MzZB8qS8WJzRi3N19OYP2Gyti1Ek1timvUzijW7CY8lg6wKeySJ1I+HTF/GNj78F+yM5KtM
bnntp2rzgjMK1rC0awMPUonbH8XZfMKw5W4MbH0gFMZ4HWbJdN9JW1twotjaBNtdYLxBpE+J8eCm
ZE07bct+uznzWez0BnjTbAyBkGqiHJMRpBPZDHfsPM049r3Il4tYv0xraIkQgCe5pPfKjn1Dd+Io
kqzDmq2379MC8DANhazx5HUioHATSkDKbT8dYckwDbg4vAkFEEa30keEQdfT9H95qkgBE8QBqEPw
drE7Dr7jj9D0U7/k+UxA36guANWosVvgCIYsctuBfk5+u9t0nXknrcNfO1uNYKL3TxKrBCiwRKeV
g7ppgWBudIatfX/pnT8JbW9bIiQKkqXceFe7N9/wMsGYyJ4+LReigZtk4Fgb1Vb6jWB3jnykgJOV
dO5G3pjhRUZBBBR9SE/fuYdShXqn12wCXZNFeYFLqkRtkEMA6T0Fd1wj4SecFi8rzQuKXmgBNAdz
gGycffYhmvTqUFpSl+ydD6fFzB771FAdY2y9aSIo5tb0piiD0yzbcmqccxMfMgxktCGH6z+Yv9pW
W6x8vgg/rPhnCvy3bpdojf9ewvYukIa6/0IjqgyzW8/li4rZtiLE1OYuRtWPgW2igj5HhiJbA3pk
Pgn1Z8/beOeJQY0QoB6h5TpP6w16gqKTRpmoIr7fAeaTOLx/MG9CY/Q0RQb2mrWfgsTfp181p+vk
H6TLYBx2vs/2wSfAjlFSEyEzG5RfC+V1nrqCMf/sN/u+9NqYUDYGQVfIxXPfLy2SvFn+idHG9Elw
3ZefVK3zVom+LgGl2Z3jCEQD669jPPuVDER5H2OfUJpqzWYeyUgsAc1u9cwXIG4TrNtG4qQLOSqA
FRKIzXa4A2ToDHlxRVOK6wPZnM5GlOq8AdYBmwuej1HRwuIFRC9baQgcRPZw4a3MJwZCzKTdzDew
uwNlzB/+GT2YeIUtorJmfcJnpoXXwtsqq6c6N5EJDqF/PcT4C9aN4uUKUVzcoBRamepe8HucN/Ot
13xZ760btP2wjcvjZ5chMVb9hfF8d9u1HXiZigz11DhXNgihhn+JekXyGol/fP9My7B4l8Aie7cO
bxnjWFDP9HOoizBi3mtFujjvPW2FQ/UAcnYThNe9XuG6XD/1JLSchRRXk2YbFOR3C7hfkVIsVZPv
sVXXkz+1yqo+qR6T8FW4D6IiWCpKlouetWzj30R0ygzE0OI/CHpZrTn3wfL82gq+ClakbBFSHizF
LJ/AtXMoWlHEvWa8ScH5aWzA0AiUGC9R22EXQleYhWm4xZ41Yda0WiTFEdXmbh8aoOj/q13JULh0
11j1ZbMNU6dTniH5VmUg+P0eTYMvtQtnD5ST3TJNS6/outBXadyKcpdghPVYTZfdlEwtPf2+wNki
+7nxgJvaY3Erd8EIJ3akLoPR29fc1orgwO4VBXGU9hcvEVvPBrPE4kZZOLOEskSvKhGFs3cgnA+r
HRJRy208izL+9JtVIZkcj+5mSkdcfNhum+xbWGQ1bFlV/DwIl6c7Ot/L5AiohQqB88l/1C51F1nh
yByNE7rxE8rbC7SnD0YnlAt42vob8ExWW6dQHGMozmCUJvCyDmgSD7NrSLYQeEptgTdlGWU+9d0F
VX2ylnJ5N8l1MzpVSqqeXtyTkD9Qs0LRCyvU9QdFKzA7AyynwGLo5mV0eCduZ+zyHNNhre0kU2LN
5+wScnXWmG9SjTiQa6ZKfR//NvXx4z0hmwZJmK5xVQW8Q6nl9I7qsOYyAiwhTubGJ9MUhMQWKIgc
Y2c9PuC7ntUuGub4KY5Dt2sp7E3y/gvkk1mZxSyPqgvu2A7rFIcvuAmSZF+gUImENAedCvrLAyuM
T3AUP8Kri+9I6zQ4eOd9JB7SA/hxYrj2dxghD6iT893dPHASSSEM+mW2999dNrvbVMHG0B/o5Bh6
TFfJpcUfLNC19EcwCrbVyqsN+H8wMepS1If3LdsISlDiI/Ns38QcM0aH5fKKA1JZJk+hO2YqRvQw
0q5fPHmtVBdBXxBtXvSErXNtlV5EjZAaO/AA4LHPTT6xWupZUZsjkTeuy/YvxvG8NdSiimD4Q5EK
LLwIxgqysT6E1NlGU1InbIfRVmF58YJCeH32TdstdHSUmJszRNjWTmsi0kBdoQB9Gc+EoKXjzyM5
OSrwIL+odt+GcZuMTzYrkH6wNfsSqLwWZ0doBSXuIBaSJbZOlDuHyJNbOHpboZdJ0CA0JY/BybM7
IwGlbS0MBw7CnJS3x/3gyW7TYt4fwFW/3r6/YzJSczA9smjsYZ7Hb3HwgPZ7w7n7L4GnZr2PSrCS
5V/3unCEP+UAvl0zJ8k+N1lPp8DZ3hIHcm1lFIjhRSHwTQy1aPqZzcezDAjFbdEq907tfY5G5KXX
BREmGRAgLq/r78d1gqWQd2D/TKfAdaLR/4fJ1wERj6lNC017CjvdA1XJykBR0lLlk19LkxKI8yBL
6xHyZWlxNFRBB/xk4rXJzXj44+F6gTmpDLcLjicZNSrQCV8YpmKlYcxhfIJxRFUyjnwShE8kWqsL
YO63Y/O5egdCC9XlvkJtomfPLq3XpqOhc0ewWs7X0QoSIGXmYiIvf876xIFJ7GZyRhrtZ+YgTnQq
++JxqByeqCq/cyxnHf/1YKnvdFOUW00hHzHumk0NZcyQdl3KoWNuWmxdsXiYlUVkqXPTXLJQO7+g
dAoZG/CrZ/ppYqhsb5TouZvMXlOLzZXOsZdjXgd6dbdMvcgXohWcpEjPWgb15BCFuNEzqQ/zueyL
hYNWhKWI7U36R/M24Tq5ZAAnEiXbFkSNsMtaQ5WxDsBSj+LIiOB9NXdA/og6C/a5viUvV5Kpw6S3
xyF/0+1rgONbvdpyXlGopo1Y0ZVjbLUhISLc7Asu0ZQOGRzIvl/fXCIvyTp4nSDccmSWXbn8pZdz
QDMD7nsbC8BsZWZGRK0BL8jaKvE7gTCqLKPgar8dN/LP8tFHQxnk5Q3nRvohJOm95hF1uRjhuQJW
bqRLE52alEr/b20EL/v1EkEWxvmz6zT2fTS42iz6nJDY7ohxzdN1vn7+rRw1dFeg7GEh4vvMgxTX
dgTw77hFxnjTQ+fBqejQuepk+GoHytoErSP/xs5GOj+jpeDql9ycHQb+QWzpob0UlJeEC24nB7+p
sxh/mbCjcaqTjOisEUtfMiLq5sWYTFxhXs8y5P+tU1Mp01UdtszZcTb5gHcdLCrmWwBHDDWwEEKq
FEvC3bhs+72EDz4lzqRKvWj/PkmEgCg1vgm+hwYfaG8vLVHaMy8uwQjIScif//2RBkdHYvZPL8Kp
f2pij9ed2OZ8iz4VpPzve4ZzB2Xv3ug5f4hr4nCx7o7DRV7BNK7tmwfPiowgt4gdkqqD7wQvGbzm
IkOYApjZAJ7j5w9F60rdOOxMm6EXq+q8xCOLYBSCMlF0z4fZRI2MHsS628NpbsdVvrJZekaUEVOy
MKhsF03OEvszBSLzCgEBFtQQa4BxfqzFnqjFiuil5OT5Z2+ADbTXWAWVJ0D6YdIq3tz4Ym399hB7
umZlrYxpg82OzTGiHBMc68CfpZtR8p5FzIAIODixC5c7SyB5KE6MZdnJqBqtbGmINwJ4U4VOGRd5
4SqBTYlTiB7co4IxPjgZ93VUw3KSWjw9w4X8I8pg2TwqA0sYTdsWm7hQ9SZevVN+V5rnDQR3pSch
EPTqdHyqseZvy6v4CaXemnTp4+r4SSk5jUIVuRBIuXUoQid10kGf3vUavdqQsl1t25UBATqqQeNF
1jrPZIeARX4BRERUF6yxjUftPpjuAPfFt5xPwqpL5IQ+1Stx9u6ZL9dVo18uOlhrmgKvxth3nXWC
VWw+XDRIrn/LMylBP+YuRwqSDUKjWQvCxv+6fdQdTzcj97Pfyp8Oy7h16+bdKv6ILVj1pOraY1Ua
lMp8x5PJMs1FF80h1STWlMOAoGCna7o4rQGI2Via7W5P/xEBnqto31XRWGE9qmhe/Wc6Hk3Dcf6P
/0YwV2v8Zo+KKCzlS4fHuskrLKkbuhgwlsa50gicCmJDR2sFOLCPkxW0HYELfVP3npy1LjpI6xLp
4k/mmhRTjUl8GjxodS30IPBTjqoWsX+Cq1w7bo7dN1W3u39PCl61Po8Su8nnbO+AwrnQ/yPZOodo
tjwVsmhqouj7D+wz6ae849PfkyCobEpvIK2bPtrLOzjC4XcLrd2SHmiSxtB9wwo9BXF++96w61OY
5nTWK4EbJsabTOQoRxkXZZbSIjEG1hxo04kXvzlk3lOfrS2JlnWR6kojhf+Gkqs/vgltCaHX5jxp
vnutBxofeV7UninzAa9cfxUPAwM0VpwReoRsUXmA2E0dJaxKU2cy669SpmyzDD1smJJgtXEz/rXZ
7KttYdwr5liu2omn120tJvUc+B+SWuM6OdeAESRYsMwcMJIctkizNBsFULmuCoXzr1c6IjpZ8Zym
9d16tG9LKB9K/g0TCZf+1mAR3+ditEZUkkpHw7hlaAGiP/xT1MGmyIXQNLFxDsvMtu4x1i4jTK2P
AD511nayVKbrF3d7/oJRcKYvzVsNbjwusXQYBcZlvzqx/O196i4HlJSLr4GAhZaqTjxw6v/Exqip
HYzLI/gShTpGij7WWeTXnpfvBQ/Vrkw5vWoUFHev3isJ+Wk0Ay2zH56pfUiYzKi0R0jPHOQ0WmaH
mWRoI5pnY9XYuRK2M3azGlfKhEG3gP9KayRyuP1PanR18KkiPigPTD+9ltVqZoaV66M195H6u/1L
9gkti28aEHtsHi45Q+WQA65jBNclwcuIpFmE4iwBq2UgBd8ICr+ls+oNZBB0I3GBPJR+r5yWFDJJ
GyWI6Z/5J4F9GBLMmTpu5gU1hzt46qRZlhywkyjoMIf7IgxCqhuhYp2bVJEOrwXRh+ue7vUZNmC7
lNf+d2Jbl9bGzhF3UReiqoDG9nRYS+/sj6V3/nKg9+KediML6Ai2S1U3+msrkJKHgDh1oImS0oEh
FPTQ/p2EHzfT/OWxidBM1gLAjkP81oB9wr2MIw2S28+6r67ZaQT6w9Aj48m2o34hM8AG1ZrZ0DOv
cSXLYmmHd/DcFNHsdeoFtgE21EjwxxrN3E7U1QVhuqSvSM12sl/vCNRAn28M+2cuuejnOSTjqCyX
2VLYZfgm3i2O4sYB4xOM1fvoPDQS//HbDRrUc1WVrRCy71EuSY2GQ6qipkrVsUz9yHhttmoImP79
wEHiHFfuaXcUmwbTWOAtnCTQ/G8U/BjrgN2Dwytl8/WhA/QUeA5sQ9VbVAF7qhcVXgjisbXPxG8f
RD4ANhwXwbrrBPg3oBvwnsjbBKyBvQHDTDa2tP1zTEEBDG9umhCIEyfuYuER+Yvauj5GG2avROuh
RpJhJhM+1f94vS5HiCfxbD7qdE+cz931sG1vtrGlRLMt1+jEQ33jfx9g5Ngtq9cw1xophz6EpggH
nCMpbGvhdmJ/f2VoDnQMrT9mIN3LcZxygc1HCc6c6km7EcTOD3xs7dTZjhuKhBBVrsFeS2Z4Bj4P
w+bfxg5hd/6ehLd8B4iv3qCwFCqjnU6r2f/56rr7+N5UKElGJGxYDkTxo18hT4cqr/f8YbXiN+/L
ErJf60GHeWv22bsxWAgOUOnKWsQ39sMtBV24z21nvdexNwsNSxVs1cNhY99fGck6eE8QW6CJTPwZ
R3UHlV1E+gwYcXcdirJ03bgXOcHj7wy+IYRHaKsaE36OMwfBSe1WD14hyx/xsXLpkO06CY4SQEbs
2x6u3PWFIgOyI/p3m84KLRLVTCyuHNom7JgEdbK9qrYIySi4ekT7O9OzoAEfAO2Xkvcb/sBc1cRn
UOknHjG3k6bsvI/iV0xUQLXk9rkqSvwv1Bw3d+HpKeCZlDzsbyaf0RF28vouCbEtakmvCpu73oT5
G8fVHS5FfMm1WEIrunupCahR7e1ViOrOrIljKXkXPM/XMwyIeUC/sBJgE/uQH4oyXc9aZrdbA8Gh
arGFxFbRKnJr7XubGGk+n7S3NBqfZH1Ph589kwQCuREJkKARknBEJQDN56NCO2+PDU1FbceiR6Md
HzPD89YHeYdvdLlIn2m3g5UNaTceBxAqougtH5bnENlvC+rOkgSIuvjMw54NZ3dpeUWNjeKFA7OU
kc1p+op/spp9JYfVhDGVAtqu6RHh1WLt4Bw6aS2rgHE0Uyu89rzyCOqKDeTNr8NzWRPsJR3d2Mnd
1iB33A+wKd14efvJsNhunpp6PIeaR+GWfftcMSCe3/sKjSK7Xi1hECrGmuwd0C9e+vbLCUBJG9UU
tAY3ws/9ESTDHTZ2X5T0Heq+FLgP2OamK/JAdy15RJh3WxPQ3OqGQ+tSBZkjsTbZud0VwxKVhQzo
zo8hyg8jU46R1Iji1Pq8Ce+Gprt/ZfpvStDj2zKSpdsvNiEpps8opfSU1v7X22vA2N0g9OdjMvFl
b6W5kbVfG6KNRoGA9LdpsUTIgRaTLkLJizKY4tYKIUPA+zscpvY711Oy8IQJy8KhkPOs77w+mQ43
x+LuCWCW1y9C8Y/LrZ/neJDm/5N5et5FMrRdve+B8UNX4hqyQ1CZ+yWQw/RuoZkBlBya8eYkisEQ
muoIJmoeik6+5+kxL1iWldVxUq5RTFMCcQQwwgs8JKNQRAZQBr8k/GRtYCxNgt/pGuA3bpYsTR5T
rP9ciWl8PftLAq1UZAp3ORyirjAqwRyTOM0WsYz6zHInoffSWN7/QqcurRhn5fEbf26ErlJDr7sn
WRNbYSTRTZ+8467S7d1uMtVMe0UAbZUbaWymtqZiB+Gi1VXpI5GZCjjbY5l6CcemM/uxFkVnI5D+
5FZdssW+QZgj8Ak3F+UYesJnHlIu7vhhbXrid01WRwP6TRD2mqCiIJSYv6dRDb6oVtiOuCrA6zRv
6uCyPBLsAjOPHXADwO4fx/B7Jid3sv8RUJq903toS0L7Q7oTZzeDM6zAHVPcCWQXFHxevrfBtD+t
FQnXlvgw7fwmzkETMwc3JDnXyJg3Y/s8KV5sx9z4ZcLL8H/o5AIWVAkeMWbkbNHUmq5qujUc2/3l
VsqPXVAUFn1bzB9gTFFZoLIgalOgKVEPXvwvdzJIdPhcpAdrr8ywxvebOg04RkLfkENE7zJDQCGk
d+7WYacfTDm3ABP3iur0HfN+O15ekUuor5hmQOf/UIR0Yvb3NWaFjWwI8uj8LHKh5l4knAOFKBbw
pnmLyBZvscKG9oj/FCPWli8vshnMC3MyUGNbGOSttcsZ6A79HjLp6RkQ3EsRmP3k0T0wZJocq6Z/
65Z8mha6nuSOhdpdvUN5Ty15aTIPlcrpJJ30LmikbeN+RvAds0yYqjMXKaaT0B0oyhvrSQMWWaBv
CxD+LZfPnmrS6eOskRvtgCZEQ5Kjizsob4Gafu3bgmlUam53JA6j+APCBUrrQ9ruDdEGPDLTSLqE
Q7lLMnLVlxFK90HgcgnxCVWhEaiM+QyA2t3r/KlAbtxqXs9GTimI80+FxgEaVGS1izT/8njCXb/I
0lWF+wKFBC6wr5hl5j4gRv1J9CB0EnmVLGqHQqiLRhEGqaFCgxvanoUe32utC2O2FnwVTiw0dT3A
bqX3e06qHfRZmC4eDxBp/0u/vtotvxJbWXCVL88PDBo37JXYGdcFFQdoMrJMxWqhnSBS2zyE23lZ
1cXJPnYYc+LMG6jYEiRw+XfeKT1d41iBFsUDEbzO3CwbskBFSVmPdDUj1mEqUk+D4WnLw+nCuIxA
xxgbjXhSafu+YWY40rrvBjy+R74ubuilh0/4qWCOMj5IGOYQjQ7ubtDBBJvYRHpmXl1o9nng7PFR
bVKijMMTWkLvqRoKj4SscCm5nYVN9chIkY7KEMHmC03a7tMos0EeXuRPQ2Q9cAGQggfwyBNfSxWj
MNLakD06bf0e4E3OZ7on0+O1ThFypDBgn4hl2KH6UX2Jn7n6WIDGgVMnetetokUMnEy0FSAp0n19
7vMNKlIVYxt9QD1ZYbcKZi5xKSAJweODjpQLtA04lr5lRy9LZDuir5G4c15u/HybzphVR1LGXt6f
3UQI3vLdlScmSrout10Bt33jENzMlI3lbFubj1JK9IccwbOkcEnhM1mzexyMxSoXYssf1TlWeq7E
ZSUtirgr+F4bTyw9xkElHzP2PKce5MfFG5QxDthreeDVavnx8lhY1vFi9vddHciYbUyJJ88EZoUK
w8n0O3EE3V+zQrHp6oib4t7glzQ6+/unxUfo9RuGDBR1SQneai05wAmh9vYgwoRq6n0wWMju6z8j
AnslAb2iEj+2xXGArOjEKwj5YVE+mFade3/vubexKzqrTHGc6Y5GY2CYB0gZeh49fE9tpCowgL8g
9zh4gVu9wCbHNYk1LL01ui7SeEUiyMdmHkAB2w+MtgqGlZFh+v+7WGX0aWAOcc9IBoAhDRvkhgrF
h1/QJ9cY/3skK/qodnhUXPoxSgGKn8JpOdK8+quVPczX83sZhuOH8vBb+CgxrAvB3oWURjSiVbnk
/C0W5zN/EjLUmB3FNcLl6OverZXDsqLplqiMfpZh7fvH8ouc46V2SIqdj2bsZe5v4BEdN0fccUbW
CIKDANzLVQZVFc4niaOtiR1lwhLrZF82mPRxocOf/3wPE1cNG1ryzffJUhBDf0Y+OgeTRGFogBJ8
0q0TltDSiy67mPcyFcYWyvU5XBCWWqrKfn8jcF/RdgXaX4cthn5riYkA/5wjZSaictfEqUDabq2f
U1pt2+sAoHdy0SZzKaXytK/PE7nhy/b3C/kSgQWGZ8Gi4VURY74Riyc6K8GHBonz2e0r7n1gnLmg
hXYiSw+eW5/7ApRQfKTqsKgxfvHZXXc8Rj+rfYt3pz7Xaq5HChIPsQbdUkEfTpjUgACtQrsuKd70
zCUZ9/3CELQfhDb3AkWEZ/gW9AddiEGtwT2dqnv9H68W1AeeRgfMssnlDz4a2Xea7C4l2oG1jIfU
7r56xGiAAb/7XHl7AfDecvWO9rMnY21RFHRiW8CExzncKCO1B7e3piMLYSmttevC7SHTUYfQXup2
CjgO8ej/L0UNiaGXdYEedjnC6PoytzbvCvLZzKdj6ukwxnQJLGqNptp2nG6CbISu6umkatDWJias
JbUmJueYkm/GhoHj/nfH7del7kHcVVUgV9EKGbxiRhQIOWtOUJ6S2Jpqwx4Ibf8LIg00EgWTtDLy
TZTY8PN1+F69nj7Kjh1XZRmONQw0/12V9AKiZw6T8a1gWKV8UXyzTHZu00Z+J6m9OWVCiJm/DLLg
ay37UPZzi3iv4KNJRycxfNfpVf2XRgUaaEVDUFOYyvbx6LlYDUBu00XRtczkwHLUbVUykdqA+ptF
AZwck265/pLsbetHt/JCU4z/JrNNv/5lY1/cNwVEV5N+HyqkP6SVyUABMwOXAyMxorne16hv+mxV
q94jiXJ1eUSgJfP7mXVN0c63ib7uGtPF0qqchaz+2D9nQbuSuTp99wt1zBsnplrgX/8WXFgNh1tp
6nTnzrzrl/RNB9eT9ivZqETiLNO71z2f6cfM81VltMqjYpY5rHSo79BZbr4kke0X9ofPfwkHTExb
ByyzFKKIQLuLtiehOOKBzPqlhQBZs/kC0Z7oxytHWH/1v83wqLV75UMwn2M2zsWihFVufN7fwZp7
L8hbCWeesgEdVimoxGZKkLbvKq+HTjbAdOOvzW5p57hYcNOKDUNun6PcsM1uX0uwGhobZZiQ/Kno
dsQEnaT3cwErCKWCs9ePy4O4ZTsLKwvPx5Wo5rhgaCM2G8VLlGwezOEfrZodCcNW38taByGdE7tH
h/LB1DZnqv3n1ys2h/JEDEzX0ixHMLQNCKlQWcr1MpHkrrseqxDJ7XMkBpZgjumSJydRDvyKrZwL
DaH98YhETojqjAj4jKDfPB9PVTyK5Kj7CHC5zmpMBm49CPyEWDaYN89jYX/Ds62HgHwen7KmMGkY
BJNIPMPAp5CEKiPA5RH0YF3RZZNsjQ/MNNvByXkmBWrDnfxs4sjyq8FCsMV3Y46AcsGeiWkrDEd3
KXrXL68C40y3suWEpIizGRy7qsYSS+2AxY51YnLOXIGYwraYLpki0vYISLDA7mfq+eoP2zj7+CiM
EX6NNBnPLKKi4cKtmfq3Hr2G/jUGWFrTRscBB10WsvNbLloEwDlB1tQoCAQOiKi4duhmHiXvlCyg
lXatLKb7RC45ExsuZu1Oj8vtWs2pfLNSGxSHZFngWhg4I1xr2n9xvICXB+8STQF/KiIVBIbK7TcC
bC9KGuA7Ak82O4SxQGmGrlF9nV9KnEHbzTSY5ap6JkuArseEVkuGxK2bzPuT0hRu4EIH7cpZbBwI
plWDiDS/GrxeNk304o7oRiBP7GaxFnk6jcyERBCX7YAmRJE1a+vQxMZ7FUoi4c2gghu8Ov/nJ+Ws
6mLbEBeSAyeW5viL67Bj3lpatomt8uRMQnxcdehjLuWC5U9JZguxdFqPCkDkDcVpTUT314gVPxDp
DWegEHQELJoVm6KJiyAnyOL89jJuESejzIz89ARzRJuyinphP98eNMxrWZ1a7qw6j3egv1zf4OUJ
I4rybOkhTzzEdd4rlf0jwE3AcDsOCHdOjFn+jOm6hOE9xhE1DR0ZU2wahFjzAmgrYQ7xHZBTKw+y
irvuAC3gDXYN8wT9+PDADzMNB/6b4Jueqv9W92biq1zWjRv0szhj+lvXJgqchqKDvdrDofD8zk83
tPHSEZdffkgIzzQgVW+YwFAG1ZI5wEj37Rr3FwB0Neg7sTLJwR2s50yCZkPkno/LepBQ9LSm9pgO
lMp7no+XnDIGXbS+XN/hCEP/CTOiZ7PTUw1yyfVX3xNVDJZAk6Ik7GXGbEptokMNK1Hr/lg4eo19
/Sk/JLXZIELv64G++p03lbB/EyVG5kXqYPLF757KWyYnYSN5dxodhCI4CHSM+PGj8PNCLMCsjofQ
b5QEldgXqaqv+SxGQjAFJul4qw2ITBwy1JLgWYCaHpANg6LZxD8MSqA1CQf8Wa1hpmmu1+wqwM1Z
jT8Y8qF5Y5DS4j+mf5Ibqsk5Ny26V0+A31gfT7YSUxv2pDwYicWXB9MVEZhydYJuZ8omhOQ4OzDJ
3ZcqoI0Kt9FcYe0KcCPt6nC89z/gvvNc+tY+GB37nyaCz33o8h7tvuw1YVFSdMeul0VauAtiA2jA
i6B2p/UoDL5dlgxBQ9juw/iTjeb3JqqYYeuwKIUFfBwbf2w9p5/L0fwgTSq+AzVAy7cTQEl0QXHl
Nyl+gAhQIeFvR0P+p4yvum+tmrhsbQS7ZmBTZUdIwNE/5TH+L7c6totbxSlSMC5YMymvHVP/Un5Q
hZyE5PiBaF69zF31E02qDJB8xhV+llnIrG3cSoDr1VlrycZ+/tSpwCw0qlOuO5F8OgFlqV06pEbr
zucSZHqpKqmKHjFo5bFEwArXn2StUCQ0DOxXGA/bX5KVN0Pzmm04yZ1ZAb7/OXK5rGVtG03lrYrw
YiBoWDw0fcjNxm5beGJPqa7kNHNdrqXN4SrcYejdKYreHPcVOorg2FXe/vk5JU8Xbjq3uCAalX/d
b6QAkw3RRzEPxm0NBFbG+D6Ge0xVlOLZ2WiXkaj+xu9uoZwsTXFRrmEkKV35XDvFo1PYGqrZlqII
kUEfEdJg+3ij7mtss+m0rzSCRy1/vC6auiuTJArIgnswPAjkrOLqcKhtOCCBI0jCF1O3Cqw69wQC
gtPRZSSQLkgBSD5zphUeyuMMp3TOwb+JxHL0CUuScfDEFLH8dOHNEXzqmFPqhdfzTAMXjKl6dyre
k1SMfN5t/BMyPiYjkzz5RYi+jpphkK5lOos21n/N0rkDRCrK2p+9QdkpAP2VO9AXs3cGwJk7uPVE
n7JNMOwmXSwX4NjAakVvolBrO3877zHHzd4jnjdnU86oAGEWEENI43p/VDR8hGmv+31TMw6eHahl
wRa5S/PiHTXlwsXgb/e3c/9r7i+vuMQJZ+ghnI7Qt6EWMjSsiW/I18SKIj4TXEfNXXwOG3ebdS2F
7AmKXwB2fvlcklHOEjKeJXC5d2Rb3oxpV+fIt6LNySj7n3+TgtXiSPdplx62NsXLDefsdZAqqtah
Ej9H7+yCDlJbcKPHvRE4tCVAA4dd8UeWZWaiSjcQzjPm5u+8XpkB4Z5WDdMNd+W8hMu9DoDxUGB2
QFAgth8HGJVv8ny12ZTnN7x5NmVRKydrIHS3fsKltLUAcg0CA2zoZgYepAcoqoOxE20LH0/T+xpu
7XhIQJNHPsr6Q7u4BmQMVVRytxGAdi3EYALLfArQBDg3U7vhFcMHcFeMUUFIzoMxTZOcyV5Ad57H
vGPkS7g8Py37kW+jvJC8P6aGHvd6QONLUsvoedwCmd2Gy0fOSHqpDEiQES8RpFLOtZ84xu8j9F9U
voG8HgxIh9vyfQfCPoSM607G4omWaMvZFeM510lD576aDz3Y0oswhem6YWLMAELGrK5jl3OFxFu0
X08gn/kMxYE7/V18/P+tTsu6REpGWDsxzM70mEqswZD3SraiGSl/i3AqnY2+KPhxtcbABkIqAzfx
HnLMNXc+j/dA9bGcPsn91ieQkPHTKm/ISDczqPPHYZJr9UkWzUbVT7lBcRQ/wmL4Wi6SFmTOmkwy
68nctlX2Cf5VRKfm4b1aecNFOr7d6HEUkSB9x+80PVP2BBc8g+dhmcl8CoJ/xwhe74AfQMYP7OJz
aY9uWCFOSc9B9zwOyyOOMRnF9ShmL8tVVXz7iT9aT4Piiu5eNRqEcsygfSN34arX8unVSkDAfN89
zAzjR19MLeaRFg1XacfWmGY7TEgeuDf5rdZYWqk2/N8E+M6Q0kHGjj9QUe+s0h+uKgKdKZh6lBRZ
ZrpsjymYXWOaFU+wPly1tjTuiAaBLAFhFKDgkTAVfllTPyrr/6dWlzMCA/uuK5qZTGlommfHB8N0
NP5UZQikVtkzFhna1w4WoriTzqMqYczrbXFOV6INpC8Pap41n+yq1y8reOkgdfvxXZ4tYndndU2y
9o+7CCr6ewEeYvKzCBKGMd85fyFA/pLw+9VPSmxQkrA8EhBPeCHlb6mtOmMnEQsm/duuYT/JrbPM
OdzVdPfr3zArjEh3Z3imTcG3gd/Qd4gWn1y08MwOQK1ijPRvWgErLbm8VKMVA4rNlcDntEuP4f1C
HdJksbEx3yOJH9oW7b2j5JH77/Km6cwshja3ECSX5R/3PFl9U8spReVkoDNztE0FhUHOb98yYvFr
L87gjfEaqHE+NWbdsE86zaTicUU0gv4bp1HkofQlLOA88m4zpbmGtI7/B8avabQ5q42xdrgpvFv2
H0G/Y5gDEeFM2I24mjN5V0XZYmAYy5sXII6zjBnkzU31VUPBO6UabrKB5EbutLTqZlSys9muM5JS
RC+Ll+De+V++FA+3fcGmYboQkJUX/qx1S9lBXPfdrAK1MkSbKQvhmZTo4RWY+I5bKARxKPQRb8S2
BayRalC9MpSn5xzf6aLVjNYOY8LN0IvdgDivx4c4qZDLSCDNdDWln5tknfO935XWhCtJEwnqwaGb
esW89HZLmp2dWFdstGJg6oCYBIoVkbBCAODb5SP5R1qGnU15cvC3dCZmnldNmLkE5g62T6R5qP9e
XdA5JQT+UPbu/ewBzi6uh7z7FzX4203OvUblVIAzS99T1wAklgpYNgYQfalrbesFHVS7wQ25pbDn
AXaZFg9MCf5QTD+iHG6qvOQiz/dB7iX48WFwPTax/DWAq3gB3nKdubakbhyTCaLH8zHei3m7E/NX
ExYFaSiLzm1rIS/uqKhRzEI1kT9vOlDZVgt1DhmQLWOmLDj8hc/gNjWUlE0UFP3JpmTKtsqaovwT
f4WrDo62LjYXlEqCvQdlvEwwlAXrto1WGde5TBgr40sxUAH20RCKVJPTwhl4nDeMJi0ly74A3BOm
uVpb/+4zvVVOnaUTDjYswQvYchJaSvXVf2N362YiyzfsjTjXLJuIRXkfnsC6y7XxRH+uPZhMNq1z
ApuXxMqsDO3lh16r3UhxO0bLQMxfvxgrK7I6ePia2Okke0lvskmU4j0D568zP/EEliN4v+AM+Z1u
pG8cMPdsDcM7lFKaMZL4rTM6wARdD6Fpw71UNMQbmvR0SEgC56JPPlounKSXCAeEpC4p0ogFwygD
pFJI4w//46mMqeF2c1nBw/RTVzR7AuDeNEX/BH+iN5NxtvSHjXLS/nZd5RvC0I1ZLBpTPAkh8qab
EAIFlM6GGpWMwgcx8pNIKXtvlDXE+q0BZmZ5fHikxQE8ArGSbencPBx5O0pctr/FY+PPpCPqesN3
Vmjh8Na7DOYfaHaaI1Dgza4aEyUqP/c6Y/axyfaHUiU9V24O3ZvKo+g+5DgmXClXxVDIVFXx+NB0
vIUByDJhjR//co3DGb7mxIbFWEjR2MSJeBtk4Y0cx0s6JCu5BxM2DePFtFeCL5HJpaZ1O1Zft7RM
chm6X3tI7btcFz0i+7HDEVO1AP97TNvZxzQnCMczniezGyuHMt9Twi4MFxhafXsjM1YLImsBya+i
UMpctymX0rev8UOkIUOWSr1cjDpEJ2q5jZrZxo3UpE6kt9ebaAGYDkxhqaSdeykavjJOdAxvlKMU
/YNUNnEOsANMzYWyXasxBkSj+lvJTV97kjSJZa1SdJHiKA02SOgFOK8dOhrd4iXNfVEXD/a2sMNn
NS+8cXZUuE1ecEl95a9PdzKM48N3L8gSvRymmmckYvyXudQDW1+sDeQ0Tkyx4tFSrV/DPCliHysj
L2oNXch8/DPC2xYnWBZ4Tip4bmOeZ+6HbRbQHKzRKYfnDwZND+pOF/dsRjjZfpaOWwbuPnn5RsKl
Msfi+dWC9v+Cn6gwrMfgNM1g0izRaELS0a3HpVBo4n9vm4+QXZ0iJfUTv9LLYpvHhVQtwBM4vOMS
pihVENj7lVswzE4E4989VUBQ7aF+RFsXxrgBZO8qsAgJo8ckcgL8yI3C0BhDg/8tWfZD6QZEe8e6
rqAswbMwDofqhoNYcggIm1QztG34wc+M3NEJRpiseBDtLwE/Ww42w+MLL7ka8K6g2Vg0mFbjcHJi
n9eEKBK0EpEi+sganKQ6kdVuSSLFhDeAd280XIntcTyifKsAIumB2LOauWgPpjhQQRoELMaP+dc6
h5STyR+fgdUuDcFfjx45Kqj9G+WMPT1RFK28/9NkPArKAlOC4i6w3SVBymoeRu8yZLREI7Nz+3S7
PtwxO3jD0PWnm2QNOBr5T5vbdtomHPZQtpfNVkk8DKWe2wjyOo369sFCO3x+UXJuctsDpgf4KrAA
q4HYxuCn0WYtPFburMzBWFvrmizss9O/LXK9TZIQMaL/wKk5TgEFCzt8bCB0iYtINFbalH1npIy3
qlj86ABxA6iOLNng9FUYVgqgEhQ2h1yKNpWFUeReXGnFYlXDZK485EYaLaZVhl8vgplp3ftqMlYE
zCHU1EuDYAoD5u13c1h9kSrOEwEfW8yWsUG//0g3VknSYxUVy9DlxOXvsX5NXRZY5ISzTU7ovQli
JS6CX//tzb+hOUm2GxssoOOcEgkpMRbSKvrGUK8SVTVLegb05mjFKi8xm6PzyhIN0KGx6z9BgL9X
T4OazJpLUNgWE91sHDRrCYVkgfOKfr9Ql7ILu8nOWHep9vhHC2gOuQUK1IHva3pMpcMogbILrQmD
sPuuR79Ggv+cxNxBZAQoqA6MrSMB+eOJJh/5+KncpJEOUZUUaZDRKd1JsfdKr1+1FAOjkDeZEJqN
my6/JHaI/Hkhix0qStSKzEKe7iL2uXrxDBBp1pSol3a+f4nYlVKQyI5lcw46waNKpsbSgks2QN5Q
SqXweneGR0NPU98TV7wDA+FAD6+Wen0YVoS4xgAU74RCBcGcgBX4DuJ0WJoYIfzg/XyxaowgVyho
5qar8pQXYKtfPco6SfWRF+3+62cPY2p+cgcBDgSpG9jSDLjy8FwmnQcrxPnjeu21q8osy5L4H3BR
AK2UYN1zkyP9DWVc/BwHlnM03kPX+K1y8Oaz2VL+zlj4MJQozOuODblAFAY9RJhBN/FQ1gU4Wsq4
Oj2VV9XN6AQelg7ceNb8X2JMpbwhV1Tfim1wWCdSUx0eBNEGb/5pfuZyCVKXOHF69utpZDo9w/3Z
ihbFKaJCm5kfg/Gk5XNQI6bcteHzZtrboF8ECrWcIZq+aTooIAQREtnLgDLJAIXxNsM+Skuxuosc
rGj5TdEKGTDaOOlalCNs7l+lkAmu6Iz0h1bsbnKBFlzq/CtaOpdL0KOwIPfm/JXmQAltogl7jNLw
rEREtvhjlTmpCpHNiYdms6A3pFzanr/1xqr1m9qlyoc/vTVsbGHiMD2SnSLNC2Wa9xMzv+pLR4Xj
QrOFHofLJsq6XrDDSHa2EDJGYjj3ZqRZkpaDb+G88uq2bdrvsFfUaK8gTbBJZELnR17goXCK2pSQ
svo1HQJKXBT3vyJFMzRBt2k2U+1YIQ4HrYUJTImskNQMbsE+EBDq1JrCPpNNHyIBwUTB0iRLXcqW
fXUQ0OzuECifalN9n5tNPd6riTrMCwNKFqcoXoCL0cIv7z+Z4MV2uSXbfgMSDmVO/2aFE5Y3FzwM
zC/OOFk0wgj6T05HeUnrvtFzz9LHaIHVYMvXWwtP7TugQEqVD9yvKS0Ic+K0zdKgYPPqUFX2zOvR
aulFyoP3qcC6Oe1wzD4hm4OYXpFiG9uoKnJuac9Urize2SSSPGA+Xvjau/hW4FhM7jvbziE6FjI6
BXbMA/kn34v9fmF/OMGZoF23DAtEQUbJZxVH8tmJ+VezJ9lceFJFR6OXdOFaNwo7vRlZn/Ftspsc
ARwzu9H4rLV9mS+PeerB37pFRLmzmwPjvWnDNzjbPFOzaZT+PXY0gwwTfL+Vip/W3/XGRMbM91qO
Hu1nSRm8/0ZQADlxq3RTTUf6J91kTJFnwTz3r26CMc1WjuBoYp8XyuXMNJWXgc2NBSMe1wdb3M3c
VnGDLGW/ExnDj6N/Uqj4TpvauSGTiBEGVDKXKRdQ+CEYeg29lmpLoJGzj/sgPfezpDOcqaBDwdpx
XuyJI2/sreLxNq4skI5Xeg8Y72H7uc7kAq49ld+tCOLWZffx4uZ8c+W0WPYOpNF48F3mIroLIG4n
pobptt+E3WdMNcr3IMviNX/hQiLREdjXHR487VWvmY5EBiVFNud4L6ILKXOwYaE/bmhQTnZusNGX
BmCKjbSy5+FELkl9UrhdUAE5AQFAOpDlrrB1EcRLsvOx8fMUzH4McD1HjfnjBJBZOagE3inWgS6h
PofcnhnOfyQ4tw11KhfN1T0hl5bWTVr90Oif0dqW+z+butlbD8d9EEqhIrJHQKnGaFG5z+q1UzPy
0OoU/im9EF+FjC5KgkGlDkjjasU9nPx5B0OeWm9ORFyWwoN8KCJMZdyULP74NHY+Ga4foTfRrqB9
eXShVNJmcO/gXJ4EaseIKI/xpTUONWZtPPF/hfeMnJHpWjI0EpCdbmKtmXIaTzaORPsS17r1PRgY
Au1z27IIeYKGmv9XzQ0rUe9W3J0BP4RquAPKI50thA9iaGSviCfkFZoeGrPdd+QWGb/kDY5QcpUg
F/JNHt7kRgN+q/EOgzJ5ROAVvY5mkwHHVKdcNK0nMuNe97vEJoA1SHdLJihlDj6ZWCHORXN+izCS
3IJEMUXfeyUPXMMuKo27CLBuhCtfxZ7kBlGQytssXnnQxRcsAKgdEdKHcsEVNvF7zz1zZp+qAMdL
1tZrCD7S2G2mta/O62BoNu8SYEJd8HIl7fPL135vlJpVZkpyGMPxqHyM3DveDiXqZm1NMIz/Yq3u
ojRUNm297yRqIwc+3HU/pEtYEBUmicc7SbyMdQ2qbZ94F5TQyMR7/UKf7DtzPPaCSXXBqRJUybrw
3F7FqIWGILNjnFSu5AmYdupc0CU+joR6fnL/VLkr/d9DMMNtAmaRfYRkzbC6IqLrW76BD+NohDwi
55snG/a8StahAmEumSfgNyPQV9Lij9dTiq5+8+no5X4sedWTDifc7I3fras/1MjBe7lH9fU4IRRs
Z/9dNWkG54x7FdLm0S2PeL+wRnH4fBI9zNbbmHRpIo+Vzdloh22iH4pabQ4HZN4dIghi0Eb7fMyt
FRLhnN2JgISHtUvriQUtisXk6VmH9B2BhH9ivfcBD+O3o/Lnt1AoL6e1PBCmj6aqc0n2fj7zX5hB
tv/EBUMoKN6iCt0YgFmDwVDw4rJac2AH9qKOiVC1aKxWcvI2OuXkAx262OIoqS+/aHpxEU3q3Uxt
mwqr/EuV70N/O7sPcgfHQoC0dgCa5d3Z8IrdQrG+3U01q+Ldc6UUP8XB0OpW0XVABw/0b98AyCs4
Vg42DUX2+bYvIVyUDbKBmDiWaSuuNCV41sw7idERN0mKttCCmB3QNcuxPdazbT7K9lFvQakpjvT3
z2fb8ScaJkBGlhJ1W3FcOGNon3WnsP/XkvbKkaH8YYbR7UKbzOiWVJgSoiI8GDhaQQLTiI5i6Bfj
ntRx7dkVX3+HIn/a1MCY0s6ZY3CMHgp8zcfVoFNgEIhZmQlbMd7tVsBbxS0LOi+JW2UZGbMXgkIF
2RCya07xO8x6c6kTAz8CLAzSvrwI8fOKiv1Zjt0CinRcTFI6SslX1cgh962glm9xj4gwZa2HdM2R
TnIn5X+gFq/Miizjv3sIdIbwn+sW8P0h31KSDl0HAfjRLzTual8YhinwFO84qRGtAQJvFZ9Yt/sE
OUo564K3VnHxjAluv5cjwNjPUA20VgfDFa6TdHyv4MNVxZTpDldyDr5yI37fOrDL0B6UCjE05OZC
ejf5EKMRXv6cs+uKIMwC79HdQ2DPcz5DFvlOvGVcnPOTbBPOqVKTMrmAz/bRCG66kxl6m1qMgEXv
vZj5oj7tN+hKsOqHwhhfr3sbGyCbrOuJBLwZCqFhGb0SW6yqAvI2EkxN45rT16O8j8OtNpkaKHhb
whJ7s8EqcWTbq4kqUoJTRrk9jXlg97MBPuyvZFH2CrmyaRLrs/XsIj5Meg8NO6nxrfBtae+XLs7T
Y77OFXNigJkxGUMshcOb50zak2O5Pq3OmjZg0yfxqa/EbE36UFj8QTyYHMQUI/UQKBGq95BO6mDb
Nkq5Lf7hzTJwMa4t9vfcUhIFur8p7hcOEz1b4tHFMhYJYptg7+p+CxUFrUDkVteh72fs+0aB+/Oz
ChDmEEtPd2AImeyVdfPDLR51VQqG9vyjQcw8NOwSnlxX42er3dYNY0FWulINAhMEHaT6vguVtAwg
/0kksV5cHBXWS+ca1WmQb3oYnTX174XtT++Nivom9s5ECLIR3ZCEeHFgydJ1IRPMlB7v5FLRLIAW
HXYLKbDZOrCgQZFQWAmDUS4G0l8Bu7fm2jwtGhObYHWYkLRjjI3/sVUlSJVeQWPd6h1pwjrCexhQ
xlWF0EsciKkh4E2vF4ZY9qJ24L+vEW8WfSPglqsT25Qda7YuHUOP5wPaeyGKchdH1qC5TmWRDhHA
8LfTg3Il1d0r47FszAEZz6PRMm1rDhWad5+u6tDPaJFLTY9h+Li5u/2kOrbm7bYm5ssmKGrFrH1a
2h+S2cCiiQXTQw1rTy8ryybT5kWnbj1pHLEUBKtU8chXJhBDCNWhbc6+XplTyeg2WBXyBxcI5+bm
9stKdxFrxW+kBaRM5Az2J0qNOiGellLieMf4ASfmk58ImNtdGp+nzqJGX3WNPxHGUDYGhBlvuczz
CGUAvAKWBW9ufUhlcoXSBBhmgHAesgMKeZp5xcipAgoPxtS+/qeU6zVWGiR4dCVu35kZh1+rku9O
aQBCLXKpDKeAummuYkkaOTEn8e3sfp5wGtl5Iq0dfIZwrgIl3pZ/MMSbdJ5sO+wN/o3d4oJCI0WR
b9SE//BcqU0qqWOplf+UAw37X9Ri7hra7Tn3hjE2XsZhaYemB0awYAWrNWWnxA62A46JT2Sx3h6S
2/mCUi+TB5LM3jWj/qCXyn7oMciZTVW8+S61EnBHCeR3c6VVI6MYyYVySIe3Yo+3Dh0P5SRazevh
UrAAMpl/hUa6yVUQun/+O8eBf1/iQcm9JoUAegqe/sNwU24tvHZfYpBOWx24oXbwpT+7WsVtg7Wd
+q89b1lIlFd83uT7F8fARqfoOzYouRB00Oocr8WM9GYYtSN/9YF/sIa9IzykN1qo/crn7r0S6o0Y
s8H7mnZsfGh64GNIZGXShuDmLOLbi3XgJsSWr2SkTNo31vM62kdHzt54bfwE0jfXkEase4h1oQp1
98F54UHwjmC9djTLOpk80psvc1Wx6okATPAYR6ehfJkmzsrFq27yXZneNUtAUgdH/wuMU01p0jky
S8dP2Q8jmFjF5g9CYKelX6m57yvqct7YE2QUCKCemlhSPz75a3F0p19Yb5gfx9IKMWgGRAsMkurL
s2KErhqXEO4nEO7MD0Q9WDnx8/PFkNGKyx4K/9G8EbE1nuHpzJ6FOuGQ160ArmmrpKNhjWIa64gI
mdKT0c/xgfvaiXvxlorBd9z4Q8eb1SunVT2jrFWEHRlvGiYiNIH/Dn7PU5Z+TLpVKmUq392uBCIk
aL33ac/bVwGe6FljaGQHfV5jhAs+9gP7kHYMtuWHbysQyxyAf/QCwXpLlt4KTYZkfoLy9bx/YfyW
vx4FvbpVIkWef5KDJXcS97nUpQsADYSxRFrAYFO3n2oC5+aTLqSjpkUgWLhWdlnqScyiIndy84vV
5fXh8drHMTl/BH6YZ5J72Dr85ZWPI4wPj18+pMkC0nEonYFkAV0mCZQLv562HcYrzQzI6BT9nhLJ
5WvhDUi2naw+a6YuA22uuTYpf+rfKIL9Yt5jZ0W/fYw8x/pyq26U7w8zENvuN/Vg9XCKvmdk6P8E
RGgCUs3V8t+8KjQ9nm0HC9o/Uc0T+dQWJBaMNRCsEM1xkVgdFQ/SZ2s+jd8Ez4B06CDFhh14LfE7
7FJ7+osllq4+MOjCDYTBb6QETK8+PyF/jcPmtRjQouv14BfjdNvnYIA4PKonZQKDbBx/IzOtmegf
hHC4MaCoxmer/sng9ObEX3boA7m2Bgv2U2yNaNBOwI5wx3NvbLr0aoXaPqXnl7/bDVgC+ereYj8n
430hnAB5Ydk7LUVUvISKP70dyxYC2XKG2nCcsOLT09Tt67ve8B4sfOK3LVYV4tLvw2YO4HIgls5U
8x8CD8bXnZhoum9c7WHv35nLgyoEmjkYs9fWwdjIuawWtUgcUXliwxhKbT10mwmEHjLWGUrttkKM
+qN51NFaSJ5gnAgYyG5VsSpjsOwH7Pc3FgDVrvqtJgN9RipRqIlh6YA1pp/Y62Mm9+SL4sLkTAiS
/fDlSHJq3G+Pk0DnpCze64kl+uYRLtPtlIvs+uPLdyriAbh+XLTBfQ329908iIg/Lh/Z3KWej4da
PJxsunr4+Ql9l2AObdOXMaSr7NjLEjcmaQauaZrw1y5EFW5ELua5p+0xg17aQW0mhsWnaVIZaOBT
owylKJwtMJsIXr3M9BXmXVB8V+i83zliFC1/w+otZOyTM6MGEdm7sZFsME5fotmXXqBOrY2jG2UU
zZRX5QTvOD9wHJelutNBvTN6hRv+pPCoQtV0i5lgujuykQs8HShLjsXkw2yFcwoR10BaHzkcarmY
iAWH3PLrPa4OiSQF6fsPKDH0fOHGUvSKzokOFWh3ShyvnOZQlynT5cpTd6tddIU8pgFPLd3x135f
ZXVD38/Q5JMEPDtb6U3KD1g17f6hHuC/dk2P5n/nApsrTTgGktV8ZYBl2R2AeY+i00iBYN+RHP9L
zXbUHcIMl0ZwT78v6/O3vpxnkL5hhKSagZCUoP5by7u9PuNZcEoGzqxv/x31QUjRsoAMsyhrSMis
R6OQVXVPMmR0mMFX0MM4X7Bx+G4XODVqugmQOWHxEwhJHqq5mYBuFXzhRIssvaR9X2w8MOGERqCe
YiGd1pyiI4Dtwgwk40baFC3c87Pi4d38vCLwoYqKmk/FW1Z98eb0Q9vpmjjMUxGIeI3NGHtTNJ5K
lWDB8LjjlVY3YU0dn45afKkMtLt7kunvaUx05pqA7V/0vhHOcTf2e9yxfeXTUnKf6vjQBUDI57Zs
dCjkmLXe1dwdJLoZKswbWp229bBIOl29na65shrcCmd7dgjzIH9UO43L/0OCdAe/qpHN4LVWV4L9
oBDTW2zecipAw5URV6Dny/n+LjT2+VG67mbjlbyDAnNgjp0ndUwXGmrpwPyP53nbCwhLT4JCxtQr
If9hXSYJe+gZr6A06YLcGJBYRxtkh4emFba0PJHxjdTKmUu2Sa4kuQEqPvSdGRsSC0gMwp/SWzuy
UjuItrQrgL9flUjnuDd53/mnfQyzsGYHMhiyuEXwiapcoV2JxU6YpSbBa48k6h7oeZuSq1Spo3xn
XPAhem23kzq9QiU+DfxbRXQRcpKswK2+ZWYF7t/+TtWEk0WXmkbwQc2DAfJK7Xve+rWl9zhlF+3s
BI3L2KsutmKA+8FnqSmxmBd3etltIsrNnDdLZ90Loteb6ePUlukFedzhQjMeZsUhg3pdxkzbmZy/
iErhTppvbZT0BDjcmbiNr7C0jhuVSnJvSyGrPI+FkJPy7jSRe43/4/E58ZkLsOM3CSI27UW1RQdQ
9ri23yiJLVV0097Ivbe16rm1sf7hLQCQtO0RjxA3LfQ7F8KvrSCrM26Xldhrb5iZqf8t6Jyt8GRC
kfTiI/lTw1Jr+ICUqjf+6ObdTEyLMYF2AreIrsz35lGaiappfLJ14NMbRhC56McLdV6PKwdL2Crc
p4indvItpj7J9uAel607+3bhfzIdcC4sm9hLtCSHNlUqOIRhnJKag4gNlJBlRFyxiTqgrHU442ta
ibMJMNboxVn/p+oiNtYzJJVghNLiu9eFyMPzIgrqxkCWfTieYMxQNN7tGN+TlVuVKAQJH5WHe4rP
a5DkXxlO14EE+DMNcu9oY6R8JXs25hmyopuOHKnjAcKxwzB2rbtCMGMVUOaw4cklCb8x7Hylk4bj
+o9i/01ou59s+Ju8EmqriBQU70yJPIGb3QJHbjqBGYuroiuTrnaouQ0+yrQHgf9mnWl1lOqj82Yl
wHuCNBeYPzaPX/8ajI9ovOgrN1H64LbyJ/uwwn14kAC9XSurSWmxyD3awnQmPTwEIXBzm9am8GJZ
plkcBluEK8KhMRxaJ7m6HPOhp3jPuKl1gqXQXzmEhNs5Y0BmeSw8uqTrYIJ8nHdFx0q7TL/kVpHz
6PDwIhjnMEZmJsH15eAgqsiH3Zcd8mgXQeyRg33lHvYK6nKs9KMPKHHnwHEtIsRVOD1n2mU8N22q
n16BJRTenQf698b0PE5VMJ1HK9ZGqfGxzxvRqmwLwNCCnGqjuOL4c5EM5lnnL5xMZFoXUp05CcVb
56dXGBA11ev3VhtPS5lFn4319GO2IA+2c8KNCJyA0T5xxo+0YBxXSnzfRlc9hS6DOdXtGQDp1z5A
QvM9RjooWeFVnDY8I2S1HshWvKjgsCBzA81XvZXZn9PZ0vIiL8L6SNBHzAybpP7KTDbwP9dH4ClY
XsOEzQp2PIDyQV8cap7o3LEu/5pHvzPorps2dCRIstvuKx/heSAPJfwktGKhV178jmuqnMcnOMOD
XDAOmaGX9ZMZbcFgNeUzlcuXWKbPlIf1VSNefr9KnHVLTfS1ULOd4MUuzgO80dJrKUVGbbIpo+Id
EffjP92sG0w+zAcQ0VOdjgCfD9azDPraDKbzPybXeP+fd/SVWxzI6Rrsk+bemn07tEkWPFy0lTp4
HLUC2gwNSsC7v5a+sKPMNJOArkn0mL2w/x4GL0B1M33Vf6FjWqPXmirAfs3APuFupPDa/3UwBVJO
WXSTx4pm9a0yuNS75VzPb26ouz107+cXazLyrjjXrwaYfTaek24m8q+Lo0ulvJz/AJnqM5WV/nqq
1mIjRaUfhewSokYU6tq+7zkAXhOZpryJ/4xgbWtisAwZEW39X7PtxLbdEVptly/UBgb21DVVto7O
cDyYdR7haJZTbLg9ZsisbBX2VkAWoKKpQVnQAG3E5nQtM7dAitLOQyPpCa4ef+fyrKiCkBrWbKQh
HdOOt8zNgudAii/1r5QPXu/ashabKT8HxU8s/o5N/dQOasfSHJAlNrwn5+CIqwAdzM3PUHLvFn2J
j3W9VaPiO5BVKsJ2SxS/FnJDBbo2C469l46BlK1XVh221tlsVaKwfdTBRj+crqjwsdbIQT0t2Xm0
z3BpWMN7q+kM3INfdA1sS/L3S7TkTbSg63KnSxoSvCD6nr7TYPZWH4YMIXm8htaaoEWtvr51XKgJ
jpabV/aiungZtN0pprU4T16rrVoS0byXwNbENIs4JfLe/LwM2on7z6Z7rKuuAVwmXdzps7R70xMW
U/WkNqaHlsLjWqj7kTnAvOO4qg19uCi19xwAAiU3oFRErjrc+4MXn2rtiCweI1yTdozEuYNUPvzc
fNTXb+qF3TXgfDqd1A1M/ClKUplh3WlfFWL57z+tYFEGp9yD6gZSblYB6y4QoiWjF7Y9t1FIT9Lb
ESNPvxPWNGl3AVOxIit4qLRW/cMe3r34zi2FbM1OwRd69//UqkkJ3ODz8rA42CXIuivon3PybgzT
fpTIEPXs8OvWCsPKlcWTzXx+UIntVNtxf+WGS5/FPh4UltCgixdOTNe2rX8CWL3xNvnUKkfShCJ7
l5QcNtUolYoWENq5P8ZMpfBhzlpwWvjrybpQS+3uo4Zsed00IR6D8oi+lK1fJ26TIsY9E2CTdfEI
ph3TSFWrY2gZIH13J48SFcoXaNqdLSndS4UtEe+R2BfqyGvcyaSjKCveTmH9cnE3teOWQim8Q/B5
vy2TJbyT1pEt/TL9SCfhJ3vM/awqksDLudIUlmjN4aYdIyySJBxLLl1VhyiBImjTKeZK8upQlSXK
46CtYmG0hfcYBdovSQcxUIDP4A5AbLitjRUfa7DpRjKyaknGYHW2y4RfN/9y9/qQ5LBcx0+WuteT
j2BSDTJav7xJrpIzVDDZlGWb9T6ro5NM5lychGHg9fWLiwBLEUQDfoK5J+VVNniArTA6gWHhypkp
EyhKJfKG9PZik7vJRQqG0jFuSoFWEANFNAiXd8pMOGWQzdMu4TPBAFH0W5sSA+KcWlf7NHvGcHEg
FgVhRZxlOMQbTGS57fmainU/iBYcWdf5rw+e+WhUeSQ6vj4VPKP1tf7niBph5/KrfUuXvC0JSu3x
8qunvrzAzsPE4hUWtVsN60Uu09Xsw/U2PIDxDO3mtE+bDzKyH0OeWWfOotyUuqnjyEI5DKqg2AwL
X6xHWKTqYKI9vb7GJ0VRN42EOMMVxg1wjqCsJ6UPP5+Tbn5FM2vhZ0w3pUe7WcvuY+kwmSXf9ifU
rmqPZuTS6H9S7w0dAXxKRuYLddeXOapmO1G9xV5e+UjalhPQ+UNhd+iM2fkEuSFHiiIU9ysdXYSf
uclzhYmO0k57xQsxicQ+TVGwvATH88YVVNIrebn8sXC29kjVhhu0Icy6rTppEWbfLrEO1+vnbpfG
GWsygXQj82/IfbqMa2Q5VND4tuBPZXwacmjxPjifkumW5pNhJTF9TMhTsj7lGstpvZSTwxTGnWtV
TTDsEMLWR1zwRVUTDa1kZJO1h3kxlsdt1mOWAfOQNvZlxZNiNE312FxY2QDInw+fP8/A+dC9KB5Y
bgSVDYiMK1wz1DFIjwc6Snt+arejbaSvGbIdwjXsmfGP0JMRQWzV4Q7CJabNVnq+PRuJK/Bq033J
e5hsTIrODvwfJ13xVcb8SEkQnccJ7z6X53nC84A6Ou3kt/7uS9Wb3Qi5wBQia29nCQCqINW3BxPh
cIKUcRXzClV2+unZSpZt4Sy1BH4+dV56+RUdW5eOFKNzGyxOLoVaAV0WUmM0d75lJWSHBPV0bqcR
NcY+MlyiTIXc4CgFsuMeCA0Obd3FoJnlYqC2ZqhXRc8DiK3BPUHd6reZN/lQ3FPaR6K3pQgoX+n+
S9fPkMdYmpjuRSTqnRma9vbKs8bq1O9op1yPd75YMyaskGIWqEWojJNwGRRugoUCADenP9ofYy/o
Dp4ICUsKiYSrIAuSvcS+8KbKbmQuptj5N5PEX+1HaDXry/VAnmdVNnBMFQCudLfd1kORiKEoScqE
KdHIBBIev1RyymN9b4rNGeq92xUcMhcKR0sJ3GUtmK3Vg8m/OMVxWI7k2Gs0Qvryke4cJSuTxAYg
6ZffsMomDxovnnX3Jmug02BE7YN/Mr2DaDey2EnJLelAsxJ/i6w+o/z7PIYD6IiuVjPCOJi9B8s/
tMjmxQ9LsoP6jVH3qB8i1wCFyZ24QkUu+x+861yn4w/Ne30FDBXxBtw19Tg4+Y9Bz92wMn5bqQAs
nYhsLVD2GV3uOcV6/PYVRTH0yu6D2pIWO1+niDQJH5uFYGkDJksXriRtV2bq1XuG1rUGpoDn2AGt
MMYJMYyX820cJYS4MmZ0QGwSuEiUB0qCsRqziIEiaBOqaovbxE3ouFpWpAftDL19f1iBdyDavdVg
/FBtKuVvwDdvd3dAejLD9/UqWCy3lORbgndAso4vvplz3Vs/e2XTaBXHtrLQPVBR3z9fpEYRkG+J
l16bhi8U8n/ga88MJz0CnMIdWqEMEUTVYxxAty+f7fJi1mJP1TqD3GtpmHqrNFYNBPEyAqHLhGa6
plcSFyIyhQmxc97dHFhDvfaf3aVIeobvTa5CNUothXHqV+h16XAM2hD2LPHUM6AcF89Bzm6HXvtZ
UZsDlx9x/3cXciqnWd+g4GlHGpJc/wb4rYxo6bxFDB4cmueB/XrQQAIGvLznwvO8d2jBtPiba7n5
+PqOM1t4Kptn89ih/6CbY921YhT1yliSvHDydVJBlzANiRW/Je7qd+q1woCTrq/u7SGIZRTmWKmD
vUhrAO5adp/+goIFxC2GgD5H7SfpO++lEi60dv057R3rGhlvwpJY7wx5mL8JEVjGabtLVvcthHYq
RsEgHxq+0IpI03CdubNO33JVkPiBZ3Fh7ApMY3J2WJY4CFRC5ZJWTIgCvLq6ZSfRYUJQAJAFeq0/
z9UThXeNz7YrBifdI735FehCHoXuDDiRlWk2t3WY2nO8/VEngrYUIG6OZsvetzmiynyI8J9XHleE
eBZFxpxa2Urbwi4r4+ebU5Zog1GLo26L2nO1ozSdxZuloTqLNCB36KWLZKhq0ltPyu1CO9ZdTgzG
oOqsNywB+d4FrfTgP9j8I1du7nPNYQdMBZgoEsrGS/Tk0dH3/CrldzS+4m4z7UiTCeuphequSMTS
YeSyTa2rQR0ZRGvXmn71eFL6eWzn578LrqucUWYHznVBckuwN443evUA72qUc9bIq3Q0oHQJOGEi
SHapPA6yJLfmdZabyoOYdqJSotYKu0VjeIcmVYgr5nPxve6IzC0YzSQYWB8e5206aUoEieQ5Xacm
hqV8sNvCDywXYZkesjw+b7/ojOkswrz1i+TyP+WJ2IckNo7BB5QH2W9PTup1BUe9WMLEmf1O0xR0
dbGF2MrGKp8iuMjQxBQNQgDwRmFgs6PYSk/NbaGkjC2voFg6/EXnOmtCIZStC0U0whKRyHaLF6c/
ac+bmB6JPrgSFB0WGOGHPbBpVXqCAm3cyuVltYNq3ok6mAzzONnIHmEUw+Eh02RdjgD/wjH7lYw/
FY7qDGh8GfkBcJvjpo69Rhj48PoPAfU3eRWFiNhTVWbpzwgOw/gJvQaG+izCu2vbi7h5kYTBiEcs
CXFSYGt25anc5UWslMfg60+FXsifhCPgDShfwZqmEPf8QR/8kQtSJeYxZtk3NWO4A6ciJMFkMgEd
vuBcF9MYZuFNJR94Z4A2tzcTjDSY5Ae6cI0n7XxdEkT3Fjv3nJjGgnxLK+HmEaGUU+cnr0keIz/d
AOCA508qNUgjmzNoe3whjrh2LLRA8x8/e4NtvySl7Y4eZ9Spz0qmXEqYeqFaAr2af/OW0dYBFxL1
01FoXklwKsRv741l9AC7HYbuh6jmSplIaU50isfdIqhs6v56LhK1uxLiFbCs6hBkPk6GiXYFQqNg
zrbonONTalXb4WwLTFh3h3Tx5R31tf/OzScOEI5fq9YI7kWSPWOMN/HUsizawI5FatRSpWHNG73x
0bzBpGTAykQsb0Zpqis+ouWppC45wjfR+j9mWegEWRM5TqwvsdQov7uSm61TUoSuvXLQ37qXrmhC
ICzcrRfCiTNoC3FpgQ6DHpJbkHWvpan/hD3oPOZ0Ijwk30hm1ppc64z+6xxbSYG6C2grLACFbB1z
1SCA2PuZAivSJzgXIAyLUZFk+RHEcnLMWegZMy+oC1hixf3vFcdcArOi2LJgUJyXva8aoJ4MPq/Y
mB3L5s4T3JJ+5VI7ZumYgS7S/CSAl7AH65wDRICF70Bf4ikIyVrbouaAL8KJlfJm4qGK+urUm7hy
Bptx1KVOFjTFKqueAXEBohpy0FAPHArJ2WnD5LJHIKv0iUiUjVmKOjmhzTWXUG9hbCcw+MeqLb0R
D5OATh58bv0v5CA9Wj213DjucuO8JmhF1jqcptCqK9eH1wWNd23A2jQCenZ/0oH0bg13jTuvkq8J
LQ9jxNhi2Bg8KJeIiyZ9ifp5Kojs5//Iv7FMtZEsTmvzjgBtgRkNqsiA67/lmxvSCp+BTeuVgKop
unJA/7/qPL9zBaj6+zryeOhxd8JyAaTr2ZVuIDsTynGK6dW3J9eq4XHurgITU2cQUkE1Us0/kALc
LrLF5UzxnAZfayUWajdjNiFc86l5Q/BHL10yylCl9P6BgijFByPOhR6Z0XzttBMKy4yfbcMY5v7h
nwAnqAZZmFttf/zyDwF2+7eWqt7aMI0I1AphIBvVQx8jbsVAlY6Ta0+BLrLGEUDfCw4E2B2aG2nb
yi1pIqsxpzqegTCK+ES1VrnehpsI6XlPHB2rxPHewCKwnOY+HyRTJWGBWZfCAKwRadIo+Rlnk8UW
n165Nt2/jDz2QKE6mc7DKSlYGYxM2FtHLQWjQ/veATJfeGBxQNma1H6y9/caYl+iws5HiR+4sUMK
zFWRpapruSLwHzTXjXEAjC7ldf6ZINxylKB+tzDi/yW/y1ueIzveKDPOFbkDJj0vtGzI/xITVAXF
s5cxEmKq3Kfvx6O9NnDWmo0DVnFyFRzfBIgCzO1vCf9xmmK+mo1aHV35QKX28/cXEoVGycGHd8VV
LJCOsKhXtpxH6Ynkbae/NfKyzY12CedOCr5ihY7zv2wCnAMNO6qNtk0VaqupXQ+o6KxcQ7lyTVCD
sKL7lui5WbzSkFePd3m5O+4nOKJOVGYENW+g4+QEuXTvUGgHnGkkY2I3xLeH9DUaPpwHZrLPnQ/w
iY3u7J0A6zOZDWOVePnXztcXs86U/0fnUaV8Ng+qV6jHlYpDRrsoZtkUouPc/tWASnsaV2YSiV/B
4eSSvMgflltMhbj6M+U7+79pkMr74M3oAsEzF60gxp1lwXwJVQ3Glu5TRDp3SJZx/lm6NR6JJ8ME
q1gDHv1LYgHpVUyi443tqlW7J8wS9P6E2fNwy4xy9jFUNoE2njvORbkPDnxeif2EnzkvZu9NA3Jn
1dFMwRoHghmUobcI3zqB9WBCx4nklE7UJHwWlnj3/qX3Q/f9UaENUDMR+jQm3YSCR39kq2Sb4Quf
yn6tcM+i9dtz2Omks1+dFenSOXTWOVp526lGUajXHmfbiCFJhQJWjoMPVemvOcGXzDCP9cHcSQXQ
VMJ2bHnE4CTCExA2ZUsAPD/qKogTKVncPpxPQHQ0yBUwFHl9JgoEvA1lSWYtuupyTU/kEwlYrdh8
N6rzLi+N80iSB4ieFw6dwUxotWxQbe/XtF8yzNmc1wi39sue8/5LhcNo8IfdP//PaUYi2Y2Gs3Kg
Ku6GBVWO20/YeaM2F8Lqg2IOa6aE4sTtsY3OR6Zgq6+b3Nclgb/vgeyXbjAXIjhY2/HLkDQN5Uo+
/DRbxzzLOkp1drmxeKV+64Q0bKyfA/XxRQpJ7eVHWg8+8lp3yZYVrCz2BerNDPdX3d6/t3iCRI5j
lO+/L2ljc8JgzzfC8S+KLmmSiah2RL/JOXxj17wq9FROqqDDKQxODTBHTWWZR++OZkAi3rdBkqwj
na3noU+y/E/iVGyheoOQMAKn4zRbin4M26B/6pJOYcTyfE820G3Njc3cMuuVjEx4q/j54wfQ2yt5
MfaL0M+rFweQYNdSFSDmRsmXpRobB7iE0v+0lK2KfoG9TbKcUx0WJF5aq8A969677pH0gxi/JKPZ
0QI/5Qcl88JdjUFYQy8dCvkhH54pZXHvV6AU6fHfAy41tkE83pZDr3jz1xV4klHxqvJLwekDJQwp
rz5vZOqV6c9X87sjnCXpSdDV9xHkSvbAx+R0HlYahkG4YBxt+k1vdT9EUlyM2xXaQZGOOqdvSXQj
4k1P/tVZmeVULPyUU/Xj/hO8QAOyR1iWi9gHy7VyPss4Y2X5vQWHwceXGSQLtfzLUh8AQREAvnXE
V2qhPT6FBjix5aPv3oDyP0MyTt8xTMeoI2qoXLqTbY8FIIt363JsdqOHGK0PwEfooQ5cvvQcciGP
iy5NRtd/+UIIQLdPDdNef3SbuW5fn/Cwj7OHK0zJOx8fkEtWj04Q1BRxBUpmMh1zRRvcZmJeqyZI
mmIsk8V7oeUqMrH+CGZMllm7B9qHuSgx+POQgiqGeJSvWafbfWGpJ509+pLkOxRnQ/h6z2QvbzBn
Cjfko658k6AAGL9JS8oOdLhQM41Zh6mOHzcg9u/2chdZMve+/PK/9zpbovx+0mlvXg/lsHLJdU8r
0d68wpFNqxhSIA9W4Jsm3S7HlT5gtjnYpajLPpN0f8Z5ROej0jd9wSOpV/hDu+UU7csijhKI3MGe
ZFZUawVxozJLoThRETTFPMLCqVGwG2t9yI59X2Lf+SpOEEpyp0jY4zvVgqMMWy5onVxkFr2RGNWf
LIsCVNUZGG/zC9G3+M+ZtaGZJVJxSsNhCI58Pqft3rGn/MQlLXoE/qJHLT5OcNEgeuPQr2dlrgEl
ziHnY9rUDXlkFsS4O19clhuJZe5seQY3Y/XvAxl+ogo+AunqRRfmM6vW08MQ4YfR04KCxa2gEow2
o8miijJuEXZppmgzbURPJccXyeE9kDQMW6QV5KsJuRhe8/ptLeKRXij8Pkw+OAUdyjFJS7XbW2fp
yf/EdQYeywRoCwYU6xjD+5Zu6e980fBnkbGnp9T1PdwpwnFqGsuyvvKJVqshSFTTeug4IbJYpERL
6HfroAuupAe0lwqylmegGcpk+RjjJmFwCf49DwrHdvPM8E6yFz4AEkm7OlVNZHoV0/xv0hlWAbid
whkW07bYjQpyroV+TaIhjw8fpGF00AX906jeRPS1I7o2NdmBvohUmv6O0T4d2ELB0SbgAS1G+nW0
ywlFxmxLGG/JhrrtjFJ1Vgw5UqaIrCoS0Fx3WsvAZO/mvePFrWCyHfIyO/9GktPpcUK6dYXeobtS
Tsq4mmwh4cXl0X3HfzshMwaXmu6EM3M/arkViC/quP0dJuIUy2+E6MX6zWc6s9tDNSvIDuA9BsEg
oFSLXGiz/kzTUkEXxIQBygi15KmgHZkscaSAYMZ5YVPPnO5Bk9Hm8CPyWTc2wGtSKyShtV0BxDOS
DHkKo1ejvD9b1Asl3rvLTKc5NMKoBDnJg4y/Bc02HV6TYLsq04ea/t1zhecOrSp815qjGaKWIG+H
1xCQqG3n9e52j50d69H1IthN4CwdmTAH1bg0SRH2T+EU51vVe5WnPPOvRSSiLL/s6pSKTLFVESIu
41LtuKS4DOJ4Oda93krI5DOFh7krxrFoA1/Emv96TlFxg1macDynd3IJdXvPgsn1vRCoA2bVg/Cr
0Pph0RHH3j8cDBw1wQXnnaNROxUTYsHRokTb6i53d5YFMt0lEfbVEaKij+kDNLd6XXoZTd1EdFie
77odbM0n3ns7nS/oYJ21/oNIjhY1zKFuTleZ3IjjJuD41x0tcxGU8sC7v+k9W2MylcCrUDCwq4A0
/6SrCno4h5r6YPTSFAuyurNdklpSayj1CXRGz1AdrT1eO1tsduJYnMIqnAFmYtkvSE0+pvk9ELte
YF2M+XIDmdA1mN4ud7PHsZcNDeSrmvP0Jdvb2BTRpeagQVT5XZhZU4ok8ZoxWi7tYEEIK5VxG4OP
zM5w+kgJ9DLStfStKcLtGo1Ec6IQpguntFlau1OZiHMk0n3Ml9ArdcszXTzHpvyrR6ckYMxuLJqv
vmHVNenhPv96vXWOroVBP4obSRQISeLaSbB8kMet7NOvdE8RPP2IGVL+h5LjJy1t8Ha78TJBvicl
jDbDfayVrph6Fn8b4mMP13UYC6NKyXEVzRZN5vTdWZCTJlDCZ9nKY+cl426kWd0nJHhXI7GYIVqw
0KBRPJQGuaSToFkEAgmqYNAsdy8j1WiKf4LU+phJBDKbByum5PtNlHKTGdZJPuQtaqC5xFvdqzy8
2r7pUwoJAGHqB5H0UUSugrzB+S5uTFB1AwU3D3JBmWof7R9lZhg8ROm9pihpHR1wuUz48hN8pLdz
rbR4POV3oucwBOZ8cUYbB7Anlkwavq2Es5NUyyiFsvhMxlk6gmb/bUscVXcdk6mVhUW5nrj4Onv7
cQcGH3vNzgfrhys0QzTB2ox3rDzKyiojIBmY5sbU5E6KBLJWNc+hA1XUZolFK51GrmdREbfsBcWy
T/jrAkFxvo5CjL/6Poafhcjve/iohGZeMfGZEyaEmlQdEiaAYMIKsm0dRKj9FRR3QuE6rbHCfX7g
McLX7juZOPPJtElwbBVObq+OxnvemSBMbjWOdXLnXv0t3+cb4KCH+UDqMCxs2NX77a3zdmYlpZBR
B7q6syDRcT1ZctZ1c6c8aC1y9CbVvyJZVGXUKcLYEScDqbecXjlUn9chK3ylNn7oFdR0Hc3TV4iL
xAm9Y9iNhnloWHFFWLTpFO9MKSgh0gAh77Y4V0Oa9zosb5TNSkRv2YBWDYm2eSF6r2Zl8uQ5TIz0
087NQmw77Jm2gi0KigipCrAQBzVs37VTBDyjRxGHKdbz1fjhVyxG7dbr05Dm+H9Yqgiyu9WbdyaE
LA+fqs+jc9bywkg+Z6vFVUy62SkPATvcyKafZbf3xq28QwnsKSG+zd3WrcO4xTmCZtwjQa2kwbVa
0IDtbAQE/mPIQrpotb/oc+1NzD7HQadVsgD5qO9D7ILoE5sEqT+h9eTzI+e9Mj2DqQmiLmfBZDlE
wfIKvKwAxFddvdNfn1hbVfx6TE6tanBNBPMY2u1iCmbpSw9YzotM9nAjfhQU5WJmkvJwTOF6pUUL
z4Nzvyk2dPqe3Ookf6PUb4RcU9YxBOnB7PGIB/i0Pmt/nd/YOWhqybODIcu2bZSKmhYGZSA3MQKT
jLGS9E64/nFmbMAe89Q6gf8ELtJ+lRd+NbOh1+Z7aJDV39TNkXkWCNCZaXy+m8EK4Qp4YUg0UN9f
G5Te+d167ykIfQDJl+fY4fe7zPNto+RamP+ieaY0oEOkTzbw+gKvPg3EN27MB7iO28V8iAqzOUa8
8A6QBnba/ctvWSXhBTyjzqieXCSQp4qCqZVHS/DPbe5b0eKu0dKWR/35J5JlTdDNMVF1pn2hqvo2
9/5Pm2xsS0G1QQplsoO//UCO11wuHYZqgyjRkZTIeqdPFBlTOXzFToYg2Fcmn4+f2a+nfiMKRzI+
cs72XLwebWehxTP0LSEi+UsX6BYYV1IpeY0J4cyNNG67Tb8lCgLDFWi3hnAYDUa5VR8d58+NnBVR
XMs+QEMjo5FYkJ5FLSHYi6WRB8InoINp9ZCy/yIarO0JYXsEWLT6eN+776Tww9y3K0XA+OPYTVr0
nVbZSzp4FqIsRmpHuhb6FnuthddyZvGEcnpE3lR782/xaKjDdb11rCVq6jN3lxdHrY6pL0VaZByV
MYk9qLDqgAnFPqxEkRhUCpEa7+FiEpX4tlG21oayaKLIPXD+NWBQj4o1oHHeYK3789gaKRHFCpqA
CZAqIugH7cPAbqiXsmDEjyty2MXSbqxLxKp84lMqRblNJsBb2Hw8Oz+9y6kK3y967wqEhwQo4pu/
895GXjWsyg38B8RrIYLf+1yU7c4Tgdo+bgr4Hzfn8cV8+yOc1vkYtOVSZjm7cjUu54y53qAZPCKY
WErMRVigONkO9+0H8gjWzreVaEHJ596kRBguzV9b7UJ2ReFMVH4AlZDxuzV5TbzPqWt0SgsbWO+b
l/H3SwO5dgfZlpXVMa08Dnhc+aiaQv5+phXQEClRkAM+yKcIlzrD+ocA7RctKMd1Um6mAYMC6se0
irUDLSWTaMz0cQg/7TN99VGcyvo1I56ryzeSgOguf3zxcznZcvMr2R5GdD/Qj2RTiF00lkh5z89c
yKvoHzXu/kCdM2IwvMdl9pvYu57q8TXHdRE5lqQdy3oC/3wTOpxtGwVzCEgVffukFLLyaM/3Yal+
8jdW7FuQZZlc5Ecs4J3MWoCMu5jZlh94PFpjuoaCLwhPVLbun5VqOeO8K+KqXtsKY++RWPK1/3VK
maJWrJ4NjV7X5k0nM/82ZejCCUPdIVFx/g5HQNzBPG6vZU6knI+qL1jQOPkDEBm0fN12bNltWopS
C9sOPRoNzLEcbI2qGva+j1NWfXYm71iNdoalvIssOKV4zkpWJGYqs9pJCrMzkoueJ0drWyyDOfyH
8AZ4bgFk+VN4pBj3lqgp/ThIlGmR4xUQ5i722Ww53aVbZCKwi9TbhMHeDcaOYRc250dKHB8O96Gq
YWIYsUbgV9AOvJ40TFmvtAVpisouY/UX5HOjT3PCYgrfFrhAT5WihEeYXTN556ImMwPtSsREM8mX
VqXItigMJSLnyi9tlViLu0HD9DyqYQrhz6URY/vhoGAefs0AbOS9N1EZVprccVRzk9x96rAClqmv
zZ7uew2tD2o2PwlHXaa8ep6VhZioJ16r8De7AEAc9zJ2XgBSyQyh8fNGPsNwqFD9uD+LqZ06UJp5
+G/BV/NG/EByixxp6VBZ9t6jfn/PjCsyUbML02nmJinma76JiuDQsSR86Ez8C72iDRzGIc5e5QXc
AQMVm5CCd8CaaGzMB2hrmYoqy1fU73L02Piw7vac4aVNlZ2yAtuoVUZ754BwJWFebAkJ76SS16wE
89H8J4bE5X2vy4OMkaBgqcXpLAWXOlBa2km4+XXIyQFeKwO76WzYdlIA3/alzynPDTrhmFfhERTT
9fPytkM0w6J1BvsQRKvBAtSW6RfUpxbyY4aDRPEDm1q1EaslXCLTyqUcZEWwzCsOQeFSs540DqHd
vxMqGzqkwII5mZ+jGmb5Rkpmr3kjbSbAemnu4X8j2SGxBZABHhFW0T6iVGi0uSLIS8DcheNrcZaG
ooiwxD0bvdzfIAk0g41ASiCSFpO/kfogSuo69eGQNnzT3S4eXUrIznIhFjkMszI2uwTFNWaFRaMA
w9vw8XF/GpxoyvJlqk/PC1Pr7HWqEW5YZUXACLGhuro94CuQW4DQG5NhizRzAOvrwYuTBXvFwSQ5
FBaut4k5BLc+2tlQxBvs3ypuU7qxZ86TIscT070ybFYEmTXkzLuQZwpiOr+t4OlaMIfehpZLAuCc
m1YSnIEVRWx1DlQYdUuHO77Y8t8G05enY98PLejKsxuygRBgArgbAX0xc1ujD/EGPygSL06hSOVW
mCtMPCYsG5Sjpr8Q3kQX53IV0om2/WMVchr4bt46ADo+fJ9fQSO1zW2LfY6sG2TWZrTXuf5iYKm3
AK2CKRNaEV8xeK5BLmfIRjV/mw5RkYN5Enz21BZNVjXLRWWKMrXR1zpguDi+Cx7bpEHUiT8Nwq3N
ZuVxNGS7nEtz5AzhTMvhLtHaxYQphqETWIcqK/uLox8uNGy7wVftge3HoX1+STkz4tr4Sno2JhaF
hqPbtkrSxI3p4KyocotFADF4n/cTYrVdhjsPhKoDXU+AYDF0MyMFYEWSRyo+4naoGNEwyj1dSiQD
dj9CMBExWDrZBTAASa60n53NCfNrxinsQfSL4NcOSddz0WuRuvQxg/bIkvoN0C1NNgkt+kticIlq
o16HplFLNFiaPne4D4eQ0DEFSQTaPuuxBOh68XL6ofQYSm2YHWOS8QqntnnIv21K7Mjzu36nQgwE
l05qJ/j/tLLGOyWFLSOGp7fWnPk0Fn/xOMJCI50Ekmd4DJmL3e7MaLycAjGZfjAmqBi2v4e0utAz
5MzcjQuPTbMhdhrrVHZFuC59LnZlb8KY5+YQ0HCdpRkK/3s+w/J1iO69OMPwJJ2/ohrcUpvbIKaX
n3DW3ft81LjCOtaLXlQ+wxMW9YBQPxiTcTegic8A2BRvMXwxvq6oi0OA+uAEoWMu/1vtyRqy4ct+
EK9ST24R68hj41gKfMB7B8cBkoRx+ybapZD4Fmq1JzmFT9KTdl87WZ6RE777g5Vrw22fyJDjdpJp
ExSIP5nRqnxipbuG4HONsY8EfXKWpJB8uTWUobbwRr1hNeBodeJrVVEJ0X2KLOHg45ihbdpqkgjs
lr99pjWQUw2jJ13FNUTYzwxh/6n472nWJcmjKrSyaoZXPgZR3yfukhd2r9XTNXTIhoae5i/EBVC6
UvEW+gc9xm9pzpQ4/wojFRb3LWMTkY5gzS5OZ+ycBXPXNMidH7b4kHkXjNnfmDluOnwNEatuqeqy
19GOfqA4UHXH53HA33BOt0ijKd/ftuDGSPLsRYULkTj1yUxtIC4EaaAY94tyl6puIe4tyZfEA7ho
JziuVGNHLOf4xV0lxjeH4Au+i+p2eXZI6SN1TnFngFSiPE5WS7C6wbmI4o1BaqTz9Q7fU61r+rml
u7+NogoQ/YISgYJSnWe/nspmqITTX/cf2fazNP8B8Ezir346lIAmYOUiqs4wsuF3oL6vwSXIYQNo
etfUM+AmXC64pgF2kvC8cu9WrXdnGXKeOxtiHH702X2UbirJY/JItnUeL0D0GHz81uv+1Ha5Md3A
JjYRbITufXT8KfLq0X38FjHAf96YcO8ZQLza9mHNXjBjYbUxHUYmeYMNtaadKIc3cgoiEH6X3OxK
cMBLfSBoXECcxqKJO/+C3GM/CShVmrxBWh5G5fqxiXCx7G8mDnpnS13X1Cz8rKqAvJRHAg8ACw9N
i+G9dWEhAi+3UIe7sqTLKVLT4teQBHWFhrRuJoWebin13Czc0vJMGIQhysy1xTqCAio+vJ3qWqE+
9O5wCdkIGdRxSRSEAYAX2XMQPnOkdt2Ke5n42xBXxx6Az1tOBcD1kHZufsTxLnGLisMR/jKxVUIU
s1p/BX9McA7C94DJf/eUOzxxQ2zOukp1D00vGikFKU+ZF6dZi8Go3E0YVLPq1EM2HzOKTwh5KskZ
7KojdaKoPWGmwaOgrZEuM664lu8/I0jDjIigJq56dWcyLMylCbRB766xnheQ7VIGb1ebXrbOEkCc
8FzLQqnZMT8MTNOQ6VGs/Ni1chLkyAaOGIKGWJuHSb9GMR0rNP0QivD8G4iXfEPpYNMFjEpExRH8
pGVUfGSwdpx/JB9ZmluoI9WkKOmSxOj9RLmhwcPdDWPifNAkRNjNsLdxFlvlMoUkV754WPKMxT76
9Xqm5keNvnxrHzhY5wfrLJy6N4z2rJodK59mzAB5OyFvfAJjuHfgBTMCh/PqislhhPGAarDFnTvq
QLyrXsxxs2/8cYfy3D6jhjQCYKEbcmbTNy+v/KvsAFZVOEeN1TyEcqon0XVgDB3lP4h/tDe+7GYo
Synq4VBViLIE8L0NFPxZl1UU8ULxNfVj0Qgyh3T1hcH72zw/9i4Uh/KCR/LmxFvpSCpkxnY6Q+Sm
86NYQnBhCnhUaQC6p1MG9nYIrExoK5i+sNKOTxONFDDg5tE/EocCCo6p0x9gW5lAMImuYEDOSsur
nYHjiLsuKxGXx0PXfQCy813OA3epeY5pnoEYMEZZ1PV2A2aQ+jVyAHmMIORYJA1QJaJVSxT3/EkX
TrATgrbbafuyl2aZUSc9qAPmAtqFVDkTetz/IgsW+cIFEvlrmUMaohSSCKCfI/9sVsSdstZ+CROe
3OubNVAnEi7HJUAh8zDnxDTysU63bLUSrDEpraCRTlNICr9zb56RZW953/QNj/zSfw2uvc+KRK6S
2PE5HcUvKFC8vdnK9IpXVcHzCOzVe/inJDHkqolf94hYVHk4B8Z04xPhLz4A6eGc4iQljNWyJ5cj
WOW61qnRMinemppb6MO26AOVJTSLpF8U4Ifzm5WmzUOfMT9OxoVrFKS8ZJ1654mDMNsrLd9sBcx3
p8SDm2PyBkq+vQJ04cmYoUUa/Dkj+zYa4lO1SHsIA7nW4PolVS0XJFIsiKDCo7K5eeKVAJFT3yoR
H6QB0f41qxEOqSAsz1dDA8m7y/4vNW65Bz+LracHeN5QqjgfYgxBTFdMWG4YBgoGSTywlAiHvRdC
HXbUaHkmJ41tEGlAXtQgBrJ19+ihDLMxLSMsBdnv4J4O0YnqHIvvkHY3HVPEuZ48Homa5tU2t5B3
a2CZJtIWhnYnWb5N71EExu1dLREw/U6heXfyofeqlIRnmXOOQ5e58L3ZGtVRuOGujnnxJ1fGiXOo
9zYkdLWnrDLSyEi07Rsad3qSC9kSujVExg0tpKCMtOPrVgsW1BaVre2qTVtOGFqOOHzyecnqUHgW
nAHU6Kt9iODuEbW15B/StpTt7vVBjQR3nLPxpjN0HvbaGm6ehST8LWqXAmWT4xNML5F5zHv+jejF
A+yHm6XqMSTdNM6qS77cHgcbYSf454ZeOIz0eWMlCOAms5Z+EdSwiYGwTYjubmKx9YVHSenVXMNa
aFZtlVUCZUNpT0T4V8+XVm3Gd/2KDaXhK5ds/IJGgtkA9RcjAVsKU28gw9OyJM1zvuq43/o2JcbW
CYYl+rUS4HpEF3SNvyuzAmtjlaOnmfUJUU+d+0K8wu3g93stYX/bhWqzNBovdKqDg6A/Fy3hLxT1
yVMZhuSnGMPdoi+272HBsq8ntbzgLi1msKZ8Ns2zE3Eg8y0kGUKRuM2hx8nr1hu2AYLlMREgVt1O
aLUCp9p0KkIzIt/btqV9PLDn+RY03HelNlY+3808TQZQVqeQg65BKOjP6DbtdgYAw+AzqcG/2HUl
KKWsrh6d/YdSNK/xlXB89jT8SRV11QH2abrGdZ9Cp0u0+ve1pQVflsdUfGkuAxIW05CQzjk4uvPb
YWouOce85CdmlE9ILf2HH/9c9C8/PAIw3uNTUM5R0ERrp2gFDwDyeWA6ccZ2SsZ8SJeMdivtZk+Y
ODWAW4wRSJhwwuTYPpEMIvwfke8NzvoIc7e4jtY5x2sCuUxkcxpd8+gG41SfokKP6m1KK97TA0gn
uDjz3x3+xettMoqFUGI6m3AhYfl8UP/I0HY9a6JcWZQHIT/OGOcZFBmphhzzg3DUEUodSKDcKL8I
pSdGTDHjnNpKJr9iPQBVoYJnBx31KIs4Jb8yAtERMDkdgNe2yh3VfQ9rWhp4V4m6LB4AZkMknVf+
fddW6ve9M4sVgtaglvk9nkJmDF7uKF6ih4fH9geDASO+x2dVnx/AUh5c/eM8MVOmOw1dZE0TmuvD
I9eRNIjiryj2TiJjf90tqJntXAP4hUASrfCMo6/U7hakjI2Yy6aQA5GAvl+OHbqUU1lGJe+RuuUB
wNS6mq5uOmtvHT2ZOh8k8/rFm62pgfEfliozHNf+Zql3NvlCbG/IxOn2sdJJN8+9wRdQAqn1EJe5
gDeJgGNubSk5CqNG9uKhxwFA12ICU4sdxBNJyoAC1zPI5WshJIPR25p9Yg2xQUUhHS00tBP4EfQz
2quGGrsba1TetGZk59hsSzA7wkIRoOdI3nlqTDxav1y8ipI4etwWc+tmp+AjzaihvMYym6cGOrYf
E4N853mlj5ACtTBQsTzHxQfB5H0QzQ5pI6TvxnZcaAFo2La50HRI6J8WtXh+CgwZS9CCvuCRsRwD
iCloLql7qEeu3cw784UpGpFu3mmTbLY2q3baiCqWIa0mqFX1KngbXtBgdB1z6CJZfM9GXKb54LOA
Xe9ew/laMn0FNbTQJrgDceSy9muOkpUHpbUSV3yVSMPmkph8bE6m2Krq6IrAIByp7PJcHh4mJQ9n
fosqFW/TsRoi0COMna2qPt7rhmFRaP5o9ts8mrnTuQyzuTnfSJxzNZcPqcxWjdvMYkb+Mmb/Om8E
BGRe1QPg75mLcYCpXk6KS00YGA+ySartPqGgqRhwVCH1ItOL2BxRGAIus+4bYMeKMq9L+k3tNa8f
BjIfYDji/CsihwbZqGIc5cwO3b+ZTvxUSgc2xLd60cbQXlxPOTw7ocRNA7OKWcIw5TtW54XPM7QR
nhKjd4W3g4okdL6FCnbRZwxR9LjEmrxdgz3qKTG6uJWvy95RfC99bVgV921UlHRWDUKiMsSqZWYD
nvomrSnQ4EvVwYcDn7xzoRxx41XdPUA82ntz1V3uZ5J5SniBxRYzHDDwjK8IHXZ8EOVuWpE4Wy2X
j2vUGDN4aJyId9EKfGLUjH2w1HTJvzh+9b183yjf9JwVZlRj9deROiEQ98gLlsXSIhBJH0yqPaGU
3sbYhhWNakrr+hKwbNGc6LhS11b84NoS/K/JDi5FyPG5+wTDG5/gg+shhYMUUmo+ex/xJ1IFoU6d
0+irA60+aJ7fvh6dDE0Qj4H+Ge6Q3UDOxqZg6X0ATGIUCBEgem3tRNvt7aEBPEkPbuabAUPVL4ip
rq5Lr7Jm6EgDjS6JniXheEuR4rG2ESeZhqErVDzZ5KWX55zpoeGQMXzNpPDEUyk3uMvFO9OErJVY
nuJ8crlQqaXPqNGe689zsBy0fr4z5yER+INtE8L2SPueZBBwvlmu4j3mfInXOVBc64kVgmU9cgDf
aiszXBymmkunOZNpticU2Dac8H48Cz0dpuRHkT07HwQfDPioK8PrHbD1vAvX2HcLWd5YRqmK6YEI
ok75ZwDB0qCdwIygvdTzp15RtkYEemw9apQFjQuQFftLy68nsmObjSNMA+cHundAlKC+DBsszv0Z
/pRdp/47nIF2SdXmN3nPOTi1WkJYm3OTw9rialU/TU6HqV17eKzVBHHXCX7tzaFMD7AHNyhoyceQ
oMXFMhurZgFyRc//TH3GSk/8qfGfnwtErdXh50Yg7DCcMDM0JKNbC8K/22ToVkc0+JNNsB34sUrY
8Xe7//Mewjcxa3amqQb06l1qJQRGBCguWi47Rwica/CTrv5UHoZbZlr8gLXOyalfydupnjoBhRj/
zb+S+/8jQtXQbs0780FIOAXIYMwXXsHpxBIMGa/5vlQaC5MSusGZaDhJj3LetxhYM4x0sMEA1Fxc
vvaHHieHwjaM+odaMANgWLmQx3EO1iS5pRrOwqso8Xr1pMCA0Pup5rq6/VKzfKIyGzqADpUt5v/r
0tzed16mqHqt3NqwcGM4EFU4E5zt3b49s6aSAa5mK9CXZx32XBep5NIpNRjKylwjaBDm7GGIhb4m
KWSk4G5a58SGNyuv0wmIG2kRtp/HvhUPT2ftNtNtiY99dtBgbMeGc/dPxkUaLYeB5lgHIBOWJrK5
ZixGNcTiKBPzi+7elXMuufdvmswaDQTxxrGveW1JAb0nzO0i5W0YdUCWk/iN55Y/PiVJYgf1TJuM
2/sxz6B2++ApeHT4OcRTl/qBMevkZSHJJvfSJMHkaitiyvtPke6dqHZyXyevQURmVeVyEyowo4rG
VhkacRL1s6Jg6/YH2WKWknfcL+Fn25ps+vK/7+YEzaQRRABvJdlo668aY+Fu6wfGEe6P+KWbgizI
lJfKmUuovxBWL/mGb1TFJkx0goBFRn776Ue/h38YqvAl4Gw6M55pKNFJLciR1S6ZXMD4B4sGulN5
ugHhRPv8wFvtc/YDd0GtanEUYgFoaW8E35y8izqrIXPN1Fg7zgygn9aHsD4iSh+0+Uz3tzkaxANQ
v6zom7I1rDyhRbrSJRg0pIp/+9dpwQJFHfQE5E6BXyopm/WGWVkjmjxU1akk/PFy4j16pQmhfJPJ
ngl1eBTJtcDXJMwxrBwHCituMbwtz9DTGdLjUzutXy/LDoADpQmvwQUpwkNJQHMKNe5KF4eE1ajF
9H8i9VPLg16ruvEzCRhdK6qUevLHeXMLGhT6PqdgH96MmSsT19bdueMw27hy6hHBdMq3b8RD0JbC
rK2etrbAnG1QunXFDaT6NTMkSdZMwHM1gkXZeozOLQOQzIcmLIbUM4SwRQPvYBF22tmVbrh7RhEn
f60RRHks3nONRSD+FjzuJDyCAl3pEMEd4brUvUrq6aepDTOD+Mjmcuomxxh94Gh+nHICWZqybO6u
HyR76l5nZksByKSh5JRZNoxw2tuz6MUE8lkz2ukozHBFP4J/s57fAchg5mrEkHQUofPGr7OdakJu
44u2w/rHYQLXRBRBIgPR44CGbaY+MQN92SFKu9FgKMOOoH8+Xa1xi93vKB4p0EXmwwCTGtHj/gUu
0Z47qJE3qkhUKcv9dYiuRwbxQe2zoT6Bl9+jGUvfoKkl2BeekqoVEBWi9HtuX/78op6EpNB/Td1c
IoW5c+wUC940GKTkQJezYE9JxYePibRKtURiAUo77EERW4nobzDpL9f0Y5BI4uAE6IlcgfXFv23B
HGMHF86A5sX/zM0WlvdXNaXLjq+0AmDNcC0Yur5++N6VwRG84DvlzO0sWOPWBSxzj+8t+jI7HzEn
+Tl8tOhvn81MusYJmljHFUpWXD2v64yzYa9pyzkUf1bsVrRytp0+KyLgCXAWIRx6TNNKjap7438N
oFVUW0L9we8M4n0zXq6ZfM28TNaCtHDSEyovaeFsYWDh9F1vTzwbigjlBb1Qf5KzjTZyXGQwlJQH
V6yO5nwvv8U/fJ8S/IhFNUiZzclkEFbvRMuV0iTCNvNXEPoP5T9Qvrj+XcccUR30VPUwRUXkhuTO
A6D4jRyRJYI5eluL/y+J8soEaTeMujucfDYYfWFoNtCyyhqjA6oms+WN3KHIrMD51hmIzxAgMTJl
J6yccb0JkA/+11WUo5i64Z/NIBfSwJIdVAoY7XnfXmX/mM29wdnIH0QRp3ZMxK6MIu2f4RNxFlvW
ISYClANlMBMyME9w9kiSSOH3jX0rpirNnYw5daXjsEv5nWBzsLmCgi4S7WLdow2c61OQ1TmNkhDW
2JSBao1jI6wwXlelo80XFRBtzy58cpZRKVsL2/2KSwqsoqJMADqdHT/1/DZSqm2iOSdyXbY2vKA5
Ha1pXLNdOhask5anvV/zh1lhI39YTtiaR4f5l7nMlYmM07cBcRNMdqidSoRJ8QJVf2LgmHsTEEV1
M4REZGRsjhfPHs1d9Vnxthl53/G0x1ly+5GA17eEgqKJYcrh9ddkvNPH4gCGNy2+b7QrT09MhXmO
gGhgGVJhjzhCy9qy3xJIr5i1pS4k1Ve+L86WugpfxAjRkP0DdHcJ85On3nPNbnRmzk89LcsSozvZ
z8RTkhTnW6borjkJIBt/PLnMxuvXrD0yeOXaJEq5jub5/uEo4fQx3TGLVGAOgprjFScHnQCXmYVy
5M27VX7BIws/h+PcgNkz89yG2H8/ydIjpW2uWskh8AxMZhudP6yCTDhxYsjTrYyicj/f3x6wDp9a
dVP9u51bN/oGcRt2+af2OftVL/1PoWY9QKmBVLMkyygEzSnzXEPE/oVZ3lEh2xmmaJYztlcZ0v8x
phcLoAiKC6Lr8k9xIAQwWswH/ECg0n+Tdtu6uHR3r1QDcfAjOlD98biABlT1+8YGllUMJszt1p6c
+OExecdn6CruCExYvuciCHJHf3eVU83txvDCpoqxH37tBxmYqxw8g7aQP4cKuEWLoC4RKnYtMX6T
vjtA+SfLmlnmM9pXb+elx2K5Ph/wXT5k4oAbONg9RBardf+7GryN0XbucPdfXCZZTy3aPxgYE9ki
Hw6i7msfyPs9EWNvDKU7U91yoSDtyJE0rz+QkOBs9hdYlBrmOlhVeA+W1prEmtovwJzCIrqtuxNc
jtJ8uMlxT80YkAhucOe17G5N3+GEEpCmYFYhWswO+AZDOIFGD+TXvtW8u/2BpgPlKy+QGNC0VCiR
v3+6qv9P3YNmIMVpWXsD7bF8POvSn4halQQM7O7WU7H5fP5X9VgixSpzbQMHZRIdBd/pyqqiqfwy
7hA/nnEDKGUlRxdWz/zre3FP4lCUfR43hsI5D8VxFvO+fIPNalihNKyqXlRJBphNa7bjsvC2c8gY
msGZFCwUvSLsZ8SlJushgaowmb+aHtblVp/nTO6vktwbbzqW0kaG99BFo1UDXxEepo41JAOzd6xa
1uqDMtuzQI4dxpUEre6w9C5G0BRRNrUuWVa6MYXZJkDUae00la/P1izukL3x9GJNCZerXJ6/Tyi+
hm+EBuDzfuT63Co1l+nB5YWr3RpCZ+jFnmCj0kWyHWwDDEX60ZD7vicxhaON1TBsCOOpAlRbttVL
1UXdetsC75VJKX814bdzUakfh0/qgcwu6mZc0VCACpW6Gnb0THgs32GWcTVKgbN7K6HaVDWb8q4g
z9I/tXXXB/VZZWbCXxj5q3ftp+XBd4shBi4uN6EQKzpywQY+4z6Y7+Z0kJHsI6rZ/SLXgi135c+6
xWQhQG1ZMJ33WRgiaxU5rlftccCVhcVJKjoEdSmVlkYhwt+Ns0VOU84POiMyHynSs3YWdQU6Bn+y
9YaMwnQ4sBaVI2T8pRaREgrivmyiyAnhhgtf5s7vPvGVFrL6a3f6R/Y+g9rmKtTJCtbr5e9wF5Sf
eA26f+YMOgMXO8wb7TX4QGAcRUEdk6+mxfjEZHS0D+PpJTv3Zz0U1V0LMTRRrGntdUeB2AhCMHny
1RlTcTHB6SL5N4YmcTolQFnz7pOhIKRfUHhS/40gpTMvzA4OsIucWZ5uRoHfFBS0jlvL9weOCdXj
wnSULOc8mqYtf4Eu+hsM6Jnutx7yZv9E53/l2ZTXikYVDXY/Uhm8ErSOnHpHjt2DmasuxGmcNCOG
8Jmrv9zQo8yeNryGoXBOqdv7PBxdmAv4r4v3xQYQaqKyDCHYKqgp2EuhrGTUJ8Xp1xc++BUcffTY
1d1946ynu5XHVPe11zgO6G9J0mrZjHE8rojbgK/hKBoItzNcyF60pvQCs2JuQD4vI3eOeK4RY2/K
hyr8Anqqc5i2y7DCYVEyTS1B0jttIiatdpir194trXq1W8C9kLYevDtm6+qReOnbrcgQ102VH4tB
Xgz9QdFJm1xNNIUhfZ5uPJjCk/B2OY2iv3lKYHmV6OZaayKxFbRLLeLmpRWmq9LbkOiTg/ADM58h
yh1inoRy/EbWTIl/73zDooiwPWjGhf+TZYNOg4lr7vzRSRP7HT0LbsE7oPjpDKX2E8aVS0crcuKr
3vfRtun1fkxszr9shFh0vurLMYRD9uEL6Iaw49HB6I+E9M9S6RqP0AIQvhb1QQDT+uhFrw75cK2j
HokMOzEMl4kkBbwRr6bmj1AQKcrF2lBdX/FEJ4ZFgYCrCGsrXYmoxfOo0ooyO3LH3weaVpLpuXnd
YNT05Ouksdl2WrMFcIFaHf4qSPDoWb9AYsT1/IQ5MTEMHsKvj6kOOsmirLwEDnZVSS9xWwXbz4L5
75yI3MAvh6jE+sQ/EGio5YgQeMKqZxSmT/sOtdupSSJxc7L0+wa0ofKbkfSaRRJHqS3IkxOsaBtl
VDauM1vkrmrSoUzhS8WNSdfBwI2sAFnLXm2Fq6ZYfRqjTmkB7htxh6WLAA4yfsdQkfUuh92gGyIp
ojDq0fYH66DqkbpqiZG//4bZBQquUQGr2LLosGQJDb7NRiZ5e2aZ1Jp0IZigPWmce3/vifskWiKc
tLBZAL5MDPKdCSyVjRQj+HVAudotRW0Iaeldn4w7dyPnXtO6aRusUQ/MPWL2d1EMzw8GnRs097Ca
Pe1oSEwK9Dr++/YYQ/BAC1IsO6VaCQ31YHLbUr7JpKrzF4hbsourbSxwQoNnn8pQeKcimfGZ2IaR
TzgdESII6Iczjcv/Oas9xgTIqRqv5TN64pfCjKFOzkbcRPequtyvbHHlkwBp5OZ9wVjNdeZhlHi8
XDbCuO3RV8pSTzPPO1OBNCR1O+G4JDv1JZL+paWSV7uLFURB97i2BVrvXrwgCGP0TVMB3bx/4oNt
E9qA8eew3iIl2bHmXZUN6wGISHOMv9TbTxEabf5qRMq8HBs9wvvjb9HRZwKJGS4xmVKW5z1Vch8s
n4UXhxeFJmRM4KvQ52zaxdf3LCQ0RM4zz1MyN1NY/4hlV/uBpW6ZvImYJ9cb+QGXkzcJndyLMMXv
fM2mlPDcQpvE+wbNsB/taXTl/TZDkkmydWnmCJt+zcLGrED2Ya/OieSQcxFt5Y25lsxtMjzvSq03
yEPPpB6Fg6ISsIA44ygpaMN7YeHL6vGl9KjFuz0CPmTEeCjm4RVApMTU9Le6VIdtM92eKi392K72
Gk18sDGjmbPOvHGVrm9BoAM0Bsr3Sj3Uc2T4WxerKxlMZ5w4w4+JOXOD/MfUVgOrFyUHBthVcVE2
AFcdNK1XjsCeADn7drCksbLVhbVwvW8VCADWLjrmeLu1/KgORaP7KmDf3H2iKICiiOz1/JgQe9+n
jReAFsfcr3cJ58YfExG0eYmy9V0EHcHMlwrj8yqxshdc1lVDkt58619sj16/jViKfQzu7jTYY58c
oObfG7v0r+0s8dr1psN0DsMSH9ChMAr8rqmQCLENBLJ6HuI9xZfdwqbiqvLG4YwAgQTEZOERu2yg
6cqtxcc3P3b/PMa/C0MlDbmAWAnNVFbByiOy6cXlqYd7E9fnNHnPz5kRbg1cO5RwR+Ckb3MMxFA3
VcbkyUfNyzD5nl4qbmlD8zJ2aZUqGDXHDpWbCKdkCFvOmlVpAAi/mxCfJZI+vYl9UTIpUepypenf
8rSGG/HvtSFjc8bIclo3yLWkIP4SS0Fjo4pYNKwMUw2ig1FN/yegUZuVvgOAEfTRKNcWO8XQgg7B
n+h7XrXpZpUsZwNxqhyvO6qlwer3AMrDuG3WUJiPC9lrRxbOer0cwi/gaFS1qhTi+fQeGqo6ROs/
hTqkxfWkY7u4yQvbqrH0UIp3woDj877mEp0CoBWjsKh71M1QzSWUT2f2odOkaA/BPOLR56IlnMZ0
St92/BPhiniwpfgzEjD2y1nZmpGS044nmfwQSVSCvgH1PslzgNfvx7UxX01Ss0EwVFAz6od7DrKt
8q5O+LRHh4rVGgeXTOl5cNetE6vpqbxDNspUpLVHek/1ylL/Nfg8cwKRfZnefFkKJcqyTIkLMJNS
vNNjarkhk2AiJUJWg3wMfw2Un1yLJ+PvuV3tif9rdDGI5FphTeDGLhjkVwNbpgUo/q1TlH5MrjZD
QRpsXrHsxfGe/Yc7vRTVmcePyN3gI7Sj75jRnAEdkkwG33n2ZcCWN5Ng+5kjpzDYZW0U523NjgaN
5BxWLEiA4zIc1HxkrSaR4M3VdLlgsC7ox/rw91CP0aZ1cSyh1NSxZHqjeAr7ZNWJlE9IbJID6bt7
ou0edndhdc+Z9hR20Cl9Ip35sUNUsjPeERlO/66M+Dz50NBrlgV6rb6pmKU91MO8fJHs4KEMtMIZ
TT+ZR3DXWZT91LBXfFG2e+baW5/XuM3bATnOUiLB/R0uXjQZOlRfPGMeylaDzRhpxwyqNXX73hG+
AZ7P5Fvy1q47Z/4DdLjw7Ks5Ka8d+dWnAvMZuu6p8A6u4q9Y8ve7pUMFfj3998n2povY0/WgtUgq
QiJ4Md3UCoc+U9G5u6ytMynAgKZjobrmizOAfTvCOMM35mTPPajcwMFxX6z/hnIPbJglhPrqaA2T
54YlNrPTml1X1m3bhIdRvsC8CCr1cEvDIB3/zeJ5nd3tMeGhRE+C3jMrTetwi3Gffibvrv2OBCWO
vlid44lYgbLWrRbNxX36wstbrqiOVHDo/6BG8xSnO00sjMquHY2pg4WC8uO1RIF5jgCQ0I3gwT7Z
ArHhI647k6mIa9gOmGYI49PB5TjDqABD8Z00P0XjMMWvWgaJG+sgpHo3kA7H5bklab4I1saFJnaz
pbqLXoD5vv3OPVuA7uIl7lcJabPvPfXKctwZqtJMePN+cvAhBMiBVVBgxkz+klwIjz5qhTIGm7mt
Hs6+978tpWKtf+FCzWOqXts9aJPb4ItJql37j0uMbBma2AlvIOShG1pEOuCRIwgpjyvlLr95Mprm
OgewR0gUft9UMpsG1JzXHXodGYu5I/VzSx2dcFZ2sQYAGVcygW+HiJdQHkz3Airkc9pAuNvMCRdK
yeAxUnnN1D1i9Cx9CMXNC2S1yurlqwK8XdwboSKfQKlFItFITqxrmzpbMQO2EBlB2tzCzU86ZRJk
iBvpc6XkNK2HYkVNO8Y5hlUh/OhxwU4PfSd/zAzd5SJ+eiE4LCbrQm8PYC5RiXS1PxSvNOiPXCZy
H/SI+xjVxhfepnrmXYxFvCrde56OUAk7XRzYoyevYF9zVtY2947F8h1mONGk/O9oa5040FqkyFjO
1UeD2afAA+o7vTtdOBNLfrwHZ9zPfWGzvTP1NtU6oBeb7wI1F2wtAxlHB2SkCGKLKfc6I7ZAlYor
J/DKNj4zjjsLXBsh3c55j2YEI43T+1AePUp2RRnXdKZmkokoeBoiRgnmMcFHsxcno71Ca+yUiMtR
/l7IYBPX285l9P1HsQo+ccsaZuq+B4XvwxORqEsfJy3fUWMFDihgkxcK+4aAi3BEb5AsHh8I9+Tz
z2f67JIZPK7hkA8jPLgesEmLZFVi2r5MA5p9IDtcApMzA8c44H4YdSH7gSzi6Uyf24zjpC0u3bkC
OZHOsufJEd1G/oYN363r+EbpFVV6kCHTI27TvIOawrGN/6O86HX0xTYnT1Otc1MJZrQXIuQrPP8u
AF7PJTsYF4zDeRH71X3rtIiIPRjAsJGNyP0tP8evTV3igcR23iGXP8I52K7kChnzKL9p9RizNPg7
oDIyQZinEuMKu+x2FmAX9wOz1eQtBZs8HtUc0LQVhFbITaRQyagKaw22g/s7nvokukhM8g1CQ8dm
n2LXqAafbJlY58w1VaCGAMBpWoEbXjYAjtk5/Mwvd6x+3mwkzDvXmHyTgVMzkntlokU1AxdO2kZB
LgJZtXOT8IX8xN9kxH3ZMPqqR4PqBHYzLlfqDiZHswgrPcVaRTSQzVn0Vn3/w9vZ06ccsrcvzIv+
UmIha2R3nCSsNc4FmlcWrU+wxn6BWn/Uel24Usgj+H2XG0VvjHvUHfE/UXi0ggbvWTYsekNOiINS
9HhjNAEyRpJVnDCXggyFMmwED050IIpt27/C2/22sRWhKiI7tqUGV+/TK0GFl87mZd3XUNfCQrli
ZQChgx8Xmts/InEmT3TtLeVcDyWlUO+7Z/xN4WuizxVXOSUzK7IBAVnuHaEX21BBS80eqF5vKDis
akCw8ymFc/7wMp7e3wUQ3F5FfsO6ApLsvtJkferoQd52gK7Rz5+L9Vs0wAMJAUTqYcFdw9fYE/Lx
lYYSWFEwD/Wbn0/ctFhDMs50VJk9LdKkPQiZBf+kaJlSslHoBkdwycdDF0R4Got9Al7oCp80sK/0
llK/c+2amanJbWr4N+erolkLDtzje8d5GwVqxrjiacOKRURmgq/1G+5EcXgJ6+B+mwqrXsboKJ1k
5q281eiYUks97zBRmjrYp3E9EXmCYJTzAMHXDQtakoBT1koGwcMAnEW5TG5RdVBdh8OW3LOpOsKj
4N7V1G4VGvE8DUiTNR/FDL5GkmEmnOj+6GglfrbIwp1/1Cs+MR+tzqVPGHOXBom8BfXoPpud4ChS
hzVbWq84+ZIxMgu0j96OIrYJhSBzjnSutjkbNaGn1DU7NXltpR7JG4pM1JOCdTIvnizBMAXa7e2y
+gAO8+AbMywXY9Smn8S90eG/6S0CX48JBgrViLJNa4UImhZcB5kkF/iFavUJMP3uUrR9cRmT18k6
p5Ct9RmzivOzyOW2B/vuxEc8EGUtAWgQ90iPsCx4UfJJ0gcI032xmChFAP2BykhiiNWjiEGfJRfb
4D4URtoNswr49VjiSoz5yOuQay1LlGHxh+jG7R7tCv4/f8dWxVltxMUSFDdXbHZRHonfpSHZQYjE
IlNlrrecKBxVxBhUIwdcvBfxO4T7o/2cS40s8W4gujKIWQZdL8qVkmcJ+YSpbFcjxkMStR/wwX2D
vrx54FT35dKH7fBqSCxd/RztaKW8DU5XEw+lQCT/1UYzMfbxph1AePzxFlSNNIVwy66oJxMDwqXg
HbKiMhNk9koEsOSuCD5ws6rC36aDSj5voLGiKYtRnLoLn45y5EuwcQ0BfnhPOpFDVGDluboN5dao
oSlm8fOz4wes2sw7/bVV58ffqFwu27XwerDjlD7+DLcx3kBWBQftuJ7rsvRTBmBOjlp3q4AjWv+L
FLtvfOcxyc65KjPk+j3gVPp9iJSoSZ2o9QW4hguB4UQaDuRx3Rs8V0clGkBW3ip1mnfW7tWm5W5E
f8vQout6m9D5a3SfPdwskS1Bx6e0NUrecn6sFvF5BijQMs9N5ZIEJA59G67zL7+IQHMMDAZl+HJr
dt9Yf/ZsBhhJJvTSA5uTqy/s7YFI8yiokMw2LFsscrOnvZKkd/ELqKIlv14WPuFHCToJrvjx6X+j
ZHZQ1gYaCbaj7HF24dchI9WD9pMfm/cXyRr+41RFBBz6VOa46NndrPKo6QaKZAurJOdg5bmCz3h1
TZD8TPi5A11jO+XuquIzPl5KWKdzcJLUSSHvmWwfMvHxmYS8u48DSH0n/clJtgbO9H4l8aKkD9B9
SiHlcu5oiedJ7075bavmbJ7bj308ncLmjHNge5fvAavS/K7Sz2ePA9LQSbXcZeP4AaWeCBpI7eo+
5aUZcQWYrPqMJz8ulNRMFigAwYAS8hSIvlNTosBVtQBvRIVWn3RF/elJwbnJ9tp61gLI3Gjxv9yG
K3S86/cylUeu2OlW5vg9pTIn9Zf7tNk0Uo6oysZOrRuvnBBOqcDzt01I9rHjwaPKW5sDEXZ2q4b+
PKK0z3dDnNX5dX+70e00WhC1ANxt0e8gtOJdiOERMb61rYZ2madZ+8NqVOEcIIieg4FuPqpZm9ZZ
JpKu0NzjgIaC9bRMwj6FWl4ogMN5FeZWV0a92DO6DmGsiqihXs3ZIrwOfd4ADVQNdwGAEvuwLujp
NhllkGDYMG+VqoegozYsd6m7tZYTYzgeVbKoTKEdqU9jLFlF1wKkdKD3a7qBfCln2Wuxli7BvLv8
P7vIt0/dg3IrqEv4DpwApkppMSiSinMzBTvoTVFSgRmRwyb8KnUpheE5ripLTH+LpR9DJzjICA/m
6UHOe6mw7+nOYu2NbqNmHVd/6RThRQo9QdpLHczxkzlP23/+RWQiyUIR9Xb6oBO6fl8qW5e4qboV
78+w1WIiPgodyjWxkISnAEuW/DAH5qgmhP7lhR+0qNfPN0XiMqJRljewnb0zuoocMqYgTSoU2S4B
fFmZLYrJpFU7BQ4qvRxHRSruW5fkr6lhv3hD711Pk9Zn/KbHpwlAhz/3XjCyFx0DqqiMgau70ERs
H86Fq0s7KSjWP5w2O/yT7QMId0DFhoZA2QnDt/Etg2Y7mru/g3LfOlBo8MBbRKydONmksTUDOjSo
4ZZkRYCzFlEUpcn3RR8T5G+Q5jwAJepf9rcLtNlHDrk2tg596J/yC9PrmroGc2CjlaIm2rJiQEEH
URyPopRL4mfVNZwAg+ZDN36OCZkITHl4vh3bgVi8M3JehhBLktEZgx4zxfAA8SJXZXmVqeJfHTv3
D64cV8LjB0KLx/5ydglkF0yL3FyVd00gi5sUfSB8J8B21zu4lF/0WWTgPv2KxSNfS0HvoBuFSZhF
wcr6UWVR8eCnjNtf64dG8U+4LFXu9erLy304m8mGsJN+GjqVVije2c2OF5QZfb1l868eUKh22tro
FlftoAg1qb4NK8jFiOMUBXjrMj8Ifw91nZNOezmTw2yxukQYDYhK+5SZ5paNM3HX7E3S9cYETMog
Cuk0Ei9AZKoNDsUj0nnfiovXb86D/MXFdVagduQGkgZxnJBGFm2QRAKQQc02qyArei5C6cgWx0aZ
Za59PJLsgs+fptgMYg4oC+fjsqZXLFO6/BffNPztGxQyNdJ08OvNP5yxJE18pECwA3f4n0Zzolqb
v+NFJxDN8XTVWRBUR86TsLO8ueu59Cn0lXdoRs5rJ3WKtCWL6WkCryXN/xP8tvFlg7NsfFzZvlnH
Q26fo9tkJNIIuJSx7cS3QpJ6IKDavTQuexi8S+ldlw9oMWOtiOYju0e9Z8mXyG0T/eRPzkrvGPGi
HgpMsQv1ONoUHx6I074IU8WYhrtS1k3QkRaqWZGmknK8RlnzjmRfCYpWH2tfPqiTS3ybVTbvAWbu
gH3iqaWJaVuJfSjH++BwbIFvxwzYA/9vKhmEofgEAsbr9EdtxJndAztW/DFimC7nCOOPDun/2e1x
7Otv/IET5eEmoJ6lxghVhpHNnhC9OIL9NrcXhP4vzlDYLjLm8GfH94rDaz+1zD+ch32n0VXrgaFQ
U0sGGxtPze37vf3LYWC13CC/AcUFR4u5yn2zSY1kk4mbGhgaaqEGBhTAfnR6SGt7Wqk5OEv1cUJs
N8ykoY7MD1qHKhvxAtlDdfcgXpNhIK57BSGCIoCdLidoi/Vb6OCzDi5mV1m5W9qem0om3CoLYY5B
H7eZEJvW5T5TC9wJ28HeWNy+Wv6aSh/K+pryKvrzJLXnKTYaO9tr5bsamARzxZQ4W8RI3RfBxsV2
vr0HS5vj6pycWtxIOxCBXhG2W45VXRpSdzKTk3fgq96PDYTMY/STH/Cf8WYuoEa4c7RFGHj6oXok
52hbhyXaglQYLVOgND4AvGQci/3nmaIvNAvsKmrqVmjn92X8TvQ8ELc5dwCNgvTyzyPFBaoBuS/N
YeF7r2TvM8uLXtWRibNLc9jntDgI+j+PC99goENB3E6FPvB2ZRh1RCRci7fm5P/3M5smUYd0CwNz
h8JuL1P/JSs3XTTOg+ytFlqXRce4oBdPWeYSzN9ZxncCC1RZInGd9I8Cb/16O2pE+9WAYqWtBXfT
XNjnQEXHuUOb8mwPoFXAxgwsQF9jv41l4F60tyfOunaTqH4XQxHfE85P+w07yf8seK9TV0/AYRL9
m2jG6d6K2CZ21S5SM2jj/3OVYesJWtRTY94g8GoCDFCxGVrWzYDJpp2N+ycSzrdG9mO++P9Ko5RD
C2kxqnm1dAlsncm+W9BhF6vAGIlhLOLXchV/H3tUmGnQGGN8KQZ4dtC8JJXPO0Fi41uTYudUAFLc
2qAvPF4hyYPehws/LTar0yRqmLVY8sIAHJGSH4DcPObD/Nbik3czxmK0Itz9HD2UuglkgST507cL
ImCLyOhq13v9DA/ARa8FszeFHPHfr+gGY2rSuFRm/4Yajht3z0INSS4UIIWgYr6lATTrAG2f4qwi
YLpjwa9Y3tWURBGL/TbIof3cpj+kC+FXIoVtT0TyFw+b0qWv1AXH7Kog53nsFj+GNb/hOqeobgD9
2bNgyX8WQ7yxvjD1F3hbZAGpofoInsgfPhl9rx7fgg7t6sKBLR1Mx1M+2YUHwhgTXjBDLvcjku1q
gualHtwO+2HQnCI3DuEvbkJXRYxe0bOI13C5el9OtsywGp3xmS5N8ZrkM7R6BQysuKWffLNGSQok
yzNOs0L+5hfh/v/apy8AxlVdleOqou8xC5MeGkkJNWANnofYAU5ETW9s0OXvfY83SvUaPsmI293J
/CkCvikNN5UGWJODbM4HiqNUfeMzCIgYhMBTj/13y2Lb/ugCn4sZuIw7r5mHp6aIoBbTSS9k8mbj
+beBVMx6GsHUXYMBlQ+fXLGcXiSAQ5vMMt6KLyZVQL6nx58lomkbWmGScc3q6DGcGekBbxGpf3MN
/a7ymOoNVmg3DTnwNgz2cl+uUwZL0mmp9OCqrknOxnyLQI2m5qjoRIUVR5ZTDWt9xp2dhy2njOZh
PETwEyFAS2b12jCEuSYCQDhUA6wveiY/i2W3W29jeY74WTi5B8jt2WKHmPiRciooEY23c+Zzxe2+
CcA7YnC+5UW8mJqERJDiv0a88A59Uys8IGovrpBha8yPqgHv+kyr+d6wZ2YeXuO5TvtrrUFlMf5N
9Dzs0K/WCJ4PY/a0aYjkeVaWWuoaKhR47hCXkKb4Ydis5NH1g48svJcnYC8bBDJem44lnAix5EIE
lN/cmb0goDZrhfMTMp58md5wrYk9KHu/4mbkVu1gkh/6Gsd8C/4t4AzwbLE3kwRhaLHj9sTdC183
pHAPDi0uypqVjUZTVvuvN8/qCWABn17kd6Jg9/S07rdWiWU3b8Woe9qGjwlLk4yLH1HBYJExAbx+
1d9gPoK3yPQ1d/vMk3Xi4tpkI5WDMEEGOB7hgxu+etRPFkGTBE/x/VI2DJ8T/ON38yaui4zVRQTe
FpsegGDZU2zNwmFrd3aHQwldGxXJH7jmnYlTqQm/TogmyNJ/9M2mU/qtHdQLfHgvDmO7DqnDrFyf
q25vzuGO+m8ti9hK6XuotllhCBTRJN1XzPuMaFmJekBcK43nP/pgwamFxkrpQoXVNCubfO9aRWdS
IpGcqr43pDT1JUZE3ZVG0Ev9iB8FSsNYwShQENbOeoo6MG/hP+tjbhLNXyXs0tqrvHZWqlf8fbR9
ABvNXqtriybCuvQ4IHrjohnE7FahjCOiKhpD08+/4p4hH3SN/02ZAWBW4ap4vqwBOKszaNgKkXR1
y1uD0sMDgKUut81OFVT1MhrJQJzgE0sw8HApz95uQTxlN4WJTPfjYOzUH6uNjOlRFTaI6hPPekwZ
WWsYpa82/pFX8uWVYN8IeyPS2hZV8FLlvtoMEmNf56dXC0uPxfYoNzuFn1FUIEGAOehsHTFLSi+t
PyCBltI1EZcFjr+eowp1ffjaATQy9BKahpMFl0ybypSvg0KLB56USEj0oN7z8S2OnldHzjGrPZVv
l7pqtdHzrVysAnuCxRzavM47ahLhJf8jtwuimZ3kFH7SpFCUGxI+r6nB/+2qrgOcr3/Nz9SuUfur
IPaBb8XvicICi+NpQ8p9PCKDea/Fa8lCeOkyENmh7tmMHy7egTX8jJySIqqWhZuxcF3QJi/iMCp2
WTYJBlhjRiq6EUPx4FbuV2bFO8dxrG3MYOLwnxulooM2PSFnVs50tHGc6zo1hTIQw1nElJDPa6/w
YHaCH10PYWr5XA6bRNVp576ujbW4ehAVEtt68hz9W6nq/oRA/n+6gL3aJhXONESeebPIrBwJ7o9D
0KRZG8/DcAMwFjCebmn8AMTFHE1p/AMLlMWYHEFHR9mGYq5kE/0f28MjqY8AKCSgjAsTmKa7/bNP
js1Ls5aPdWUsi8AOOU9B27CsnEHcaQ5afxUD26Ir6fYnZ6CWAonxbjb+1KqSTcsGsXgJn9wexunn
IrU3nUqwJoYYBbrwK2b6SbD2OtpA4j3MFN7WYUEelil8+v9Dbk5CHrcfpGTO65c53/jGwxALcMYT
qZogpHZP2C1+ZoCQcLnhrz7ZxPvSCLVJzQtd9c7HKFjb8rltFg5LCnUWBFJ1ufxos5OnPwh8R7qY
iURjJbAGEsRu3alXlxG0b15eEKRhmvUHhpDHMFElR/XoUFg8YN28lWZceguA9a2r3QIXEME7nwQD
SzblTzGdcAjJ3eJmYM/6kjr0mUe/9sjp4K05G57GwaVju5ohtLqe3FlSuPviTdetnehtANp9/JDS
kElv5dSu6XAQMJWu6NF+jaUTesCjFzWsu+UyqJD6w8x4hQ28BbtyfktpGbGctDOCQapx0eK/BV9S
jw8fN8v1JNcfzCM9a1lYHzh4EPI/MZkSP8kWrP38zO1gJ+Rx9nGC5pGJf1FY6FRTWy8PX5uPXMBd
Str6yPwO29eNoIlVDq691KEwBztITAEAm2/1VaoVbsl8b9X2ei+VYKpyIA8oZNwNaQumZAPloaIj
K6C0eI7Lz6EXMK3Yqn8Fb3EQGho0z2LHS1tC5ZaxOm3eKSN4KesLcwEwQnYHu7DI1GixKItX8xiC
ugSvxd/OjCOVoekThQBcFGMg/d0Z/ylEJGjQYlm4Z0abcCVE5FZ3/PQoCGFvrbEJzJcAAQOEXHo4
+Sg/KmBhTZi+dzNCkf2EgywUBlwi40IzqG0fAyUuMILR/AyH+yj90mTVhcd24i6HejHDc4E0mCCV
yWC3PRKqHfCRtUlR5BAJNaortBLtjSSyxZFJ99Uo6dyhhhlyfZZJdn7If6d+lxqf7XgCBh+I3DI7
aVOaJQzpa/pxN/ZvL2RHUKqaCS/CyizNwYzij8PXu03o8r0GVTNZg8je3VRu4XCJlf2krP4Yjq9+
lqR62EkFtOA+gmHqpbC7lppPPeL+EbQk8XwzAIQp0zsI9M+guQlX9B8Ec/SAAClGKBZ/Ym77QEyD
ssnAhmQO0/wGk+zDPFjzmfhkp896NHlUnUzhVcLPOenYEBETKfZ9pZlWxIO+PoN9t/zf7WCN/ja4
P2SjEoeOMympY2PR3G9tFXpuQLYbTRrZshoAkx/txkvaSbA5ais17LSbvBQtcGR4TMdog40S6kK0
tWQ92u1yP9DIb4hOcim1gLq3sBo7TBYBNcIeyjAODieO74URm5xgcTtfBUXNLFuAD5IQHv44ejTw
oxBrVlQTg5yQHks0Nw6RgYFXDyHNFmPXNTGhFhn+qNwMpVM/hdNW4PhF//F2TXyVa9bdZlqUGiOH
XNVzryX5V4v7d1XE1x/kl7rNn0oPMoxxCCKdx2THCbFoHG/JLudM0XGOAA4xrceXeJ/l/k1+amzg
BgHLXY+bBdeALFDuuT1+4ximZFlT0v+laVbpeM70rrwhqkR69DVJ0ZLVbRjasfCnIs5av+BA4ie7
wfvYiHbv9wqH9C9GfP+lqWJrmRmziTH51pFVlTfN5w90f4wzeGWPz65rx05BqGUlGbxsRH40JSBT
ZyWX9DZL6CMhIK4qfftwOfCxIG/Jqta1xVuYn9gxPA1JWkNFfBIs4+rXFYQtp3YCoBG1kZkniFxN
bvoGe2R3apqTQ0rl8Mt4QEMz0vFbH8MZiLnuWMm4frzco5Y/azSAI5yD3ipB5dvkfp2Rtp0rb0ng
yFl9qc6PFbkiQHnRvyFeAcg6HyDUIv1oakuOUIphI7wC40FjFTi0T8bgB0og3xZKypwHM+iKeE/R
dkoO8LumL2kuYdWgeeT65Qt9hucT6suVJIreQCTUCQrlrr5Tm4yYMCEXIbnaZXN+nis4dLjVi0Z8
hKSHLmIZvcQeAynC+c157Z9mDSnBKXYy0S4xoh8DwOnjYZpQhOotDAzQsZKF9NaadHi4oMKPiWym
yz2jYjyDF0kQvaYo/bVD2Vl+rP0I7ABNbNTPux0VRANM8UEeUYs4K45QrKVqWkv7wUji2OtUPqUS
0aalQLJjwymp6CXLSRh/uleLY7Cr70Y8YN77/62TPGZ84irLAAKcoSthEqfxAwSo0tk8lmm5iXu3
dVLbqrkpNnr548DAU3tJ0K8h+tFmccPniSgti+rsPGwEqHDHlhLqtCiaITt2duo7Xtc6jO9gpYYA
ATUsnrndx42kYbo3oGpWQXci5YGlRV9K+VlHgmGuhs0547uUpk5a8ffadyolchb2xPc9GjkI7fc0
RVeCtsbT8s+OanhDloTuUuyUDWG2d+Xdv8McYaIJ7LvGEOdmdX3o+5GlAi0Y7s48eAR4Dv0kmrnV
erspECREm13s2kB/SbjIxCIqJVyIXa6F1+/1wZ0Zew9FOuFebiHbwRUMb7quRdW249bvt11DDHTi
VQJLHAUdOiPEa4ThB8sfky/QRZ9hsLZbG4slVlQErAoxaF7U/D6pf0LSgDDKVVYP007ZmLGxP8SU
ipaHXCMPMU+3mGenNqBA8MMXBmutb1V6I7hnFq0POUUa2LHHSua3QiN1ytxOjlttil+j9p7WB9Em
ejogoHKNc8bAyAzrfNd4qL6BGfmC5JvFo79fU8AEJHNYnzYfPTXTQ7vOvzBE6hJ2IvjzY8bQ/Ic0
ZWbql+EUgzK+w1SH3R1R3qchwghfBfd67ziwyevl4+lfxSxibcsqV/pa/jxwc2xkvRObR+8LAM2L
5xwXB2R6dSv9s0VlzemlTXwFm6y+ByvUMsF7UaBKi8aej68zIVO0vN4TiRyBah66txI8aY8yDbzs
wmzS8mkc/hXArLVMuAwsSY5kqQvYDFevYq2QOBtnGYuoe1VgfR3YlbOtQlDIUh1JqBfEmtl3065n
rXz3afnO3qj/Cj7BCetW8iQxUBt427Q/pswBmAL95bNFbXg14+m3ijp2iCFA9HO48X6UrgzI+pyY
RELbEvgdb8LrQ5GCpWCVjfTTbIQ0JHrDwXklFIEZyuhu1hXWF/Yx2DaDPOMWQsCwIJ4V7jXEFmZC
tENcw6+LX2d8ua6K1xccI+kXQG0hnbveA5mVmZokthtyQgo0uFJjP3MaZ/guzO3baojuW2cmGxmZ
L3ewYX72xNtOkPyEVLWA57ftsZLjn1BCisPo7pQRwDhy3zU6lbBdWU36F/c7CbXYToTOpW/pOjuZ
Kf4/lGUEtveQEAdfKPcar3yLY/yr5R/B1W5utlegcWfjX+WjgknhCWpgavdBLQ/YwsICWZlxi9rz
P1rmy6DGAAtqlM+demeC3JvqUEaXRRC8Lfnrafm+VtaqV9nlFnALzoQ6llnuPtk+FkRKCWfQjA+O
gthUDDF6i5A0zZrCtECcm9fYe1l0PNi/Up42EB0P5DEv6tS96cWu6Q55F2MRUturVbbClQem6uYr
yTHwqVRSUYSU0yyUVkYUUzP/v/Tjyaz7OokuRC5R37hpXXeObJugBU6Pa0umJ8AXhMm1aaiqFXZX
mL7yVBspJIoD2a9t+CzO2tGxtBtdRT4Age6b5qQ9qqI8KN5vVGFh1b+LiYYTjkNkbBt5EfF/Dmc1
0VaMrUygvioMbT+kJB1TBBq4eeoO0BdDGE/f2MluqCzgQ90dOab3vRFOgLNrpGePFtvuCvZruO0J
wy1hDWWDSZasv8Lo9zvXCmJQXyQnSf1DJI1W7JEpbYcZoVkHiDEifdbmrxvwlQtZ5PaMhtGTllSF
/ab8sMc7BaTiSrB5if4sf5ER9yYPCiDQaKG8rkKmz9Uxu7XsojtKUBLq7pzBeXNGFTjB8HJwOG5/
uUOS1bpR8ks5iHn7meY2sDtmNJj3RLfuGooxXO+XR67KeQlh9txZwgLml0+TwwOQqI2D5t9i4twX
J0aLrVAd0G75Cz6KebAZ/9+ObK9qu52Ykox6cAeYuZDsmX2aPcuSrLustHIAIH5hWj8YLSaeuA0J
ykER4vgdv4q8m3bJ25CvC1iR82nAcKOsnwbeyfNY2Af5EL4Nf14k0h1K2taxbpxp/0brU+ZPZudc
IBHgov+OhHppzsae0AdalMHAvlcFUxu/Qvby7+KRGBVMIGu9h/CSxmLo0jhdu05BLcPOEnJ3LY2h
VSBAe9qOSRuxVlWz+TCd/6WRuHbmKKK9WylwdzIYuQwZZT0ZgYipRxoMnKSI9Rul4lI+7AYEh0rh
btmB/bNpXOKwtuzH9FEhFH/tYOxNCx10M5w6cteW65Et0Mdhffx//Us+RotfLaDW4ASb6UBrgXQp
oMIvOzq1Sy4ih1KejqrfDp+8GtFCw/8YXbee03mK9pHPQW6YHGklWFzG/IQ1+oHbcEWCUDKdxzJX
18WhDIQ1l1CEsaf2gCu1c9KwZTt2qcgWw2PkjBytZ6RhwGyGl/Pe+lxnyjU14P8ipdVRYkSpHEJF
nAu7uSb8uUPTFKdedOxtcSKQHu1FA6bxVKqO3/lgSnMQMe61lK9SD1MaRgM6vf0au5n79LVyd+Te
7JFCH39a29v3aUJteqn/z/Naie4nZFWMjnmC1WPcfEAl11jNiIjqErgd1NumD+T0xXWmw4snvxGe
LmfD+Hl1o4+PSfwqORaewJVzU9ZhhBeNzJ4MiQu/kz1sh9EtGAt2UDPXk1NAOtlghznypZXbLpYo
dUIgQtuquPDgHWOOksygKQksbrJwZzpZkRGwYzZ2MrXd0rRi5fr4ixj5P69R389AyXoKlzgqWfJn
x1TcQYLQqaot7yEARc8bUHgygrMfsrkgQrRzcDnoM4UbdhBZveb4D7sJ2HyjaQ6d+Hz0bpk/WzbS
yxGQswgY8gKyYSz8JnswKwupievZr/4XDz/vLJ7zYCF5ImSAClQNkoXN5WMc5/HUVGqLuZSTB7Te
tTGgrZGNF5PJRra83udpuOwrh2C/gUE7BkE+4VUAtKCj+Be8vlF6h6vjod+xJSZS684u9vDdVLuM
22g2srd+7iSQ8DXPQxJ777R263sPE2M1ftFKNFerNIeSLRfhrgk0tyyJwY8HRtI97nhIdR2ZjAR/
tnP8PaCtksb+T0vGS38dlW0OqzQf3coGWbRaRGvX+IpbgzN/7dqAWRq+dFtgJkDJ0CjjZ1PgPkuL
5/OeYDHEVpXTlhWuY7P6to7hsue/8gvnoa3tBPFKiHwMN0J5jrLceLvtnpiebayZzxkH+q0bSd04
I0pAwtzruSX2noJwyyhsB9k3BoVNQsLmA97Pny6zH9+2rghdY8Va7F/Yl3HlMTh8Xst2xgo64LUn
am6/IJa1aV4XkliGLns6Hs4pfiyVqYERYLGFZ9I5nXzkMfXDgIUZ8Tw8WWtKOBRC5bVtYuGQk7qO
q6NH9y7cdliXNycgyWz2GOlrNj/57StzQ4ZbCdWjBmk9roDUsT+HUALLoMXKlrWqALZGAm4oR6xX
CT9ztDISpHrRfYf2GRMqakEzXZS5TWvQcjUuZR9OjIfkAa2ZXjlukSW8n680OnKrhELEZx/zc65e
yB6gfx+BSa5wXVhYo5xRRDOZJyLXHecsytqyQmi8cPx161C1G9PhjLLEMVv5Z4u2PiXa/pXbxcK6
rU/zH5q0jcltCcBu6H89bSHFc2z2A7Q4Vd0q+c10yMiXQ17qP2MT6nilcUncaK3DzozS8ibtx0Ns
8ypYbORaPPL6EjG+y7l41JPz0GBmwD/6248SjPtIpUakrhkMuYhf9FGXYW7GuIn4GfCoILJuQKKe
WXgryJ/THZ+FmVRG9saHGu80y30w4t0on0lzvPDDojk+EYGWyQqRcY2ntILibVYe/LROHZl7diUH
6wOBPYoQ0AF6eR1ue6mPbytCsJR91PIl7fus6vRJvwubdtlibnieBEXWR+3nVCs+1WycLp2EzgSi
iNGUzgwwBc574deMS7Tt2RXrSY6SCYbwOsJlevjI1dG1+Flra81VnzV0VOc/Lbwy8GBVJlB1kutn
Ti6OP48MaQzRoPbuMhkUl85Op/h12WJIXv6s2B+BG+YIHve/wAhRT/Cl0EBuEZ1nVBEWzILSEL8P
M0kpACZaLKGXuySoX8Z2VJ3FvJz0crCT014/z2H6q+E9jHSI/gWgaehRIj/pkHg+kedi1IvbPoT0
Wl3llEZnihY4RCaUEpJJkQ/xZVDCnDGzBjOzjtptd9S5nzvntSYinw38Hk0JOSklGYaFvBJgqnd/
1JNz/Zh/2vNPn2W6Z/wrAnrveYUJV8TQIBv2YbYyECdt6Yk/9WICVIB7sqKHgJozrAX1qp5t9jsk
0j5IUjM0jlOXz2veGjnMx+VKqiLhK+CKCok8c6N+yBMa6pY8kDRLuwSdTB+m6EISUrDmMO6IQd+o
xmgiEtYk1u0ZHieD05r6QGWtUekYQq8C/6Kqrcs/uR1xw4eZNWOuvkstNHgFaAbNPAayxcXex2h4
5wXAOeFgKeUPfFZ+IJOKI1n3YEUbYveJpnNcUsBX+QZbSdot8Jp+1s/PHauVcY6VNxRPLumA6HbK
8S7W+SO8XmZ60aLpXpxkWBok3EpZv/YdvAwUMpb9Mg2hb7yCW0Ev6baseQIt7HkcDSsRl6hr4YuS
ACs5cB7M96VaTFSIWVE3nvcfgGROiTwIR9IBWW7fF27IpLB0Wg0pRiaR7SQPx1WwreYBZkAep2v0
DPZZjcLobx+LtfM475bBt4xudNxgOEf28lz+Rxg/7fVTsDsfdIqTZYmNRagCSWZ1GlfJRDNFdJqg
i8lOKsHMcYWz2Ikc4AVcwezwYOl4SXwQrwb4ruf/C3PyckygLovw2+m3/r9VDTC0CJXumMMPXCnI
ZcEviG/a/63mZgDl7/67d+4sO34iIjDgbbeK1fPwjaLBBBX9umdLtoto6n6dGDzE3vZxy+1RBMR6
gBIWT0uMdiR9VtyTuocCNNMAXoFXgq11aedAuTFNEmWs4nu/lHWbQBstsEN8LUKRDpoxrS2EGcIe
CB7yaAlaOf7uSN+euIQMk791kcSTCp4A8raZgF4NVP7cPN/u1DKddvHjyz5nzg/bJE6NTB5qSE8T
KyAuMHTBY2SB0WwSTALwkSLRLWuhFutofbe6WO46QgwW2gF97QLVYmIHaOwRma/NHTVFdbqsQ8ys
rZgMCOUNsaNtagpZDQ7N4nexndu+j32kHOK2Ex/AQQyPbu4dHpgd+cghttl8fGr/TgnDWIBtgcDU
z+08Dkooyz0i5L+6YQJIFgEF5ypvw5Aby4eKq/TyGaUA/qO2xsf+qkVPtzpra8mzKsYUmKoOmzRs
onwwTrRur8F8HN6g/VQsRjaaoR74SiBfH/FCrr6QmNaMDI60z9bc5LKPC20+0IcX6087vA2DICYD
lUthhdOPYBAeEkyqhfXlCQ1/NKgsPHHO+XmTnLHbmuXyKnnrBh2ooYsQaFDvj90HOaZ/vPUIygCR
R6yz4WSqrWtvLUGmmuBTCwzhOYglss8LsiBuVtLN4NcdZ+SfbVdAhST6Tj4YRsvy54fFGONskLIZ
j9jLcmTGj1ZIoEMDOMyCiCEECD8/7JfkseiichRhWjtk3LkAiyP0c+yGajBqxUfmugxNUdrX/mzh
pWiGRr9i0SO3Ld44N7V/zBNykpbN48ycIwTr4NnSu1Mj1pSb2ahPhI35bKR7elqPrPWJLLsi8FX3
ja5CcJPc5MOWNRgmCC41LABRUk2AgL/QP88NDqFL7kFWZ7G4ahkZspiQU2JYx7I/bL1LOkthqXH1
7fYCWRp7R2iqLn5bKbA0z3m7UV8tCZ3bBEe9ZCXkTVt5Xz1FQjWgzDCxNYFNUWQ0U18HOGGofsDH
1gJCMNf6stOs0YriR+spMv/cTI3lfnyonG3bKCveUtp5ox+OD1y0Iy177YCozmb9uA/46uqa9WvA
eAnz/wXpmfRjpGFNbas1gfgwmXxa1bfOSrwY5Mi0tECm8kRRzEiX1p/LaBya/GbjDJOiZdIqJadD
dTAjbVlq9eGExKHjFkE5Yi2O5wegtlUikzBO/lrSlL6qDI9BMQ9oVcodSNFfo0H2AHDNmEwm+tl1
o9HaPfF5twassa5Nvfq6f7ID9v9TbphHhPvldeBPeWRwBsPp1SrGeH0RwWLgTIRUeN7pGpOkTYCV
cStB3PPmPoUM2zAxOueBNZ/Ej2mqtEM8M05krNyhYLrGTftBEIiTs/yhV+QzjC5/nNujixXP/30p
b6oUJ/Hcek2y8GyF+cETM0I4rMOYKwwOXG5TdWnsPkmoFTlZp9ymYvfTeoqbcYqRG8tGi/cLDeKE
zX92tXTLBoNa7tJIbNJjEABrfGaT9Du7T9kXr2LtPEbMp17p7OCvBuC91XOxbofYd4ShhlRoxZH0
227UJzl5HPCbx+qDpFMD2iyktLSzhS5ZOcFn6yiicYd53DIai3M8lmzZujoIV2ehKSGlbV/a5OIb
BDqUz74P+84yM8AmNigEEIAM/4GgTaaZVYWjxAF2k+8neBgGHnKZJ4wiajBcbM+7acFJQ87/wCuW
ktLs/5WczdKJedV9SmXXC+9n72qdRE2MbPjyIBfbJHkL+BY2CiLs/nwI2KQ6U7uRR9d/o9JVxLXp
32SDIyeUM3XmrPTgsnkyzIpFekthZLTdlndySUc1T4BH8HkBC5fI4oa9r+rvXB3C1rN5+3OI7plV
ApCwaTwUR4iNoXrBvgH+EnlQ72Vtrq50vbR9asaWX2rRl9Z5qm5gHx7OvTNyJrTPNIHVYLracsc6
IDG+nY58mqm/+InuUK4XYsFdhbpkiOGmkXEeb+DVTCrX1NplVOJwx5tIl6eNjBjwGljHYaDKedB3
OObRdi/8BsK4wj1Hgs2yTanqPDFfglBDDddJi3OklzxFn2HnQFN8MVzmS6qLkvVZYrr/T1/kY0qj
zZiv44EqanEtwumr0igMeb6TWwkEQohJ7b2lYBKDH5UH4erlfaB0c531JctUMgOSSAotm4Tw4R0d
FTOUfz2kVuEFOkcAjK0PEHNVPAL53N5daUQv6veyoNLA7CTh67uTiXvZLdO89Vod71iS1etm+K7o
eQAb0Msoh0eUTBVvQkL2OO2F9P9u0iOLCG9IxEq48pdFCvV2wP5nv/4guaTb+wMkgbb2kGygM9Jn
dvnWzk42L8wuqHz1F2pZwcY7HVwXLTyoFlrGm/2LL5egzVBFBg/FzgM+SCoWMhlWgKF2rLMRKALN
vw0QoM4tRI+krMA8dmkmNdNYpfcBemXi1D8+UQDrJVubYgdxj7T/xRMjxdGUzPWPIGulvK+s/cpa
SWtXZ0SGivSBrKolZi3Nvwit2kEtsEuTMOu56yLCh6X61+3EIRiRMqY005a4HBGqZALtM4BhCLWn
387lK+NdQ/cPQgLNZiZINr9k8IToL2Fe4RKYVPEfK2JEAzCt7IP/FavPAGBTzvSLw8qEP1Qg0PX3
R5j+N+6aITfIG/BmYGCuznDju+QanUXPM8Cl9yWFeuVvk6xwV1UOrjmXRzfqDG/jVIJOe44Jri6D
e5mjUbX+YAu8YaibqLaAKBWfxLmCpPe3BdauUuUjMZXIK5JSltkWUFwojOUpsqTOevIjXu2Vm0AN
NteHKloyR+Otafn6swZmwdY9LkRNvSYY4M3wKuWzEHdz3XbcXCZtkc0SyBj2fb5NGRTgOPyISvrC
rwrIknJ4U6n2PQtbfvMcfqlONgDJdqX6Df0enFBcTPqmmu9fcUW2uHFq56KzeT/4+YoRPQQvGTMQ
9lPbcQEiEX3xCHZK32DFZKzVJSx3xuhOcekjpmz1lc9Ryed3Y42SfZhLI4oBXFBCxQunOwdTzCjq
eP6vAohKBnL2EeoZPJSTa24/etx6rmCfLIyfULU5E/BcG425y48qoqCkxSvWiNAymIoLN692plWd
tUo0RntRol6U71mS9v/Pom0qAixVAPYPfaQGhSLLknEUGwb2y/3+ulNUsksZLuZSrrlEa3bdfUX5
yBHQIkGzUHyjxlQ4Jf7/MwxaeK6kMxG6x8LDAqFL2CmqPmZM98viP6pHnvP3bFEVQwigCtfWbLtk
t3pzXu+dovultqYk9xe+XqlEotc9TF1dP5EXBgNLQ0zp9dVDWV4TvIAJDfDkJZydQN0gq2XDMs80
bb6CkJBldYGyuLEG4yWDhkJzo+y6maz6S8V59YS94mJLygDwkW1bce99C8qQpfIY7Ywc6eRK7abw
hO1tGgSxtUEMnPAcKYzvVFFD3+sz9qk4a0QqxHr9EEKoCh6Vmv57uI/7zkyuW+IztGWQZFOZeyEv
WKvsTq48RF9jXp37EyqzZHcYmbzmR6LnETnk4diuMSpcmNhpj25UwEY+4uMFYB6YPWVn1izvG3aE
v3NBVswayWanNzT+3vs79NdhCjHom4b6qXCAAcGr0hTZQsolyfUrMgEOrDe0EihOnjIryOG3QBO0
OM2UKLzraJVVrxOKh42B9n70FI6ixHjZsoL+pbKzztU3zh9GitM0x5DmWz4MA+C0vhse9UqL/bzT
0R7uA1YaY5cf1otxB42DQZHXOMiz6pU70kYunDmWcbvcD0URSBAWWCF7OSqoxe0j0lkW6V5oIAIw
oMiGsLU+MBYlDdmSuOf974qPaWHwicFHilJwGZiXIfIXJAktGYMkbvWhqJC95AbSiuxPGi3Pe2Bg
DyPxo04ChVU2BSBG88eUoviV8MmWHDwh7wwV4gUZitbhpplkdySPZ2DmpUdpO8VikWEQynEdBMS+
FDmvBQ0I472jcyXOndw7nMzxTHHDaLuRcWRQDkOBTLYGc2NuTaQFiyD6XZ0jvPMYvcHaQka8kvL+
4KU6zmydqgMcqEtM6+DS6wQEghzraHIgr6IeQmZkY/XFEYclQ5yBDBkd+KhGkD6RCBfoaNKrjWwR
CXmkrw5+suNVMZcoWQlZQRPUwsuMbL8xh9gXHdAO5p2OzISAJfdFZdeMwibFGxGEGIwkRhSahW0M
fUHMO4xePvP8RLTva+Y7njwrTN4kgh69v0iU2LfODD7atNOOPZbVIF6MxdnZ2fcQxOtLRy95HWaO
NjLV+09yVgjA/N07jrOeNDivJOrCnf6pT37aDGY1ITqToo+g8vZdof4/+jO4AhBG9PtqZcV8HXGu
bf0V3BVTnmYnGXBM+r5C5Wf1p7m+atd3UbR5mdk+Z9aW17KkO/QYg3tEAzhcEip/YLr24KdY60kZ
CflsjSOX8DnCgeLnHcde7oc+12amIBPAW7hLrYISO7WYKRpZCqTEat/CjLQuBw/IO7kDOopfeuEi
QzmGviQK9u75GNdVSASAF9TIRqntCRGLsu2R5obQ0p8MlplqWiOgBWdAmLoEbzasVi0vmzsJicuS
zLhckYRXDGew+lmrZ0w0Zlq0/2ebcz4E+8sBzZwSv1iRVAZjMg6TPbiGJkU5OAlXaP+fM3xYY0fu
KRWITKQaNHhqHcKATFOBDd3RT/EzcNCOyhTPnQL2Wj2BwIuJJ2HRKV06tCCId/HCyp+s9zveUmxp
ehuDeCFsWURhpDLviZKriC1bYvL1dGW01Ud1H/QL2juYDXRCcch34SM0YhOurV8VlCvQbl5/n1gG
3iSQkzWDlx5ZshXApdIOP9fqhZ0TsBu86hUuhEB4xgDmQTkom1TxZq4tFFmA3/7oIN+h3bL9YVdk
d2s8x0Ev/S6i8o6OzYwn3fXWKyCRzdbeeGuUlxVw9LQW1o2CBLQeOgNOHa9sSa4Z1oMYyGhdSczj
X+lnn4f6C3ME8OG4XWr4qYc4Q2AQOyIbN2xwAYyj1lue14OhUTbfPCL+kkjylB53xph51/HUcWg9
arDr1NsG88Ce9X+k3y2b/j+MzTLMSdXzxdOmG56OkxPIzp4m86zMn+ylNu80KSVugwRY/9Fc5a6/
1VU+NScHtOg4okjCOYtrc2grmhvS0xWtblVQLezQzVsJxla2qzYkZTsOmDuTlbf75SOpXl9p//sL
i23nhVcWk3deh4OssbOTPBpMzlrHzpRZnUILWIDa6ycEZNe1HoZZQWRPS0Rk8y/uj4q0jbQ1tM+J
8F41RyxccvdWx4LaMRFwyQ+ivWFnrn8CK7JP8Jv3QtPR2fgcaPiKAMMrE/4iFZSqzvDiyFsdsfo3
tYwX9i+9x2rJjUB5rfitkxdo/IvLp8BbQweb99QDxfy4A43TANzGJHfnSZMYEMYX9T8Td73Kj+i9
coxTDCb5z22Yl2eNngB5n0DYsNyMoXl1c8N6oBLctgSPFMSPOuquFwO1nfdRiwST+0OymrHG4fhy
ro8zzOhwy+qmWEmec90Vxn4KEGGQY6hgzeVAqAkmHevMU5eqv0XudxXtWmQWSbj92e14fNznme+H
opcL7RhrPSaQPMLk+D9RdrYWMTscMzov3cC6YywdfsZ6LseiTpGcw9XDt82P4u5n/Hnn3KdtlQ5Y
WT8XG2WQ/Sv6ho9zrD/+KqXHCtnI19Vzbop2hX12l240qp4gswU/9sSt5QQjDlpbUxefpMlPQ28e
5IrCBZCvAtCtzRr/Zesz6NS5cu4VScZg+uamZgypTNO/fFmLfE1kbZY0vGJ9bCU0sjVrf0rHwnKl
ngI4ELz57dT4m542d95qmcH2VrQmZDFxPXeYtD0XIkKi54EghrPVuHXEmxDcPundkZTp9OKsxJxW
GSyGV97drDtWeH1/rGNoKgqng3FhIGXqNSL/leDVzsAsySNUgA3IAQ2G6flKo6huY1oCeIkDGuwc
tsdMOZXYV8z/sjNQ8LTi+izVtXbOuB7UFcVq1I+IleThOWZdzP9wP5d/9TZbCiYRctQezXS6kiwS
oGXTHMk03c2TMYkeZXd8yOJ30+ExzNft4bYW48mX/ud4RhWiJMv6juXsKIsjtZ3zDXqSSdwuybO1
JC+KKFWFVs0delRo8KscQChY9qnOVyifUj6tzC0C7dvJ1Ix3Cqaa6mX4ZY9y6i/mtXPWh/6tnf2/
EdOL3WOQ3G6lsIaGiblxs3eXw8dv08ntI6yNJy4Pw3c5VMHQkdheYOHRvWKQF8dh3da8pSZM46sq
66WfkMWRLBi1UOlDaoggnyfLXk1loNM09mZdK9xeORINq4RlcVRs2CIxzliO11tqBAaB+IKTSyaO
Q3av1Q5B0KqquP4rBngc5vizEm4GlTXYo3JjQxU7OgBtzPLeq3/cxA1TheZB+CqXD49x8gE1Bj6B
slZgJPIazRrNJ5jqhA5E+TNDebFCGiZmy7lhNA9i+9OBOb4j5qEsZbV18FH39vhZ6k6iBOIniZlN
IXbh2tjDznYlPq5hPjwNMneH7sX33+if/6bv1e/l6v/6pPlFQFxTsBjKRPQda/DqXk/PXdzO6BaD
Ng/vMzh1Qqx7OiahZj95xRpO87ET+hXpaNT2wHdj8iBO9IFJOaNtS4YcqH8sCOS/XRuWKp0WcO1i
6l8LCfnkrhG9ojp3s3bMTHaOPjes47ymWwTJw7bRaWRA+yQ8n05pxU0bL5GU/DmagZW3DZUK5tvq
PbzSO2YseZLfoOzRKZRcqXEpHw84dBwbDgiGrBc07toidYGcRWt/p8VPb5668ZK550WgelucFCKQ
7HqP3jpduVqftBNQmQwAHZvSWrye9PF1C6+MUUHtWnAgupmiCjG1MCpJARFQpLdgZyDwOr/5HqNH
2WTD9Q7v4Fjgg2CjHwGNamvosJzzqR1A0UZK4tnLPzfjfkmWA9tUS73CDQ6v91v1L7/+gaGnvzN4
AJok7NUbtfVgerWZDdfqaj1Xu5L1j4PdiH9dXWEViaDkOAf9xSxbH2PyaWNNrOc28lg9J9XgZ7ia
TbO9E9c1mooQpCidfay1b+MhPHL/N1QBBIPpWweJuTfn5MjLakZldHM3j4dKrg7WlL69mjs900zJ
Njfn5hSZrMLDgkAZ8feddeLL9z6Z18UX4fvCy71a3DxcC3H8sjEw8B1iaReqtyrLYN4jIe2K8pNL
+P3j67jyiCw0Dt0eXF1GR1hb/yzVo5QO7AKk8bOf43FLjykuM/MvOVBrNvXEXxal2Ys7Ea7z3Qzt
Fa+mo1fbaEpQ1xkkaHuZtQyr1mHbzsILKgf9HYTS0Nae7vw9hP06t/PLP7nTuhK6zoc/ceEAznEk
CYKrECXTcQXzmfM6yUo3Zm9ldqajWv3IvPTCeT7Rmqp1SSSVCnisdSSv5oGBRUop9BMD3lvnirjE
xjVHZ41oBkGIJ+q35WGlhpCy5U9CaWyo+qNS2ZgnTUid4cWpXejED93wwZDFFHeZl78az291IlS5
buDMYbitShIh3KWQJZPcH9zxrHs65T6iH81cmd0xCmtPb6CpANiQDwlj2LCPnGMZqwJ9lmkvEFO1
WhMVZf61HMHS1S8L5ZpUIqx+A2CcuNm2vX685JVluhi+1S5eSexexMC+dKrIw6ojv6sx21bWbiaa
1R4W1UPsDuy2d94sS8rFDbgrxuCpN5tYiF5oVb4v8EnJFVKqx+EmrBgK3tXgKyjvnvW0r4zvhDyb
2gSnK00k+OOV9gPlOromsGanDJvXeUK+/Qad0Ra93/rsacyOSKQnmfh455HN5VYkcTOkNY9TKLF1
Lb5VDo5n4gnA/4DfIcnrRyFD8USdQ6Iur/81xQHZlbwSMsas/rKlcjY07U5A7bF3t932yHpCVFla
QhuQP8Yultxa+9FSCoHfgaV+o5zplnlJ/6wuLCSTpFs7lhOY668pKc0fVzb3uYx5W2mK39R2veHU
OeHLzXrIgGm3XtVWR3xipyFc5WHpbkWeVJGhWHukg5WY4u5b+LBywyAK/A0PuV0XU+SMKyGUBl+k
47OLCEuM8DcQSPLtd7OxVU/U49JTblokxTevcIIEkuC5w06KjaZfx0z1YDq+9Zv19TrRsxdXkdDm
44dNdtBDn/mBf3/1cOSJX4mi+QOr1t8KjbkatOnvAF/+z33nBIrsvyM54MEtvTjjuHexCDlZk28x
IS3hNGEaCJPbKHDeDlfbL99j9/AOcHbT+57g71Azyloc0Yj7C6EmOdpN6vI3pGbBrbWtcVc2+Uu2
YZ2yWgfEy4QaT3Zt9IloDfFMhPmYCXVA7n3YkrNuEG/Vq+fddsFbSs4HTKr5jfnitxW1avRpBmQE
QuFzVKh1kgnuuZ1pcY6PO4qTxVv5zy09J1JTIAwngReEpDFFRy298cXhVF5WKNf87XuOo7MNky5s
u0dZmP0uXTHM10KCEhscryi0/aTOADmyH73jQnigOzSILQrWqR+ewZYNE34+4RqM7Haqnux760zB
PoxGyX72F/g4iLq2ZPOh5uNSTvUDAnbof3j7O7Z/VN82zVV1lPnVA+9OBieN7r0SdTzJpcSZ84h4
+2x3ZRjK8XmUSfbf5K7MgKGqv75kMSxn6aulnq8hAMtK1YMziIoXBckqEw+rmOfIXp3CS5rTHy+G
0Pl1Ul50v6AYDKD5QD/OKOAcn/MuTTDiBL/+EmDYfQ/VKef12muYjPQw7XcaMaEa3+RdHIaOs91+
rHuHU2DgzVdlEDOE3ClAxFNsdWWVbHLUSobVeBzs0q5UBvuRxrDjcYtQbBvrLMi7OT1zduPVbe9H
YqAP52tv3ehXEIJbexbjs3OM8cBM1hcBU8cv/w7Ri0IBA64B2KaA8jCq+dEd8Q1pzZUjtpqQHT2f
+uocVPrgcZPWBXvG4B7QBsZxmQW3mvfW3wx4rCkubjwAyALGZUv3f6Mz+fg8U/uDZpBNpQaqbhzE
ACRq1q1ULwqI8TsawX1aCdebUA4fSwrEiiED4pbJkkFjvS8YkFPmKbU2puLSrQAKLVKQm/3HT0+I
YL8dbgwMocq+fD3hvVlEU/9u/Hz1OvFrFKzPgmHUVWRJ5HJ2iv9YsGotgqVsqZLIZ9BVU79J1IyI
X1m+3tBZkbCc5V/SToZrEPxJCq2dZ5LUBmOc0L75WvXL9XMStrMh3exKswKTaSl/MsYx/lrdnUuJ
yvZFdUYL0c60SR0WDBSD/ToFPPLLuvM8GgGc95zKjNJa2D4tkyra5jLEivDRtZgz9Vt4YyXLy7cE
PGDp/tkHLl4F5dyv6a7n0gTEDyp1p3fejAoeS/3sB/boMuk3qnDU6M+VfG1eI5nrjd4OPz1G+sJP
B+LJswOD+PI/ScaZ+Y8QqABKh9u3CZUL5mMkGEkqPekA31xxDn3OdtDSbDPkD9uDY9aloKvwJlQ2
Dos+UdJZoKDCpcm2MiiTJ6aWRxauRZGX/Nsqan8C40BkpEwN+sssq0CBXVKYh6rHEBY0pL/1gA+V
03iTvs2zeR/1ke+R0XicDnJVXBWYs4vatn3TGmgCRstoyh3jshCUQdcbaaTXhuWI7eAnb77kG/Ri
dka16UHMa8Pi0Qg8+bzi9psDQVd/x5UnSjn3UD5oOajxGuBiSYnLie2iR2YXJJYcKbniGXWumLv9
7DPxOOkZ+lbPFnd/nsz1ixd+dxxkUBfK4u6e6Ht+Vy19pSqkspwwz4HPKOyfqpawAjlRu9GeTDzl
AgDlfru2HRz2TCno/uSIzm49GXBoxMendXPck4ttaDneBgkkoAiUBBGPjpsbXrstgKpyCoE4WoOq
k2JUaj7FkBqk/PNJRqjpfNJT9/ujMuXGvrLaQRaHbtQtxNP+oVKiVzQOGyu1QvbzRt3ZtpAnecM9
JVa1sV728po9vaTq5kPaxPDBkhuyhv/8ZHcL0n/N4tYd4fISk3yP5cJhVHUsq/mY6w5jcziqp04b
tIK57fwCkcWfB3txL+p00YMO6XSaikFhIVlkITm3ScfKT2jGEKm+f1l5NMLRCZUyDUATNQn1nsRs
45gFDpKXqGLLWVt15jTFheWAJH/3yFbZqAawcfwhd4QfXXv+I13Uj0ujxWaf9ON150T8ullCCVcp
ZzSJ5TuHvohbeOXYDPwof3AgVpscw8F5lxQplSLswem+ln2TnuHhGSmAdsIXZ80Wv5wc9f7R53F5
qyub0NviNaRv6W0oRVXYNVjHvXrZ0uvEUcUUWmvvcEtOH9yM34idK3eR5qbt5X1kJJzoLdAlc8rx
xTbyYoAweb2H2D782s0OytGrR5vIhEZRhqStgo5ydN/T9UdKeOcJB/Ky8niztGkIMDtrOg/dzSGi
C9Utl+McljddbRd6N89TdtY6k0+WMKsTQLQ1VTbxwYKTrqKXpb4nq3uD1rxzgnNqg5kWFUHqwYlG
60Fr+DTacwvmMXiFg91KcJWgBvATEhynMW7L3c3g5Th4TAhix8uo3fBLF5Bfy6T5q36sYyiVQMAE
a0MWzLzLHjwE9lb5ByYBwEfPTkSrepnb0qSTwTknl/rt/sd/oTX7pc5V1G+2PeJK5qzRc4tnXWbb
ynJyFfNKLv2rQwmZ77XE6CWWdggv0hYKojo6TXeNJaH/LWTd2mgRpIVrJAGrb4tJg8UDbH8n4CPS
sTGN9L7fHrrcm1xJRUHAy5zS6afvd7HLv68cNvk5DlsR99PwyJm9tMOkSLYrZWMBiwvqRMhRXl2x
KzXQQ9lAzGs+OC84uGNswug5K3DL8hnETXaEm6ecX4lOdvxhXEw3c3m+kXTT7f/M2N18il+t88sJ
5yV8YmMGQYPLskO/np/3dwPzsf3CvfeUbij2Clm7wMo2RYpf8YQRCDdA7ZPrr6W7IGDHG6DN8uDJ
TsZ9/GwB1/P9mdKrEXX4LHok04ESlhf97KQ4Ka81kNRoZuFtqncwRRdQc9Tl3zf93u4HT/P7aSKM
kEj5bzHiILlNp9hQ4VurcFETeuz1Xucf3pp4WnbPFpHBD8NgTx5INzyRuyWiUvvq0UgkAGd6M56u
Jhxq0HxdWie1/I9JXlK+0mSo+FC5rwr1kCUZVIquhn5RXJTDvDLsplHYM0JI1Ed9vsDWNf1Uj1MM
fpj/eGAvnu2q52wSXFz7DmHFlkatpY1XZLXNTcPdFfDF8gnKCHupfNI4jNFVolF+ngpVDQQNRafn
pvevSfyk7OH4SeDexz7KoAGm6E1iRoNEosR4WaG9XVp95jMtouq5uPyQzKTnF5Otuv48ekEsIgSy
dE0gK0s9JdYZmhnPRetw5DYQUdEl6j10xXGFmBZ/MQJT6kNKpXzStsuJdNrydIYASkJzijTwUsDx
T/ScHY+1+3LKW3WS3EMc0wkZrQzzNdId4ljtk6Q0EZEZaX9J6HwZxGRatEtW6dW5In48RkFWAZQz
IL/mxPPF4LxZJWDg3RTk3SpxQMt0V+Iil84FH9QG5B8A+RohY5njUn/ldPLvjW1v1HZ9smHJOI1f
TsUjWQG4M4dILVqb50FvdwzLVevCFtAluiUB8nsRmEHwOhqhGxakvhOKzEVcB7j826LGNO2kTpfl
0HrQ6jn3fAMJarykF1LMWGVLFPUGbi4BC8HRdpHiRe1kenyC41KFshzc3TRFZnDL0Jia/skdcsyx
rn6vnr3pvjWW8DhyF4JT05ZJRdH4dOaLNZ9NDI2vaQhtl17aOSvNSogTT0aw9xXlXD2fH74ZCh8q
AnL7KIBu6AB77hOeCzhxAmc/VOGFchhYxd2rrsiFSVjaRno0+IwT29B4SOaoCK+tsQ67viOtZB6U
SnwOhvG+ryoRtjiRhGdlVFpXtctvdI0QaUYwbDgnVFhx+OQ+qipLkesTN6v7XJUKbk5HoZ+0dUKW
8js//Y6+bB4MwGImIVlu9zWof/LuFUQW6+mjsmFu5LDcOgG3BCSU9Dx3v4V/RmrawyCa7aTe2QIb
YE9sjpew9/aWkBt+4eyWdtAUdy94LPElh3cFlJCM8ao2KApYTpJKGXF5HsiEfZJ9Ggs8HXB13Ob5
R0x8IZlUMokmkq5PbyJkJZBO/NOj8tqFquWN9DWH/Tdy/R+O7jl6/av4NnMP2plfC7zupKkKYuLs
OBw4COB/rPWS4T5Z87cAyXwkPvcFAof8dUxulNLE5JY2LR3IGaTAAoBcU+XH1siJDXYaZxkKaA3e
gUTXQxhtjuy4ekP8pw0beoi07/EceOLs5K/lgqLuXX6/mudmaD6GuDCe9tcNgpZqmWz8HNLexo7z
hjIIv9pL8mPa2fXIXrlQM0uvY8p89JAUXn6+OShVQvOwgyWnz99A+2GTvZpXkeIgpDmLB7vrN1vN
JN3D1VH45cTk2f6YWuNNHTzCRL8A1bGXwcFV71fts99vCpPxnLkp7qke+n8BEZxGSU/3ghTOWVvq
imo4rrzgE9FNYckO3EMqHu88axLoRYR0bEgtga3jGcOCFSaid+/secDYH0JZwa2EPmNv0GGMzxW5
mto9y8OjlmP69vbQmGEFtC00GmdrWQmBpnBYkpX1gWJdnLs0ecyxyMuU3m5XLv1ZfjXY7iG9RtS4
RGvR1QNk3Vx4lnF5HKJjdV8BJD59rltsdIvJFl7tpY3GJd6aJ6t1xx18XTY3xyRz2J16mcGC28tt
a60wDTKdMeSZeRegE/E4dvvFLm5RkYOnpR3988WF7IkCpS/vTPE5CA1+vfsUU1cEAOp5C1j16Krs
j5WLZy72wz4B3C/veNWTwL13pQrfE173aporCvUTalZuP/jxsr+HgrkAjA9WfN6F06nscw5brSxZ
P2VWetnoWDfeDVZijrvBXTTHaNR7myXvYdx3MNiN7Ey1knHH+p7d1x2XT0no9k/80RmwQU5L1e6Y
M42z21QEa1NFbvhAkytHg2CIIEU53ZoC/q6H1TQh7fcpjywSrqMykiZ+qfhn1ShftzLPIZQDbyvH
TbHYKV0mX/E+FyoftL+snlJjOwrd7ejGNVoppRO15nfrsYnP0vQfncvYScjHLMzj5uTRpfs+zlEc
3Ln1mW2Jtw/0vqBDzYomqI0pIj7vKWVmmUEJQcnMFg67zrf1ShlbMrBU59dGsD6i3ZNbT+e6bnkr
kidjO6C89GvJHRAR+NHqAqy7BKMFEnyhJ331NHYIDfTofBB0sMuM1NFN0DSxuCBOe3Nwb7EMhGX3
Lw/G2SnWMHtCHOxYf9d1zN72vkZ3q6uBDnM1wvbKYuiuRiZqOEe7RmWUQ4cm41Gx6xyJMHa1iN/H
zrBD4SQ8aHeYwmAc0DoElZBQtjcO0EXMyLF95UkbNmzkk8erBp5a0cr09tMoHSt4RxJ89w78JZu2
w0aBxKATOwtcSWmsFmms3J0MlSDoR9HwAKZOsHBSCaPXezrIgiKGzNkeB5WFepOKNsyvYfnzzSX/
y5P1iByNioGl8a27MvDc7juCb4rnepU6kuIzXBmBf0Q7HfSI8NccHEm2mdLufOUHV9SR4pYhqQ/9
QNvnpr+f7hDUjw3Z8irTULdbcchoXuf53vy+DdwY9T4B6aqTrTqi+TxB8fMDSg7eQvY0Aj8UdixO
sNxFBua1mAEtZKZ+pl9rNu+iyc0ne2fAsEEPJm2n9c+0EwQ09lF32jfLG/kBYlSbM1DMWvg2pINK
pP8uM7lPSS5AnNpl3rPAZwzQypYVZ6IQYzs1XPeX728SFLNI/iCI6YQo7XVkn4WwfM3rPVKa6/sf
G0HKqHo9z/zPD14YbKB8+yJsfMyGgom7jfxs6eCWReMd5E84MjibExvcWjw41eChRu7DUPfGnL3h
Q8rSvWi5kRmnIe9U8iIqmXvgcUhfuFC+ny53ZnJdHnWg0gQvbWrIxC79j3QHAoVhj/D0N0t4oD/e
gTjdB4g79+64wwoTyA3U86Zk3sx19EcVEjc1vCAAesoI8/Gs419zFq6kP+fLc0SLAuxyY2TU6qjh
4cRFg8scfU+52yJAaj3EhUZS03DuF01WtNvsuLTgMZuV2mCD/Kq3JJ0y2p+ZApKnGboeWru27cUF
soyKYW+g2ywSSaQrdZJvr/yr4Fq2ETQF9GaL8hIiGua5B1SQSiNr9RNfZ46tyo5KSvVl3cbm9U7h
wJWA5GY3yUmZFtFMwQBDMdyv8rWiAqsFdo3fx4lXMTXoD0KVD6LGp0K0r0M+abWn1VAx2kanKYHH
isWoAuU4cRsXujEXPGDiYK0fsTKAKvKvWJSjAqlwAk03ARSU7ZS44e2KI08SverWegawuqyLvAT8
ECNdoipoaE82jMslRBtO7vyOEPzLVzKI8bR+URjMHUIF89CWcK6+FsCGFRg2NMitHXTsGXeZ8LwP
x9+QFVv+Oc6rCD0XL9r28owto6eScyyfiLluZoSs7v3jO9M2l4llSVZ/GEs5w7YhYQWk1/h5fCLf
JLv3CduVAD5dJTh5+F3kSjM/oGaW7nHIYR5JF/Vl4cuYslGi8Yws5tgoUX2bWpuTkexlHCFFFphr
N7omGvYBxc7BiLDPbr8KhZvS+Y0pRmix2DhwDsUzPvHROVizL4yQBrUCoSMMTtTaasF71U4JmzJt
k25GzCDnGDCa9OMq70KDxxxCnY8GZcDgH7GUO52DQGJWmuiNHiZG8dA9BlVBiuX2L9Bwmlzo2EZi
yehL238wkbzQ+BCfNyS6HFTAILIAzaUcOK+QukEGkXgh4sZrrLbU9Zt8KBa6GGgnDhZZmg/4ZULU
PlBKQSWqHIvlKZ+dKJz3vd2RsHZDe3HdHWJDDIX4FpQJ09k7iskV45vjtPB6Rdlrqb/3Kh3AShBg
9mFrXDrN5+LcijkDEZxaprrYVoGJ91WEpjYthFDFMVpISaUCmpRYJWaCBtfGOmOeSeemaET3+YiF
W8YbD99Tf+hsS5KfnDJWXn6W2Hw4o2gYC90XomucMXXK+IHu3pu2JIcI0kVRtxqdULzYrcfEwFEL
iqFpHKNGmeS8EXTBeGXMUkazWi+LeaKVdK+VH9QSg+QK7m+Z4L/6MGiIePwwFxCf3vIY1DnizTMG
B+NUvY0H7tX4qIVMamybEVy2dUtJ021qFDxtf8yLJ+3ceJs0NtQvFaIIif9vqjaOFYs/GnD0y3Mc
FpjThB0VnUtIV+yNlGU9MenM00A4T+Z+zbmpVXkQfI1C+i9QN8f1Vp0aVYwCE342ksvinsilrq/S
u7/Wp6gQt+/4Mg0e/0rodjifoF1d7GLcR1mpxM8sW5McYK81tUYImey7mkb9HuyX/IkBpnpFJzIm
MPN8LCYwiFhLGSpMt7eXAgMg1R8utGfLj+t4ErsjyMtsPaKIu3pr3m/QCN1XmLftFd/jRdf/VG4n
cWq7GnoLuPFB6w10Sx9QEelsACsjt8egyfkq/Uj+TFzsBzL2fcgCuqWpQVV57d4r8ZSFxGL3KxH0
YYXsUaEXUaSkzgyBYlAPzM+RXwS39MtUE0oLhLcJtcGKVK3iDETyTw8Y7wL066Ks0fGFRiNIjT/H
ERMqQO4U20fsAhmKr+VHMeTiCCEEEeARAqLHZ5rMMsYlYWsKuYyLK8L3NFLeoXp2sIlKEn2QDrfr
mzKDuJrCqQYYsRfOrz155rWxhT6fs18RNw2IMoWq+g8X9P7uU5rJoxumNqdvY5xqojxZdmOAnzbt
LXTNq4jwPl5mqt14egW4ckQiotrmzkeSaWXseaDPfG10lG/3F0Kae5H0idz63/6B88gw8hg0U4mQ
Rwn9VPeZyjNBLuDI2Kk9291+89zWMciaTvvU1OWtRlTY2b5101W4liGXDihwtKBB3GtguA4PU0SE
yDyUhGxhpNRFXE3r7qun047Egcu5qCMbbUnvdraCEMJ6hB5w8AZTSSCWZGcXmXSVbYovul9SiYPK
/0vZcihe1WI6X1E0sIVIkcj8aDEmlPntEHEBmbvyc3z1R2EuDEu+fSNfYWOq22V0HQpiJC4B6deh
77otS3eG7OhbkLdPMZz1aGxH7oyp9PNI84mFNg+oDP+nlU5ZaODGCvKeJjb+C7TgefGGjvXdlnS1
7znhPFGAhstf2GT+rodOtvsFcAsDshzgYxF9ddbpQyMVSEs40h7N+CMMrW6oXohSiyxQz+5btAU6
/Y8vIa93Y9mvD9CF4dJ/mRgtWzzWJkxV+GH9Yqi6yoUvv6QW58Gt7Mfun3xFDR18EPQK9Fd5ccCi
yMuriH4NnWgweQncT+0slJAVbpOuIro/bZC1fUpxq8VijeuLenVGWkfghsvCEFxPs/C/E5SW7BCz
EG6TjJ+KiPUXOOrHcMBzUqlYFfGAUZEgCxd/MUJB2K5WSo54Hg4RCuzeXC8vfAtw355bKZw6dOE6
zXpQRw5srD0/pFNLT3e/QCW8LD5TrJR/AuRXfCAZ6n2UFSi1sDjRNssh/ClTyaG2wOWR6Wqvy1C7
56DdHa58Rw6c52Jt9EWSVd/Ku1izpSlcLF2YbCMOp0IHqEbFrFe2Mx3xsOpXx/BOZQlo5SOVn0Pb
3NiN5QbSWQ5WUyX2CiXezWGLeryt5vfH8RFrNVX35EbMEZ+LNTuKDD2CTflSXLCB0WnhHsVtnvWy
LXjm6lFWHA0UQ7im5V0cZt4DEUdf1IBFvTS9ABjKMI+D+zLVRB4VUxY1bnnmk5MwV/RBWcuDiTdH
TKnQx4wSf0p1btSw6PhrWCvVHdEUWkAgHs8Q7O8Q+hZiz33vXlDsNWYk6kGch6gkyOJdSt5g2zkb
u04jAsRYGwwCgLmzjNMYZFwfznH61NGzRrU9yqV+2Tdkvr3nKJtbhew231YfUVEQ+YAVRX6Z/0b/
eiyn55nVp14ChRXSJ71HeAOWbEnAZLpi3MTfUaCKRGGimjwrPc7qKwCVpmXtkDQSgZrH9CcPfXGp
LCuny+m/ND84PMFM7iuvIHkQseG89fsxU8bJBSO0Lw0qgtR9YyIH+cM6qJhmmZh1Mfjh1MZvjdqZ
ByaS4W9NyYaRzza2XaDts0gJbITOjRbkxchyP9cR1Zvd5CKfFCZpGHMyOp/sVj3pLN4RZM/5rWg9
zWOQ5olRu9WvFPf77OBqdnZxb9oAHEGbDtoJElYgxzjkDOnl+slST+gqvs3RyZNStQH5f6+LjYP8
dpIDTEsIRFAjXvFWr87WSPqHyyYgsMlJlO8BzKTyG5ZT9gyUcIStqTCCFPrYah6mQWUtG9n8pYBP
NQgcAYI1yMJmTP0fDTh+rpfXHBF6rtJg7TTzbTkxg++AHwEl+eLMspHeby6+K5VFyLy17injIOXP
5M18KtBHTFScOxJ8I301O8mx4Mvpem4mLczPVNrNWdkqnX1WKHZR49Lw/iOS0u+poL79ouUdQrB7
U3LeKZm1MD2r5KC5Uc6aOlGaSoNPeSamKh9C/dRZziwhFeQ+z7/wx8JtcFarRonS/gX8PcWCjZeQ
0tqWDWPmZSXBnwGOQgA3CN2rU+fIClcXhFWUjj7PIDgzI0dTD1JJpElxabLeHqKW6Nb4Sq9rvYjx
a6FJ7dEzEU+84JMmQxYKtvwuWzRRcqES60Uh3yc4zjqxMYEi+cPCQpQCqqsICTAsiI2aN4+7h6Rr
p/kZUKXP9/+Kx3DyESO3X2x9isWFymAik2hkhWNk7cRBGCaURNgpbZZ8V+MXlUodU1bqDiFbItuq
fmTV8idDerMEWhbrhXt1P9WLR1+DHwRZqbyoeB1HiK4PRLm2iLXuoRcQRXSWF0YjDNGPA9CBorqw
pr6IUIuDc/2wFESh+0XEi+7mqdOlH5TSjIWmupBcM4+Nx/cBOM2j9WRo1hXhUjYj1+tDrX/NUkMp
52Yx4A7t0YPYNM0AnHgokPM8vsh+WtXLgT6Y54nJYE0xyWtXP79bZlczpGRMyPwiNoQczz4+g+Da
5ubU0aoPurQSVTyVz7ncySnOrAlrb+nm8/GPo9Lf9BKbrZrnWX/mEayACDvwWiBqhTsS0ZOwfO0e
T0UMR94NzOHQhZoaej274SMgaIOdSdsSC+IxnfoIKIigCemw2Jzwc65OkPVcvTVKYCljXQCc8/J/
9dpYg1hJws/EiUO8CA4M+EaLSMsq0GMEq13xpvkZNkvzUIm0gOI61RVgJuHxFIX3DKiMFCr1Rmh7
cSFgDwjUw8Ik8nxHGS0y5zZNLRnNCVJeznInw+FvbrjmrrrGMfF+wrLwC/GeFMs+cWcI9I2LwAdb
bb8Cmj40arYz9Y09DSaSSQPgbiRW10kvPElaBRj0LpADOMgKaEVP7FH2G/vwEunNfZQRg3gIFnlN
dwc/J4gcCQKIZbIOvkyG70aMEbAQyKx4m18zALffRI6iY+nldMVKV/eh3uMI7UV4/T62e+H57Tel
v52mYpOgJRk9uRP/MUYT6PqNVNhVVIQQSdNJFaj/vNt6mjOwm+33P79JDNPS49W7biKcKCd8kEfG
wTok1Ha+87Gn4NG3m0+Y/iYO9asyf8xEV9ruiuggcgu1qzgVjAa+1J3TBOWLDo9kDtDGhUcqIjAk
Kke9epBpIh93wKe6QQ5UACeHyRMDZFEU3TS4+Terky4mYsu+IJ1hX80+5Fj7YIf6QNKM9MEni4B0
C7JsSJJIua58sWetDtieh2oK7gbUS+fSVBjtvNp2rMOlomqhBR//IZRpVeZRUwtVZY8GNn7qAfk1
SGv5BxZXuW5UmcMWdgpF2Vqv9GffyMYan5NN18aICr6W/shjIvdQG1OwmjFQ+W+R4KPEkdTL/pwQ
1bho3dGgVR6jhnUqSpLLEOwZ6cuyYXToLRdTAkN8XMFtEZya7kTdt/G1p4o5PzkeRM2EwTaSiJFh
XWK2vH6M7zmE60A9QMBNjHntTVsdKkONDXzwWv5iV7l3gz+8u14gHnNBorP4Ib6mkFOJi/tL5/9M
G4Di51Zr9IOp/gD5kjisvL5vQLBDmff5xmpk6aaVQNpp4rlZPImUzzG7RMTKQ9RFIsLrl2D9ac4r
GKV/+FsHHHyfpRTeDiaggvXlLqLiLDdsrjywii2weW10ClJNSmzTkKMhkv2+4ANnJGl3Xcq0fLFq
vXh5iKigqqpmQPoq3ikG+EUAFMVBkF5jGeJgWp3itj5K+V76fyJaS077K96IFY5xVTXFK57c55hw
PwB9SAaodhjX+UBKmzHjcWDesT0loFaY6ALbUIejdWWGhqtpL+PGkrf8lxaE6bgWWfF7+RRGykcK
dYk+FeJrW3dIWpF0kYthf9AMWRfxE5k7XtC1qVGGlSob0E0ZL1Cc+1flxKysXI+CywsU2lUsCOLI
+twYJBL+Jsfyrf9ycyUGWp9KkjHmY0Hu86FyVpLsHdEAwKkeE5FF7azGkdiL1bc/pxb9+RexAl77
MTnFS7B8PbNzZjex/mPLpi7oDs6rPuYgAngKYbOUgOoHEpF4670MM9syrWw+w3aJcjMOSlOkO0T9
lAZo38ghiU6IFuIqVXWaxlTKkJMAKHnVQmhJxMnKdi9fz9+gpzYJ+L8uV1dZ/5Y+msFDZ+fddarb
JPog91NbS56BelaWlLpXSd6M/FVZ4iK1JuVyPlqPuZA45f0s7611O+f8Kbth1hT/08yb5AhZ+OKL
rqh9npDcOM30c6gaxua0jtLisHEnoTdPdUcVTCPCq79Vz3Pq8oxZe49knwL9vJr0ncEWesCPhH/7
ChKH+BD51XnbYx7k2QlC03W+LjhtHQ1KCxYZrHcPzAj8YlQMn44jLQp94no0R9JILtriYgdR+1Jn
lzAH9PWoPo89BlDcnLj08SpeT996hk3zP4NOklg2DhZev6yk5KHvVDtgWOkh5MBG4D+j1Uy4EdQU
t30IZRqzjB9ORgA1HowWhCJFVXKzgsfVZRhHWBwGvDlFp2c185f9GKNcO2BZTF5mXylhCor4oM5A
CnEInNZ6M/AT9AXvOkJUv+mXO0N5kYekE0Gy6aIvHKWtvfbjBh1DLVlSs1b8Qd3OqJS6P4cSUIIp
lY7P/SvvBhvqsOxrjBEP1u6zpSGGySQ2LLEG8cE9cU/qiGm40SstDnwo/o17JV83YCdTj4T+ggIf
fEfzVvJEFXD5j9oD47D887pwtAgXvCvtsKzu4CTb11ku6RVKmZBT7ZyopORMNXpmQEdmZtJTiemp
pCVyWvXIKyvMVV2MHGseIpzWAr2ycSF2PcptJ0avx3csjgsQSI/nQ96/p+0iiP9Yck77F+xtl4TQ
lQdSSXiWIXwm57eRlRdC/wjevkoPXCIckZ435erV5poKeZrxHjdUUstrnaWjSv1ruc5gRIbPc2bx
WfXTDNpuSH/Hd0zyKwLS8cMKMylkzrzAJcwnyT+C29DLEC3dnDWJa4FIt9xFCTicreePGXnDcLr/
8R4/A5sPmULmMOe+7PVYMAfFvDU6qBnmD7uEbDzO20RNyXZWU+hk03yAj2GmV0lwxu0ltDxUXXHA
3gOp+AtnW9Ee+DlwsdPsF6y+0xQyTCQUFXsC/NWdIt9e/d5x2jD08L7nkkN0vK/QLpYQl5GDXOzT
CJyCCBgBgcLghb/zcBP1XrwLvYslkBRC0OiOe35JhOyEkP/Vq2wVvvAgPwUN947M0gQhnwydpKQG
nxhk+syaQ5lVkIz0Vy102LZ6RAshkSdr+E/o97ZO2WPZLN9d+45co6+tQ4KPa73FBDQU46WPu4aL
H1Ui4CPg0fpb0fGkKMESZuEYSn2pFikc7NMWvccbpyUc1AvQ+O0QLlnz5fCFF6p0m6gu2+WV9B4R
AQ8D11iIMPd5uwZznqi4SESuz+Kj1w97kmvRbNMJ+XxHQ3rpP5aqn08le62Pi3xCeeZMfs/k7HO9
3AOiOrq4S4kv0RagO3q/peQLnlCF+Ms6ssxdKGBoX80mzZSqe0VCSJ8birsTxK8xmcziv3bmv7GH
dkQczvxjzr0HqKifRuNuNCaZFP7alzG1WhrkIEOd1/Aae0RR89Mle1HgT42w7ejvYoyAB9QQjDlT
qD16CwsIRX33YhfnxJdE7tn5jwFR6I1zn9wbVqnqnGeKtL8vNUe7Xk4xfjF5+ZwHYZLQZ0EhJZbt
1eVaaJLDi1TpweJ6yji0n5ADRmHEY7s+3cv0FIzS6NYSUN9QSJYqaU1A+d80Lc8ayBNDS4cERYBL
ri+cPjb11tQlBoYPGOOfc7B586k9rAXcHgWInh8MyF2mWLTYymcowA3nUDfRWXo6v7bEteRURhoq
3d19T3tkAxnenIFCN+ECPkB4f3Dggt9qWbA9pA1ArP9mOJOriPu19A8sT1C2nZ7XCXukspJOWG5z
xB7sM9yA6VWTOXyHTsB6oHUxe0h2MswGEx1CDq/4iApIXn7/KE9vNhCd+Q8OXJnsiH5gYJAPdKZS
p0hy/NM2iDwM0VrtWRa736aSCoaq8gTfBrirnKOF7XlJfb1dhr0vmMkVOaEg+lHJmBTTzGWKAqP9
VcF0jzGsjdt3Rzn1/bC6Q6vmHH/RaIREGis1r6IoH1DGnVxqS28wkxiL+1a7oH3D9I0ucP/ZV5a2
SEl5pp1Vguzlgi/PLuUeihrUz8a/TZinKgiYwWDmOqXLGn+nvbufduZAu9tLKjqlWgZ1FMbjTjpR
LwIg3AwteT7+oO2SJUiTjH9OQok2BpW19yFECEKvsjU1/CqeAUWPtuBc9FP/U8NSj0Twssi3i6PA
LzDSOBrH8e8zg1aVNWDxo/Nrew7e8hzyFjO0R7+8Iu2hu82DGyISRdZOw/wT7xhMNaThk8nwNa5e
uHbVkP6Teoh0pkWM8jJ4xbYByKLRKC72za+TpDRjS7XJzTq4nLiQDdrdW/WV7t02bwrRgTmcUOn3
XqdUc1PEScB5M2hVkgdw3OVsoGxTbXIT9fZJMdWtlmTerCCNin8ks+hXRM9aZB1qL8Rr3X+EGnub
J1vLr78ZQaPCDjZu7JXD7XkktoZCvA8KiyxT4LAuUq4W32OWelPX5ED8xAsxlooNIDEkBk6aS8eC
EqRKmsUqm3950GP2cTto7JosKVpLYaHVVz0wQePLMWsaDvhr3LWh+PB6keqXWgfUr4KtibIdjpjd
Q/0RKlHZmVjE9ng0ESsFX4frB7Lf1rq9RkXRvMuM+puTS5FlU36F5zz6zlrLKGMM3Qs+8dV2fS6i
N6Zn2rn8KYVO02V5qCv4uYld6amh3oADx5ys7IxgXbRYNxB+pxcIBW+Qb63vQ7HzxYuP/pdChPJ2
8BAC98eGreQokeQPuOpuBDao7xM3L2H2U+D6z9muZd6g8OdQOrA9qFC7z9ZBV+QypGaoRBqcXDiQ
rys2d2CPLylBlJS13qLnJKtY5CZjAdk2yAl/QsI+R2ZBPenuXhsCaO/LbFp+35uychK8DmMxvOF4
YC4aL2UszlzIx3BnxHuOjqH2SgKrpAmlbS7slv4xhsRkxp1iSDC2tJnd5u2JqZ/L2BJlWrGlrv0K
A/BcbCZprufbo2lqI1GJucYsnlEqnQDLsYmwUpc9jXbC1ra9yDjJc+8J0DkHBsJKEwckUDKniKtG
JD4XO20MpQMEa3cwnPLmwfHuZYYZUvLVrKCXoy0ucmJClkwuv2Prx38zAhTVZYg5x+d2s/PvnEf3
nPN7WEwm9USfb/AFjhp648ZXw0qrQv3D6zffxeZQFDDyR0LTC6H2QPdyfcpwgRDwpuL/WskVlJE4
obmMKI9T2GiK+MqipaHRvXDyWHwBgVD0Mez+2cUT5GOOiEQJ+cYlVSxcugVEqs/xtYfxj4tojaR7
SZuE5Ju8zLodapGmrU9T7dQUKtdtX/taL3Imh/Gr5fjI6l247EiEqIyLbHyjeRZcQjWWrcb1Oxhw
Vt5875GZyyhVrfP4mx5aMqz+87iXKwo/LoeeQA3MK+HsdQbqQ+mnLT19qCC5/UDWM4iSYrmoxkeY
qg3aPvtrjRvTGphBwCl/1zCgpcHavaYHC/BCnLVj7DCGlVZO/RvnOsCyaCfm94m7MeY/6jhJo60L
Cm4gYUNFFHz6GMkUZFdQ4sXxMYNce5A/jM6rFvBuPBs1fkXkmVBOFZcgvpSGGsM77ihiTSCo3ozL
4UjaEM5HhFGK9PRDa8DVO8TbpLsI7sDB+7NQJjjeq6dZjPmXSuUMcfhQIDlYNtJQaMP3F+jraM6X
IOY/XJBzSEe4GSQYQ8LgiZ7QzIvQKtx30IravcO8JfPm7MKV65YiScbvt32K/4NWgSA7VinTCsrf
EERs3rpCkeTPjdXrcP9QlO1gCaGjEiJcrKeD+8ckFGj/+1sm02ej1drW8gg+pUi6dCVMxHZFghrR
VGAeLr7lfWTv+H/C4PU8TGKbk8tz+qr5m4qz6VNi7O3xf9OHElTXEjG5R0BeoppIOmRJSVQ4J1Hx
yrEud+7lmYqHC2/FnrFqaWeurjsNLOfpn1da4+MfRa7dL7LNEERCHzUaZXQlUFhOzFzHpzH9npUM
pM7+YAMmPGRkU3VPJZyn/66XfFKKFCOs5O9tyFwzFKhzBzXV6q053hwtsydP6Oey7aKLMVT+ubfL
hOJsrq/FKmizgf7YBRfzilegVH92HNt1VweXZwEeCif/Ek++o/FtrO5x9LP637HXnJbBgQWmTi4j
52fmSe/kOnhOTxymk2RdaCOhLbON2t+w570IPiXDpMrc1zLsWysM0gMGB77Y9KxbbD12fSBjhGqH
Axoq6lTwRnnBEf9nkiouE7Q/lQMFSsaE8dV34UQx1fCKbG8tze5/z8Lm1QF5UJ/dc2ayyeJ76eE3
hJ2atEmtmmncqxbKpY7nzfdA688AHjGuEE0Oo+4aSkOdu6A1ACsa7LCyEMgvlwsnumxhwIfat7/c
3b5se+XRfZyOI1XcBZbYd9trHu2g27YzRgljW6jIx4/9Sd+8L2p0O8Wt+B9hAOVDR7Du50A3FtJE
OeCAQoKjqSw4IN4ke+wy98S86ChomGGf/12S9p7Z6B1Ivvdg75pQ1YFvPUvfb0ZmLTEAUQkFqnKN
D+NrrCe5VME3Hz6c+42GYHmKiBQoeE4idd3NIUWm8Q81hEY0jrob1KIVn56tctgr+G+A4Ltp/u25
Lm3/VXqVc7wGrag6XCw7CMF7KPcLkdRPTX/hoXCdakGAcfRWPQBz1wLZqve93I1fMDjBxTCYbwne
FLrFlGcytfCviFDteLedH5Cna8PRY/zeIJL5KeRT9CfAwHMadoQFq4ZXU5I66SyDQAZ6pfdGAVSh
WwotDmjz32Fiw5fNjK30NNRtW7hkyskH1E+ZZeCim/tb+dK25ZGoskHMF8xWVOdt/Ju1xrRgv6UV
2hq9T0ezpp6PM6I2u+37s8I21Y5RQQjml3WabENroQFVoiqJPCeM46+80OfJqmmbl/6pgeV3mabv
rRgu4x1UPueN+5kLEVzCTW7Mi431Ag7g2yw5rJCyxtBB3QNZrUX7K+Ce0hdYIUU9ShBEUSPo59gn
IKwmKcR0TwKY1pBIgCFs+/WqR8TLFtoGM+XwntFIiZIABrUeJ23jq5PgJ21TrETr6tVoFChuYgX0
vduhncwDPLOcUfkccgcqXZKWTMFbB/8zTsBwKPtSwd4IAQ1pDagCfcsx3MhyvzgqLMfJb8z7HDPP
qg3AZYby022WdP6W1cdPQl8O4QkDFmcOOViYoL6rpm6olyHX3WbsJvyjuemK6u9P2ymRcBI1nqxr
1NX0ZOQauMeXqxUeV4oKxPp4hDljDN8WHl247KJq3/GaDvQoYM0twibtccZGxYk/o8MSgFqHhjkM
ZuU9B3/z7zI4TbTA9DQyAaWsK6bkVnHWT+Prng8nvsBtnMfX67Dg5Tk0vGeByVQXEAm0xuLFHpdq
ZpAYRkQ0u7OR8Kp4QyVQCsR99GRb0DhDJmVbaV3kLNhPtTn2eDxgnX7nzl1aSpdxLvq822BTLLOn
M2M9I9gAHscLTxNsdraUJZTxPgCkksNrVuXPdTvp0NrRz4hZoyrsNHvKIkS4Zg+mW04u+DF6ylHF
sQp8ut5Ca7Fx0QVvjzMBOHcYQAQxOWAhry86srFcf+KpbblxraK0GriXVh2C7s9CtHmyn0+F+DPK
5GrSGIkcju1Vcvkw4E65i073gO8a22FTQQ/oONiqcJPPWd7G5xTHi4fi/1VS+ZEpZM3luMm+ZL1X
nB0TFy6xFLLz74be8v1HjLkFziq/QYqgtDgbQViT5BQrBwI+ZkD6+AbLDW11Df2630pffW8AlXQ0
jdq9byaNAgc1O+Zoq/sS/8kK3t9GPYOS2mP4ZR1yHLxHYtsm1LLGmBRrKX4s0APkW4HyKyzCaOPc
B/PDdXLD8aWTJEOep98CmOS8QsKePCdFpLzo/FD55R7uMquQtqGQViMpIK7i3mPBDRkbAPqZZT1U
n5aqYA2Ts8VqUG1Jp1QBKseGYg53wqCynJDXeylfbcE6hLDyoaoiAu/BcG7H56PA/+rm9y7Qx6AX
7sn0146brxW9nAkBizxh4w/7hsE26ejtZAVQS6f/O7FPkVWI/dKNCLm+TIpuE8sXKGktPdu5rr3/
gE/FTFv270d1i8p6E95KDv5RztYpP9hJWUeb10ycfVMiEWPKNSYr1BYcMXscfuqUGUpHsbf4wAbB
VXTRiTjtmHdUWiNWJx02yGu97M1sb1BSyf8NKmLilb2Zez7HUaaD227CKR4AMKMwMt0VxjOLEKyY
tpwvQ0OoIK25JExGwL3uXdzQ7bayP+SVxAlxlaJIP8duM97+upKuaFC0NAC5JnYo4LOi3Xn17xgl
gjtKVADmyUd19Nk41LLrRbdM9GiMfPLWF598geOouIsz6NYgXg2u6wSJ7G3bVzIDtD9pJcbxGrjF
Jw3KOH69PnXqwMLI7C8uTPYxmSZ4OCbo7qMcT3dk71+Vi86yhFQqLrgyDMSVEFOR6SJ0usprsVpO
IoVOnb9bJkwgHzfqqVVTzmzbpR408smxBZ4d8emrbKHyI/siJKi7cSANgvWljbn5Jn7Ys/lwyvVK
KeFm9T6au38ulyuV+OiEbmGby8xte4ZHpcahLeo2M5SJ0ZTwc91lLcnCweCRsmm4whJdNfDqoxNq
9wwAU8TbVwjF8B6fStGu0cVGMcGATkRDZRZEOm4EUyrBfGN6zMN6S1nAmwPfMOfWlPNdOiIa2Kp6
igVOyS55xj9GWz3lWt7a6l9o/t8qzP9o4eUh8Q4PXIDX9Ipj3wMZBUC8JqGf2JRVbvCIyXGSN60W
Fi6W5FVyk+nrvA3vj97HOl+0JZc4jvUxXTxryDbKo5nNEXk3M5nlSGX/4RUgnVnquPw1idv/q41m
vRQUTeiC+SK4EZcC1alhrFeugUsRaAlH8KEjgvXp68Vq2h2fg2vRemxiw5ZvrqFomCQiEZKNvw+0
Ui831Cu3IiwcTAcTmWNJY1SFI5GowJltD+Xz7hIzW5Ux6JwnIi1s6LusMjaDLWByp0VMifXn09Wn
seqVb8fTgXSF0X5sAegN/mVMAjcY0LVb/nrgLOTJrWz4/cS5F+YVjaa2OG7XQr665VZC7pKdMmFJ
k8CA5ssa19BGxCdQFYW7+YY/RbAem0zoXL1sv1FoSWX7o6FJ+vnwhxwIePp5xpowL8ZRDXu2a+t0
y3gHzxa0DhYYTJs1DjfW9LEzpoYgVFLhJUheBTjYQV6dV1FZbrBXx+/zU2zsT/uulCR4Akux32OY
0KGTppU7fgZgRDjpzPs3Fn7ps3vQYTgFhXhVtO7lP8XOHiEI6M5S6ceKHhrr2A3InGoqn9ORPOTh
iaGROs3YaD9i2UvMgMmQZk6VIexGevOZsl7nWNbNjavR7CJPWfLaqp9LtM8CCgtmhY0+lm/JMgLh
L9YOZN6k2rzr1uG92/YgQMyOtJQCwnkqMmG/Sdzo49r/1Lu5ly8NpTUy/jUOzmFQM7K9Uy2rgEjP
bW2jppHaWqNQM9X2z5SFQrorFkdMuU3PER3GfS8ZiwpIEMigUbIDyTnbY7zDtpgmBLNjwk+opU4k
VKKeCI/w0BaiVf0xqLVQ3iCm/Ji04LvgTAbHyUfbnKO6Cc2sQi+HiCagy8l3+9c1487kdlMvVnoh
SMtfErayGB2sP+89ixXaHjZfLZonsPCZJWQWIH1Zf+ypKX1Zw6ibaJI95aMyE5WAvJas/QpRFgR/
HX3kgJiczSmLDwGZGKy+RJu5PdufxQR2BbEOvLvRuE0uMiCkGlVwT7MmlDMXROJ0pDHI/XtglgsH
hSwbtXl4sNgJfyFeB9otj1KRAJP2TCH3YlcHEXLxH2qcE1xvdk/jF0U/r6E2qQz05thGePstqTsw
3OF26uza8rkjAeLtxwzQV6/EhBKlz4HrOG3FEo/l64ZMeivoSLphgKv3g3xx2KFSIvOU8uRAs7F4
LiOwaWamhPlX2NrQg9coRf+KwBiwtmbIXE3BHWZ6eulcmaLLnX9HcQyc5beqIkb3KPFdFodVzShB
ZgWJ670toPkXDbCvthugP87Ij2VFAeYUSB0tFB5Zp+U3U4NzgHBBXIlovfCy1kRVTJL2eBXookRg
BQK9f+NZJkwqvmnWisToJiAGZobkmkQclU4V1XCZn5NsJQVqGrs2qlnSSnCJWk7R3iNJOJd+VwEM
5M/NdS0YqTqTc50GP0xrBsuxWaumHDg3hcofeWaxPrjggzUG1c+RcIPtHIgn/bzEguJJiGzfplFj
i39t/riFLueIpSB/Dd1TgqJ9G3AoQEkerVnmMHkTEP/3FWOc7cHj1zirir2i51Ijmk8qgxbX0eOM
WuDwL00CJK5m6FHND7SYubwocXUOV9wLpTVo+xd+K3y4LWfMPKqeOKx3MC+d2YxDQMLCCbRt24Md
uVHEHuDVZr1l+GDlktvLMrX0kb+GePp2tw7a6n2RgfGx8JcGow143tS7R7Gx/L82RDXQ31w4m28i
kEF2y/C4UAk52pUk2dcfIKBiyngOrxJbjUqcEwO3JkRPUrfipu2fAlcChRBwtTk6NFZVXU50zfCu
3uebdFaPKV68U3kauox7Bsc8rjVPLWQ/zEz6OCsDG/YiXPW/QULyBIuaG9yXEsr9KxnCELWlrXXL
sgyIAmEuCySwb62tmfOAF1BCzmp9UzCNxlvr3Llvgq4dq2dqjdoA36CPxLsR/d3+hXk/adNj8bxx
riSEHGvIY36/LkS6rSsX2Zg0a7v8p7bJKy/unI9FNv5F3r5LlyquUVfY0Yp5OD5aUrWa6wX8Tzz8
ey6siVoc6311hOUKIxnCINEEZmJWISUiW+Q83qyrOskQECvTorYkq3SzOtDOihXArGomBlhF6aCJ
y+V9tal+pleGCEJoLsQmI5hwSAnBIq6YPNxc1EpxqLaL73cCgU9b6z00c39AxKwOJ2k60y8N3AjM
zGdmbEBSGrT/ocVthh/AlmNQPkCjo10UsXkHoTaVdDCdQ3l1fuJuD4JpBpHsGCkbYqm5vq6Aw9Ra
NN+IrGW6o2UQA4gz4jNvCrpIGoey2yqzqsHx5UPsxXnMfCJSBw2z7Qa8Yj2N1sJDNgv2zQCL2l/c
dewAex1GweWadQXgPDH4gOnwBC+g+9Xc2Lz+q04RP/GBcCgvGFMOJ74NnM9/n6nMg54j7i2ojbwo
CV2lIUxDJOLE/12/c66EgJrtP/qCocbeDGjsFf8wtuVd+/UPy6OfE90SJPqd/nJ89eAHPf2zVBDt
UXlVXalOjR8wCqC4yJWBHLj/XEI/Lilg7J9f+SexLxVD3nmEa7nki86XXCKJjnG1arEupPl126F1
R8t1MQh1sg6hjp8FxVWkIzRUeW3WIXT3I5N/QO/rvYmxozeWREflxXGSqLJlGqRxQOqUh80orIXF
fDFQyQzv2wJD4cQel6oCS03wHAabZZDiurrlGPNMWkWC86c3vnWLIoA6RErg1Fo0ZcoBCXRuHVEv
VcuOyVEanh8+59X0BtJIn+HiptcxY3shgGjWovudn/9ndUBPAyGEHiqSuEflpOqYRyXqFow7iT/F
G7sh05x2A3LqD7BNOpaVAKB+Gjri1G0A04y/i/RpP7+jtV+VEG4fnT26rPiUgL5u8L7OXu2ozVPK
L72AqwG6QQ1dTpV1PbplETTxOg7mB4+VHElpg+xCQDyITpDkZgmohXLwhmEObjdqxXtMpAceV/Dw
+c2QdBd3biozisN/Tl+cZFg0PztunsQKyKUn+I+Wnsw0r2Viz3lNtpBg6+v7TUBske6SnNWk2QWM
c8F86f1WZHCVHGMBz5SW/g84X657qz/dz8l8mXYAOq7dqk6Qsl5UoenndiUl/KRibcFdp9gbUGkT
XW2ayqoYRMnIomXrAemCBxg1CzYzVSH5a6XVVSZwo+E+Ohln+YN7RzcmpBkABr+bEXeP5zocElmF
tycPzhaKypTmAIl8Vgto+YXTYErlWpxNy5nk9rbPYbM66R+uRLCu5weCOYEOHg4JtebFV3H+TJxR
ABnKvl3KUyyciM0Fzh66NMIRA4pkgoLsKtZhDx9xmrqjkbz4XkrGyLJ0kPpqVbadls2n1NUyAKRp
V4nsbRs4yBSwM73agb730HTXu32BVtMNeO2fQy2GCQMptYnN74nNSYEnTdCM80124spjosuq9ZjD
5J/hFukTeVhsjUtZ44YkS5+J7VpctpJJjNAHCvVOM35OMusZAfc+Fbd7A4mduht+LPMlPNlnXrZ0
l+EqejYj5S51XGmAh/ojJuaKENVi18B8Mo7W9yb+k267CDEV4Ytj+bWby9cKkFuiZ6chAzlvVFeB
tAeZPuR0WCprAON1uCOniFdoK/uXkNNUbKCC67Mp4Lmi8XkjCKxpVMknkj+A7xX4vPPo1xs6RXrj
gLv6s7ulHY+hBjtNprjXBfy1hJ0lr3CdCcpuIdskdr3UkOAnQ7hADw/Y5KWCdm53E7qGVGP4Xrax
50sMI2XTyMhLGnaei7RLNAfU4MyzQoBu7Yw+apQHp5Y9S+xPZXJL+nrFv867lVY52KNTMe2xvPAc
VagPUU6a41eMDou8OyGNVJuh/g0xq1NJaYSPcVZ0vYOzeruyC2sNNiC4SaR8jk/zbXNKEz0g9OO7
bjcKQy8X+r4qNrLh5PFbEzdm2RFClB1P3X2PpFDsNH/kppBtNAH0nL8NKzL43VWPS1AtspUNGF2h
1wmpPf4fJ/dov2keJ/qSbKgPoy1rJXNfaLSNfWt/te6jsFQQJJWIQkj1jLhG0sqJvtrnI/dcvuuh
GK0rjRQxTwVMsfRDxZmYs1XYuvBZdalpznlpQizpBF+HmGLzNdZeMDNxIJdgjTtubWeWDpIB9z0D
kpnGsOWynYTtqoxhpJUq1Y+o4VX+6n4wyQAymOMizCLTkNcEQ9eyph2QtZH64w5orF0+C6D0p8KL
UTchZ6Kz9wzAWDjlRZcOX/J1wNDL62RQgjZQNKXY74OGugG0+JM4Rbc/S2E72l6UoojcGu5S1eAQ
pevOp/04HWyVjveGMEiNTp/t5Lq5xMBMFeQ8JMhiXJX6/Qk8vjNAXsBNTbncxQmduYUkUWTQ8TMI
A1SyoLqnnPRdB8gXKTTPpZUjX/bc/4ypkaL+Bb9Lp+UrnB8taQZucG+3wgRwphBwAT0dYL+ybF48
7PqdG1UV5r2L47GGNsbHImu6amPrNWREL5qJESt08Pk0JnzO1KPJFZkuyrKw2MMD/4f3DnE+NbCT
ZI4PwGvtqXg1I9WIFd338IObrYrFDPwjRxkgJbhePCefEvat3mW9+wAGdebbqKJXCfLJMWzEkgI9
IQyUJMM5FfQxSPkBHq4yB9c9RK1nphBMjMY69wrEH8194OHhyLcNt1rl3+9MoqUs9EQSO7dZrW9g
cOQ3DBadyurYsdPEziwi49m536HRT2hWvzR5O4Pdm4py9RgEuGFKuvVDnh/EHtxD08vRuhVoxmbN
wfpueKTY4Mx/I8AH6grO7wE8gGX5d5Xp6GvcTlhYTqJOTHigzz/lqdTNIG2OjAxendQ4RfheoTPX
B0gbvRWlnkD85mx0L61XSsPQ+m+IrsISFvskl4DiM5VOJnA8O77kQa2/DYpzH5gDFKXShEPnJHCF
ZKhDQX88FBeqMpQxOWWkarsNSG6QPOLci+5rH9BSVmulj+NzcONb3oLdkcb1z9HBwPDcl8DuIEib
qtRVuKVXjubR2EkZiMbsGqmrDeveHFeWn/i19mDJdb5gC1V0ZWX+u30SlwaTWc3AueKn5QM93xCe
Onxy3D1rAHE9MBVwDquAJC1mmg1FcvofS7VKMc7EJy6uqTpBbv96073Y06PZTGbdIq2qUG2FsLdL
283NArAieDWZ2n/Rb9pkhutCOTQILh/A9kghFvS67YHkW/ThbCUIRn+ZkOeS3JOIH8Voomq9qNTf
gfoxtZCORHMi6aGskbVyuqRprNnpup/xSYfu6Lws6mmAFzSa1FuXrsmvqhxgCRYvHc9fL1bArfKD
uRxVAgyfBVzo3LM+enBPGuNxuBZO9tf/uYlhJ4ZaRbZODPWOsXJBulSfKe58BGhvtiFirT4g0GL3
KcaytyP8+Kbm3JwUWiQz6qgdvN999NIi4t9AayaK0fbeo4MIznKdjjoHLoiPbE3cPN1nyftLlYhJ
NBizW1Qah/4tsVnf36ReLv+Vt9RAQ0/5KSzoEbJvWoq950yQeeiCI6kQ8CohfbVEAMtPgNKB8s2o
SLGEG2vYdTkFrPvwDeWfqe3zUDIQyjpU32B3ODDc7eLggtLR6J0jBOX75Z4kqoFpMB5zOgVYJvHz
gml1Mt3jNpWie0U0Cx9mj9464+jWhkLYrkX/oqFcUn5sJRxS2TU3Wxx6lDm4Q9XU6YH+osV5jimc
yih5/etUVCUQM+sD91R2nlXXOcdmmafCM6K1T5MAWx9H27TKlDTZHpaEXfYTHYD0jAS1Gy6spPD7
COs6fz749E6Lk0PvBjO35mO3gnBwkiUyIGkFn3xFoN9SX22DLhrDPqVQug4CnFalfD6aVd8/XETD
6YifgelcFvy2ls+qP8zMrcmVXD7jsd9CJneOyv+cFuOvIYjrJn2H03HbAVawU8Tn5ok66aMHowbW
RId7Wf8OqnrMVGMQNlsM0FcoFc6Hj/v/ZsWdfOLsJhDl2PQ024PEaEF+gaDb7hHoToJ0fLTNhkKt
hjWO9p9GR2WlRYkBhijpkZaGnfaRXLQTCLU7K2vYx/CPTlsqmirR+ou8aP3gwxPIZL9mzEmE5lIw
62xFT+Jm00s0J9RRc6eRVDbRGp+i8nA6UedWVrIOENvVkQlu3+uhGu5ATRY0GgXUXEWCsb5l23OO
Wut9a78+MfV2R8uOyNsp1iCSfKnuFWGJ6rtlPy+ztDKEqmIQpGGRkryMEO1Ww6HCaBQ4vclLU9Wl
EI/BVkRI75WOJSL5ZEjWePoRUu1P+ULNA0RmA/8aZXnGjxPK1MWw9+2X0SID5q5dc3u9S6fl/ZI2
Oc1DFYgMmzucNR2u5V8rm/VstvcNXnR3ry8cj6eyq8iYuZ6v3beqODBKd8vato/mLw94Apl4GJTM
zQv/rr/NE+RbDrySd6a49S3tn+pe1iE+GtgK9GIi9lYx4gVsg/iFmn+QI9x3P/VF+VgeGVZfSNjQ
jA4Li20dBHOAGxQnCdKCNIFwBiQ9zGUN/7Qdb60FwNMle8kF6XCpApsdIHTWCKR57KXSVcc26di8
HYr0DJcxnx1KHLzJHrHUrytZWzuRF28QXfPeUpidrfqrPjNzX0oIxJ1BHFzGOPapFoff72GCQCOI
iDlZYtqws6p3mXNWJ2uU6RGagSc/tjtBoTxzshR/QDNSk15qP0roskF2cln3Fdq4ipWQdJrnitaI
8f8knrxE6kX+NAKSSqOfPlUbLa+z2OZP3Bv8ZcYmsj8ibHuCOY2LsWkI+hSKeaAdFuUmc2Ps5U9e
IiU/8xKSFn3PYKaxml0cYPNu6fDUaoLapn9+vtqvrRIvkPNPmtjdj3McvNaO/bSUY3KiIp7lEvnY
+/wQXrPhUANU4FSFsIMdxe9Pv/2XhNHBwn0jagDgar+XTlgw0cxwoflV1GMaxoghz4EeZBf/TYXf
t7mxmimH+ozkYWoCnlXFq1x/Et4Jy9+Bm4J4Ncu45VgAOWWMQgNOp/NLdI3ggYJYb8RIXwK9qFJD
Wgh0GGTx6adc9XO/ZwAqzxqsgkTJXIMFzTr25zziD8lrldFsfFNgEAgJhYZDPsUWR2wbGSrY7NAK
+BpXgzGQ2VZc9jbSGx12c15uml5tvxTUnaOJDBSgKhkrGgHEcIfQN57vsoIZzm4AyLdc2H5oc3DQ
ReDdZqmiIxxm4JXjdrE4XNVTt/xuAe2H/GLwnsVp369spzYmc7LHhQcEl4IhPY1PU6K2EituV88S
CXbBYVY5nN8JPjba1ciWFtWfVj3DksAmKT+RfEw+aoOApG51ndptV0vzOw+Oa6I33f3OLP88EyZh
T9dgEnBQ5KfKDk3O29CyGdQvLfyTLNeY1hwQ+o+qpyhJ9QUE90lsiU7iKJYbq4x32aifjAbPWyNH
L7+adYeRIW89ZuyE1uSCxBbS+ErIG6o8uK9HdlqsiQJtAAUo+mYvwCo0Av+1lmnqgjiSGiUFvgJG
Uf6CTJcK1cW6GkATkdX8aUzc+r3wt3UqiHXDki7mAHZ7Ck7M6619SEayvpw6SVsxe1u1WR2iJuqX
JtXh6HmNxTU1KZVifxiyYrl13AN70fr2lVzDmiQ6E1YDh5JKXW+qOTfWHczIHEUpirujz+RMGtm0
XPXoN5Rach3H0UKq0GpPcQrxmkdgHAoI/QAMFqPqH5QtPPMaXydpErieebPNE76btF3zxQf9g2ge
+jEPKe6GMkHfnc8CHDuOGPb1v1rnDEqKMNEukIYT85arKUqK96GBMZNxNtkIEYqxqrK6imzk4t3v
N8m11EfEJZaiGxcoioyNsv3Wi5DCeM5gp34g0GB2Ewjjm6DLvxChGkHn16jzmHq/5ndwtMxge05b
WVgfantwBESurERuFiDL7JLN3uK1bwoRaksFaHPMnDw4LMZKcEjTe/3EOI60moYeCJjoBcaleLLi
bxv8Capg3waRYUc/Iq5jhd76l+/v3u/0y+WAreO8Ko9WI1ukRu2F+XOixxMrgqsLyY8/c8+fRz9t
dIam+Wyq4sdD8lC0+IsSWdd2ptNbScOJKqR15eKms5OAR+g2OPMZIlmYgvsXm9zkaZPlpf8EpCXC
4XlIBZqgWJiTiovOvOxnZ70IuuR4/65cTF/SUwrpgS7QadhSUFiBspzIoIzOCw5K4HVGqNMAV1E6
dxf+VhpeiGHRLxuWpfoUAyHkR+LlmfDQY5cs6mRHzvZ85pESsEgLAHN8XCRlR3UF9lnVmho6mOMx
pIw+Qe6vjTgnofliqbXRqC8wQfDIm9p6JOKTeNbCFduIKiIC62YiZJMtqvMrVnE+0OhqBYrVENPq
k1+YwVBfs/zlXu7bg50noUvg+0J3h9p1+UV70RDPeK3Tr/PNQgYriJULJFGg+jYLpjI2PPaa7Kjv
E+ZYu7gXX3GXojWanzIhs3Hzflq+UNBLtFuA4vNbW9kk3z8RVhzMaxMpqzmD7lqVelZdH8OHqAon
riSEl0DrLarquLQfsKA0rfY+WWxumwsBT+jQ3k1PGh7lniT/ieOSDsKMcOtkQV6vQ1zChGmtSFJS
pThFFm1g3HonC+mpVr6Aj2cO5j6/rreB1PqQncZoJoZTjEB371qWUY3fw/01hRY96Ci8iaH7JYA3
jzLVPBQmKavI4AxKUVyFX7mJYYDWRmTXs3b7Ka/2YjalIVQT89ZR/KZR2QzgpzTOhPLTTdcu2p/P
nNWt0MGXk7vpKCRp0TXJUPPFHf+BA2X/SCoD/aEemclyQwUUYr8HY38A3Nz4ZJ/QIszxMZX9w3x/
P49h0NkV1N1eogh69nIb5SOaIF9ewZRn6HPsn7tVxyYSgL1QHk5BRmsFR2RMIQOTh8yTgnO5kwhG
1Vv+5jwyk1QX2l1u2AnWjTHBIgpaQOTO/58BUT/HznPduin+hjse7qTRkbR6XwMc+6OBTtpN5Hvv
yxoCDQk38J5UNZv2HorApaybKrcjkPFrrsUrI6SVXDItXJYDaIgY6QCsKUX5BH4CHgO5lRuihHaM
Uw6gyMFv8+7biq3R9KsvNFWGkeFuzsFNu3qoA2KtaXllufFcWLP+A0Za/ILEgRB30LMXodyUj1D8
gHXdyI3Qn8LyW/6bAYC38BOw483nd4ApaJ2lgg4OXn3Wq0oAOyb06a3LXnwWtB4W3teIFe/H/Zsr
7m0rWkhIAxuHDQ4uTeD9TmdGmmjk4KCjw1BvHSjhnRmejTtLiclQVFHGQp9hDRwJTpyt78ZWT0AK
Xe5RWy2hFB3l7V5F4OhqmYAmz0S4UYGuY8cvsigEF6ny6Bpw171QN0vEF4Ec7GC7flle7BZPdgHS
qOS0Wh+ZY0g4J/nQzqOrxo9apbkQFsoemgrKfCoPePisvDHcUntUBv3Z5TMeqH7dC0ph4SV4NMfL
r8PAAWiBLpeeYx1zLObL4giPNs7rgMRQrGTqECGYmkpVB6Ld23rJJJ8+mSYPoPmNixPBSPfiy3D8
0ZbZGilxT8vvcibvdbNQF08+8olhpAGReW+nEmUKQIcLGNdOllexeMbr2SIcc9YsC8aqJbRKxsDt
js0mzpTu7RgyswkraGtNFVNLDg5qFJKbnkptpYxoSZTiPWx3FIXaCRkAIis8kPplphB1kt5cJBR6
U/aCUweFmWRjS/brsZxxAa321jGZuTdKafjEGzlY7VJ0KjAURw7TObLsPo31tfGOJRVXb4MfBQnM
JGCggupdTAKVcbwTsvMVdwkdLNlU6tyUHEOqGBMr9VL4JrBHiub3LHMw0NUDwpIGvKTEElS/FjUG
uQoWIGoCWh4EKnfHUc1KbnFrMVuK67N4bCv2yMIVwxdbxg1Nr0OckSsSaYr7sDm61M5Q4sYeznAo
uuTDVK/h3sym/xz+my0LYAENpsq7O77AoFfvV1qfwbwnNhffd6wfMFLjdqgk3zpElblQKt1lkWpV
Szdb3DJpDg4EkR9C0Ot6oxC1Cq0ceCoo5wKNvbOUUIQqJg/6CGspSjnXJ3012HKe9WgU9TZwDNDp
D/ADQX29JbxF35AhWinrXE4gN+VRhwvqxLNp1i6RRjLcPf5yB0/h0MKOCrbbbUdKlc26EobVvaWG
MIBOe/RQFUBWJuHsZ/qULJkzhbAszw/SIzLfUbEiTOWpGflr6DUlSNd4dCtmSvq7qRn0llgEFjOT
sfnJ2d91/aRbU0m9ipjWBCQORzk8iXoHhnY75BW/hWcWJ1FmoYkLJ6552/zSrkFTuPCN0Q6l2k1H
hjOnfQ5SFiSsgOhnZu2q0bg1ln0FFlM9ubm+WVACRbbcQuIjogOdETKcLnkrXXL/UfNoAY7ZFUmm
MKJNyRl/GYt6ui1Ri2dEool2i5rzGR9BEVR7TM0x6FOQlhvcaY2rTuJ7eNszjTYZDV+sAvrHfwPQ
fXSP7VVWPVDCMQ6jvUx3SLh6fdyLSnhp0IkFXaMw84SdMs9kbsZbZ0dieFTzf2GK3d9mZjgHBLz1
D/dXj+yovs/ijpPxJVfThzqBQ4XBuQbjnNLYzAR2R2G57uO2FNwxlp6W3A7+qjk1FcClb/uV6Va2
JuA4gl1kfGWwvdWCdNti+GbynEcSHqjJRWJdggHEoJhrFWgwf/+6MS/5yphUD3IfzmjGf4WLHIea
WC99XrCBL+wwICZi1RTsV6jvCuy5XXFZCIc4zpiFBgUtzWeM31zYOsYyfteAxo3oet583qGbeGSS
Xo/IiejKxr4z9DJV9R9ySUcj3KDX/JwyPrJuLp2bn07I+Ls6fr0mtAB5nE9usjndqwZyYYgW58yd
mcoK1mY07Ye32skENjSJ/uDZU7UTxFxZSoadq6P9wwKabo8FcvHkGrxafuCuBqTafFFrdpeQn3LE
qsAHG/eg/O2SpYRyEGh5a5jlxT4SODR2/6uWGMrIe8nAfGzH7EzSrLMU2UsjwJecAdl7eKA/Gpok
N9fVQ+brKcW4T7LcryqRKtZDfBLoGNT40bZa04pDkm8FWlAlOtdvGJTJTSG0BSIYSvYMVmq0sI9u
+NUISlYNmFknGy9zmG02IVoIjuuFa1HYbNYNarkRyFuSWn5VW5WcAFAahT2F/vtu9aviE7D7zUpl
+fSGEC1nqd9Ag8f/6jSqI7QSpSO4jvCpAlLlb15Vq51rIB5fLiocnK32EmNzDCdvSOrfFc1LEhBN
Frl5cacgfnWjQF5oaahSlNQ3J6j7zU9Lb4cURUWyxXlbDgPROhZTg9kAyLGUDuEK2S/uYiR5KXiQ
bC+4rewhfmwVH50yM3/oOUk4bDUEKxq9O7uprvhLh2YWQThXaqQysZVvHQeavoD6ZfEXtzi/BHGD
pY2kIMIHXaOmBv3NvVFGb/YKGXFYr2iujRRsgMqvDpYrh42srMCy+1K8uYOHFEkX6f6WyICitz4g
wTo7CZEwBgvlkedyYlsYZAzFIz6puyH9PwBnuNSEr1h0+gZU8SdSuFnSCx4ZaCJZyV3Db1EF0lVa
KQiM/jYKtVJm0A1qOK3ZTftYiggYWIIu7K1sJyNHE8nDHzCawKQRUh7Vf+KtpC9NIk0QtcgogkRq
DFFQqTO1vF1mPUw5GC2C0PUfTA0SVH1+XQSHLrUd0H4Lx759FZJQleufQjEvqpwmrSz8XQPxMux0
HqGsW+n7r1HptBwZUYpqtWuYkUeQ5YkCIdkGwleMP0/wTGbFixkVok2mxqvkMEUqyME9i4i8Y2Hc
bh/U9sT+JkftdVC36X3gLBV+LjhqqZWrsX/PLfAx9UvUHhymtbBe+IdMNL0NYvGxUhHBk0DOKrkY
6TRqhMFFc1lCJqe5yvYU0iPjmITySs+qLswRq7sakz7mtIPZ9Hl/cJSwE/K3LPcospTjF1Bu0zo7
jubzxvkn05ef0Ufa8RjpO9m1zcXI1WY4+5J8JllUkqCYFXv1tGRRau72n56IUiu0rGJoNBJtwnYX
zy+1wrgkBGuVSHbjvP2x+rSm75aLyLT8FQ+XVmAaKL2g9mw/kaJlDWzUZRFgr7DWHJvf7zbMBrvy
tuAdS3c0dqJ2mbU5Ad+Oz4Fg1QGo75jeX2DyHTXal2+pB5bLFDefm2ohzXsqwRYl8lY6RTNNAVCK
e5r93zOc9WhrRJ4FPKng14EWBGZeyVcBrLFvKDbry8Mnl7UWPi3318kGG9Owf60ndRJMLd5Hg2cD
TqxMuhclHaS49vbRu0rgI+oT2aZa4YNj1jDaub25mLBOtliqC87X2rYK38xGfwy+oce8H4jQowxZ
WA2Hif0kEO9G3XoDVCDVvMmmYJGmVeRRAKFHRXU9FZyekcGXbdAOYg1kgfKbM6g1c7vK+TvZYFQy
jeTZO8WA6yw/IWsEBCsk6bMQZpvKVDflvuWtgfdGV3FemMjRKwU+c58yLyzsG1HHfSBPfsSmwWEx
hOYFWDEDBjF8/FSkj/JRS8Y/jqWu5SlXO5BJKIf/mO4P1xLDMAuXUlgS25U1nYwny44xtBZLcst/
sPueZ+uoCunLUHt6UeRwcvz3Dx0wiYW8xJQESNKJXCSnBdtS0zVppA3WToEwJMqJup1hysOL43IT
m3Jaa0CQ6CMX6tSL2ldjBzCnjz1RmsoSHU13fIrfL+r6tCt6KvoHcBvLb0rvxQwMosUY6ZLZcmZK
UKrYFi30pesEDklPT2fpLcUJcZtJFPy3/NZwlRE8VTGZgSyyDDZnf5XJCeWMJODY74PtSC/IBpaC
DknBh5Aal4DOw7Q25tHpFKIvkyRWWWP6VE5J+e1M4ZVqoRhauWOY+tqJ8JfzeJflFH7NxR7AYNr2
n708pkyNB5A15hucfLmmf4LZ4FIlz6tvSqNTa0acCeYqw1iWUs/s++DrPRaASkKPs49NSvLbuxgt
qtl9JgWHbx0OhDdMi5EgX5Vlk8YNDG9Glf1Q3iVtwmt3qYzOva1o6JrmhqoQpHgkntSgUgsaEzT0
KoKUWcrr64oNz9foA9GB6AZnZndD9Bi65HxDuBr7YO2W8jg9P8iibz55mfmlTwKxDE1EbZPfgVRp
WGbAiXUtLOk+rVoLnwS2IrIFEeAWroD6JgNzAQt9xim/HRPSngZcwXSmd/VVHR37pyffim8f7zK7
GZyO45RRyA0rhMIjGB/Xa5JD/jvu4fcqXgcPU08V67lyV742apuPiDWEPVxarhwJu9F6+ZCbrBh4
quA5eMfA+IxafB0RwZJZ64TnOXsoyK4xunOhPrd+SuYmmXgFsD3BtWeRfDopSSd/QBA/j/QSBFLy
U66yYYYdOQO1yClMKPvTniNwoYyAJ/kAneSHVkn7WGUyKawIwQxQ9zHGOtl4XB7CPOfcdYlMBQlo
381pHySixDfuqxqXIvcpMOXdMtyn4ihhh/OYeR1XnrtFmy6ojPguPon11bL0s6zQPhkknGaujYo0
Najjq+6kR4xP1QUxx2QmcI/imfHU0IPORpadn+VajHd1EwZrHLSrIpJvbNRofwv1i+9dcnt2V73J
rmSi+E4Vu+ZQ7zv9zhEujVn26vA0UzRDTF2cs+id9RuaEtsqA/0qRytBp2mi2bLlOumzMTca+w6a
ZQm8jEAmfB5n6BAJSiILXq3Go8+CGejDadVCV0/tYTJZSlS6YaYeg5Ah6K6IUNWG8vP/9Ij6M9ZM
q2PsvOgpzT9QAoP5qnSpfRrb09RbeggywBf5xyFUpTunbtLibqdyWMACMem37xXAyF9pSoLbbM0w
1AAwgG5Sh/CPi59KBNJb170YZdDgf/HOTDLhhtxa0onut17TJ6+ONyRBIv02ld8smmTTiti7Mg1Q
BuVato0veORHk/54qjhxlfxNWY994qpYkM3swIeR0B87dLduXgMaCNAuuoiB+R7Duo9VLPBMRP2T
YR1jR/2EOMyTE5CA436bVK1O6UTrIlvgltLaxOrRwibgYc6dOr9mWc4it9edh9yK7egCAmoD42rw
Yr7BgT0Rw5aGUfgenuO3k/WPHce5b8KJei12IFKC90wIwKxbD0DccbHVrYE3eWCBXQLBihUb3PKx
1kk+yuvR5y3UyVj/HIpdK+dpJfGhDxwwGRwcX6SXs4uGQMJyJmZPVQMiXKXALbuvuh9xyTNpwv9j
MjYtLM8qs8yr1AIyHaxbbY7jqzOUt+6u2fx63Hwd1hlhzrAGJD0C6T3P8qfnFZ6BI/5M8daD48x2
vlbUg0GqBUARJRsr5JqtLiBbEDAsx2c7kGz14jRXw8xNLjYqV38vzcLCWjPzHAlvOEEduYfDN3lt
8gGsj9171d6YMbg5CqA3Ciwi9omLmAdhn6DrxlHMaV7PoDLlAtGkm5sLFnwIa95hHOWATo/jTGVX
gnPJ+z+6jqGWeV8mmx4W+XLnkLDGUnKiIAMAFcM5gmhZYF096fj4Lk7mN3ANuuOQGUaLYuqj4Mv+
fClQd+gGGb+I1i92orkqDQMtyZs3WrgDDpHgUJppl1ZZ/RBtEsNm0Ka+I183NtJcVivy4WAMf0+v
OTbqM8kIEOrmu3iJDQNFYQE5Dbn43RvXhBCmqj0N47T4Fwlk45G4kYdV3F5pfermpeFpw2Eg3a/t
6t0/DKk+TL91KI3ut71VCyXW4ywktAzF9rde/U9i0hxHqecOrNtmODm7ajwr6Zel+5jQd7vtcJXE
MmZB2WsqLlf5EMj2u0+e1ahaBmiXpD8Yt9i1UCtkLr8cBs4dmTSMHWV5Bz2tC00FVBspZmHYesoW
OT6+zUR14ftDTuyoKKRKvgBTweMpCy1ksPNGIT+2nm4DeLLXMOOm1iXOz0nT37eH3I2QFJlKy0Ov
R5bNplOjQR25NNbA9LZDypItfBSiSnWSYlAmpR3BIsmOba/o1Vyz31R3VKSZm6Wqtwcbfs51gHk1
YqjEIbBWKqEWMemJw64o0L805sPMse+bLfWxy4j6KCmEk4t7W06OCyXzwvb5L0DxAJbJs5TUZLla
A0b05GJk2iR4u+N1fmr9JXBH4/qgl4ZU+UcU1Okz4AQ1kLU3WvwZr1di4R2g+nmx9VqfBm9y4XEn
lYLKrY1csfydEyH9v7buV2YJT0LUjNxdRcQoeAIAYGDpNXBnSfOtCeWZC268joWYrgczSIV6GUcJ
6O+eZoFTDbK4hH3ZR5JRdrJyc7Yk41xYI7OVmR5t9Tr84I67uGPtscd9t6CdRliXaofJRtM7pWza
2O5qjnBxKwpTFniP48a34lseZun3FIJOO5Bu+PjEz0woc8cXfTOsM698WIq1SYCZm7P7ctuHV1yz
jC+Vg0InkPMQG9o4UJpiPiUI92mf+fp2fKEPT7mym5aet15b0PFtH/Dw7OZSppHXAQT73zt3ztnl
67vZG9pWc7PHvnRs0XJb6ispY3jgGykwUjepfW/1elEkE2B33JGRC0pEvktXD1MF/oEU8iED3otq
GB8eT8c5thRa8LPrtnsqqV+AW3dzECuZenxQdT4qsTOO13rEHWy8i1DBgdw8YFM34AcAZlldL+GC
Bray6r6oqoCngruC7ghyFf6zO3KcN8GzpZ8Cn5Nw72+jKWmTbVoCX8gXc/SW1sEcdmPz4jchq1kP
cTgIR93fHxzwCaeJi5h8pI27VgpcUOgq0m/7th/c3EzTqT9LlHlcb2udmEO5CQC+PvRGh7mrwg79
AaqNOsB9W4tdRRXyvsiyEkU9OTMb9okUmOD6Xaz/8IgXgPIgNgoL8+VBRNCGwHAuorHeuoR4tQSd
23+b8NZVH0KnaJr7aE19BLWAPwkF8WeHXJUDKrbGHULW7tPf7lxrYWqwTfHj5xDSf96Sk4A4oR0n
ybMRIcwT0m+JTBUxLKf5r9+8K/KvAIyz9OZ+MCZR8PhJ3ULxE2crCOOuRdzq4OSyCpsJDZLYw+Xq
OHB6qDSwzVQQXURcdCs+oBqyzh1856btZN9uwPiLU5AqcauX0pecBuY8E3VjAsQD8juhAdiTbN0V
TMCR+uvJIH4GGzk2z/BjRqL3nm80BUYhG7FwcQDS7xmyzO7rhEmLaKrkRXOulaNeZVaOWvoHLxmM
2/PXszUAEbOGqSsq8k2q2pRqdFPAq0Zl7mSJrSVGxy1R0ylH+y4UBtb+jjPL1XpiyXPtwLHXfyvj
fNmHJ8uBbZoEK8UUL380F4L07JkvsZMamDENIrFihfH3ZbcdW78+K4lvVUJRL3gFxApC81b1qWph
azCp3fZCN+N7PQpg8CKrKbFwgRj/JK5yqivmWRu7lBGnQ+I9ONLkgtDTBvWvjgnP8dyaW2JZSZ5d
rVZOKfXWegMtaJQH+hHZLaNhUVRSNYuLLrG72QecznqkBr77g2l6WOsnlWzRNPcwJhB6AGjo9QIH
7lxf+sMWj93uZwUgnmHKbKZSXOiaDWz/Ud8/RTAuZfGu1wncWnfyIfzYmjGwIfhUBKOrt6Fg6cNW
fT9rclbNMZ8FAXM8C8W95wyyNkNfXOIHo6jXunB0/2JeEy9Vc2YdRYRV88tIeTMcy18euqZ8euHW
3dU/2Z7hIejbdFUk83q6EYjf770Mw2qXP2cOmNIWdWkg7qQZ1Jl2Giy3jpuAenslPGhULNkZRlJJ
oZI0auVRL8TtIM701pji424QWGRzHWTdXzVnGYpu5ctPIHKDRb/lUyeHthjUqc5iyWbm+EUPur7y
YA01BIynur7Uel/kHOf+Dr07R3EPmo771cfzRCNKMiB3WRdkBLFmBG05BZgaMVCdYwk0ekRaE8vP
d3af6YyIF7wzotaaBgpAUWL+lajHYOyLQ273xH9eMlefePFhTnCVVq1miJoXoVo3Kttyay0o0O8l
ozRhAoyQUjxAb6Q9iVw5m0AeyaNtr2J8Sl6Zmt36/qz+YLLUHqrwKoiM/Mnjl3Y3BBztC+B9/GuX
NyQCnzv5R5Q5+WD64P6maHRnp9GCZ7O3IhibpFhLCnYOrc4BQ2/GBmZ10VdbwuQ3YPRpBrkMVR+z
/9TLwrzq/4NVQVADAsHd6MdaXpTlC2bJapXWlTs2ETeD0piNiu8XDr067JPRWeVLKMKuPOvUN9mn
d08z4DwkndG0+l47w3nt+Yb6/jhg3XpqC+QoNYVNcAU1OFPZuj8J1hK7txiQsccbtfDiCMmJPhxc
QJzzBmKNZB3mcnCXOs6da6rHFmUHO3rBvev3YueM68wCkHpNezGfP8iI7cNEboI7PnKPleIzwciJ
KypRESH7hyW4XEZCDX9aiHAqGe/FZ2Uph4hhkw4Y7g1R/s1BJPoS1ADOoxKg7nmwOBQtDJCxcVqS
8dlSpJOa61YyRxx42Kf4AaZCmvf32jGJv5CVLMw/r9uM7Vx7CFKjHQSHI+kNfAtWn8KaOcG8NmWp
8m8x/Iqz2ghvdTaHMUvavb+ysbP6rtxn4oV1RzMweqy+XHeb+nOC8yujk2hcTrf2cx+c0IJzxKUA
GwwV2o14xtogptpjdnc8PquzUBOjRNrg3OYrEjCtcLE1rHVSMGz2SlXoEY8RDU3b/eLMihgRkjg2
w3NX9irdBfMCxUqw8U40d52qFY46TvQsSGQmvbLAnL053zRsv6UDgtTxb99OyY36DoYU701Pqmgk
NAjaOC6am8MG4Msauq8w3bVwAYkMgFQ73Bm1MJk4uGrHEkrC4BukagB261LJTPEGHofB4eiIwQSa
L8FTJcOEQ4AIo9HUhkaSlSay15x1ZZDphNN/Pblh29Z5veTVmI1bHrcDhaDNAPIoRbu1xID1QpvY
rVql3cAzCWT16vk+xCBlzvVoR9kxADMr3AUji0LlnMkDJzHTZzjYdooFcMFW7j5DVbR8ZpBNURE7
SmBs7jviu6Rv16g1BIZFlXuQcATS038nrYKq3ueiwzziCw8JZg/Lsc/I0XEEco6hj1fx1x9HNCmP
9H8IuNlt1ueiSN+8ydbfUVt3Go+t1fZaK5iek/hQYIqhp+/k8Brs+PN2FN7c3O1DvMtmgmuqfKl4
sur0Rb6J1Z3fYIViSerVPbKKRjJYHOixGL5zp5XyOLcQu4puhie59RLzbo+sUvZlep1QpugVbDm3
YD1IMI4vrbUETStdEDAW+xo+e4e6REdPLrfkCLFBykskDCrVgkJB+rpTdao1uPRWpRSRuYWF3kWW
+zIgvRrFgJvt6tIy9OqjFzWv++UXxRCcmJ4EWn4k704H0DCmGMAP3BKEuTsiMHckm4e4qigtF5Sp
UtltmcQogn5LLYmd71rf0D9mSoM2M3UHEjuMP2Se6ms4H0+rdFFFXapzhwe3b6QVELGfcAUWqkd4
hghsaTkQJ/ybTNE+rfWH9OX2/MAuiHznxoahRdueS6HQC56qYm+3af+taeHhfAom2biyczJ/ai+3
jxGuFSi7cBexPj5x9kYOM5yXD3O1lhFQPYlW+8ShvniSjEAc0omRbvuFL6eAImj8sIyVbcXLpLcJ
nfw/JAYdknT6HwEIQSvzXtP0fBjDhTwiZ27KUpMm1/tSGRDhxnFH33DBxv4foKvxnkvMc/T7Dyiv
nS1JFOK3lu+/9FJeeyAK5iwH7ULE13zUF1RMQypcwcAe2tGUlcI3OBsVSpaVehPWIgF+/LrCnFT5
Oprwb0Q/6eJwNDjQhbc3Xc9YjrnaxKRkusjCIJdZAPKkjUzchjxx9nfkZDfwJcGd5uhvk+GIb78D
sZ/os8GFKPOKCZ+9qFClCgVZv/pBkm/HeS7XRp1MFtCpduNupHvrgh22my03W3i3yNWcOfkWFlJ8
O3qyiUSc+cDzRsWYusvFbqsvZAWItH3F3EZVTCne9NHttjeAd30IFPwkT3+AxsatE+njChUHN99F
Qjz0AQYi8cxYcZHvTNfN5/ENiV3stVOGUVIGucFUpl6X5B1EU/OnlDcPuTcOKrqTPqh1rrhjYAW5
h+w0pRxv2gcThyeWrM/iuYXd12JtfPWW9ABYX8QT8o8uPJ0tBJAvsllE+ykTtRgRIWVcZq18t9Tw
2nRtmsJYZbp6X8fUzvj5JRdoK4gRkocqe2YkH6X9f7gvLxO7hAAJI/zELuD0LhJRZfuYS8kDTh4n
Zd+S9k5klCfvNi6X2jYdOhY4JQIwT7NwJYilaoRORTK30FYKWaS3aox9sXmiF8GKOr9qOlNB5UBV
n9K5qy8IJMkJJZBpcSemU2RPlb7icLCrbn1M6hCX074c6Ur2FD+Uo5d1DbbCEDYnFsJzVciNoK5n
aJnrZ9L6uQ/Y3I8wVt87KsEK2PL7BFqQYbCQfLjbOsMRzOMSqgufJZc+4yid3Jbtwm7XZC+DlZpB
NPSxUtup91pb/nFXk1YInlzfokv558sokbss4vWSXJqAVj0P4EKz6bCH3kNgobfVdfCLifaDNFzU
tzABWM7QYfFi0dwfx6bK4FIY+XCmET0G0zH8FozrcnGblVaREA2ygcTSBeUGq3btQnFs5c+Mzj1g
8Xw1KG3QM0br6dYHglxrMh6FSd2Qi4rGLUPkwYOsguP76LziiBZYbrsaePWZIrR6fyAMnvn4yVk1
MgJoCOcHTZvEy4BZQy5i/FG5z/Fcquhfp3PYfdRW6H8gXIICy65gV+4Gm5960ktOtOoMkK+YL08M
n7hGBa4k4VWwbswuzsMb43e6T+F1mzU5/dw0qXw0b6aC2rebTKhX2zh2fpBhMl4UjxRYtVFZFVsC
sPYAAN3DxMghF8eQRcbDFrk1V5pGPx5sAB8fp2hAdFKhy/BFo7FZclhIL9UP6AUwvJ9gmxksnjc6
48+8D4WWJedtzldwdffF6s5kkBRZ7Qe7d/9BX+CJ42fT+3vXgVbIUX3IU5SptdzFV6fpHWqYkrDn
J6JGvpB/7ysacyT2Tw5NM9ahT6y3MpyUQE5AUFbH7wEu08lZpXVYw/hC5liZeH/jDyeSV59wcE6E
WvO0BeAPq+klN085GBcEWcJ2Y8sLdSUTqK2lpQNXLJkDCv8yhm/rQrBU3SRNOvM2jPL23MusFSNg
y1SQKrK3hihjWYI3hRIPofXaLJ4tfdLkNwYixr+J1CKWzR+tug2YDlSHjmEC88WCFEuRXg7vHmIJ
+V/GtYFMb6cK7WnrDAxBPTWSUXvQ3dBLL6l3hiip1y4kB30w1br71lcpVKKSXBRyvU+mkrvHo7p8
yE7xcQzpIo/Xk5qlcXkL8ffqD0SIDIP2m/H4req3wuiHMq+4PVs2H7MxIUlqHZdp++m6tWnGF8Ud
YfGl6lNQOQLlA6jYHA2J1ScNgKsbS6TTnG+iRHwIjifVkiB5LFry+HU1C/tZtHIxfrGU67qTUClB
e42CxULWCct64lYFCTejYQ6IwMj59zGrgPJhqSJSHjqTiPP5tNngRuNLco/ZvMeNWeqSsv8/CWrV
iN+Or1hc/NI8q7Dqq+sVZeLL/Fc3GnCRBYzWFifIh8Ustv+/SoRa3hIzzzhWcjXcQsziufTT2Ush
ErWF3bhmuY/n8o3A1+aeBvalqxec1wDI5FWZgBu6O9PTb8+b3a+37MGKB5dJJAyTMXfn3lqWalaQ
DAqrKO19/KQmssc74PigVQPlmcfF2D5ArwARbuC+OX7Rk5y3AR3zLxAPlIY00wFYfMWJiiYQMDeE
tpagipxj0SUwxFOr7cFrD1Sczno9nk6Z3eWWZhDFwVnEllhy+zhx0SENOh4Q3oxva8sOkPqBOe6C
hDVngKPXsXoWXtDY1qkRMrfv19BJxsahIvDy0qYN0iPoZOWMGcYgWy/daJGVM+sfYqQ7Lxg/NCiM
P39DTG109imLhGrNIxJxonGUKqbn760JkyCHM67HwtyscOYAjk1ZhSCkCK2O+AFoSM6Z39VEcoau
2ADxbLQdietDGOqFx6+2FGDtcx+ZyZ4TegH6pI3E5SrLC1DMweylNkIpvIGI4Omy6RSHDq725zf2
vpMA8owMEaTgdARV+esTzbeGcXKdxyY8Qaos45JXf5xW/SyC24arSUp5uCJckLjtZcYcJrp3Tm+y
Z7r9NUjDCYnaGLyGgj9SyJtZx4dj/J1NQ1jaiICbFd280PZvwSF4Cx7oNjC/sSxX9fTK3QOsJ4TP
qXnOSZPrEcLSuMSgV+xGVdFUsU96Zs84T6+OCkI3yACVqWGNEFTHIi/AFiQfIoZf09uWCVitFoBf
glGqHl9bXkp317lm+5Sl8mc5iX9TWVeBZPHbxsKU0gZjuoeYhX/RL+G1dF0RNmmSlnPUyCWY/5Ws
O2GTxsnnR9znvrjn3ZYlo8c9mdSuwX5Wq05+a78wPjMwFxQbM4c76WyzkEmLF2oCtktyygKH0eKD
+n1ZzoSlv7CK8Qhv5cY+Y9KQ1QOGtK4UuGbMP2dsqGBSQ6gz3I8azF3E9hd6WXMJD6COmz+2nmTN
aa18+LL6DZkHV0Czb1pAyskkbwYb8ZhPYChenjvTFQImF3td5YW4Isgxx1mVKAU48bkWso7s8xZ1
IYaazxk59HsJVQiwKKpqBrUqFfXHGvkFBdhWPJFi+q8zsEqZtBPdzPNOnc4ckz4r9DOKwC0h9v+4
K7+0LL2/BivkkQ+2rFvqSWBGpm5QsmvRXa5vyYy3O0CRj8as25YknTfF+lAFM2eMygqpY/mjj48z
TX7MbPQSVTQCcxgxJI2Ip3GbORIo/AgLue07UHp9eEjI5VsmKkU66krmlzgsSFXMIjNB70PEfirp
XOjVEzJCLklue7r3tljlU2nwjbyflcCaHa0lptOELjQ/nT2hNCzjxumjFbPFxzcQtLu3HxdDF1UE
32NORXdQgyx1XbAAFCqLyLKNTmhpH3gYBMyOIj05gtn9ntKDwQrLITA1b10TLfM2pbgDfs9gx1bX
Z9tEmmOWUWCEVdSP+rs5eqP1qREoGweeeLVYHnB1oJ2gGIBhaeO87IxY09anSTmuzEV+nN4xusDt
H0sfg3zDqI9vVDHwu0Ctr8177jz6S8rR/5pTvd4718yog60Ey12RZzVtK8zGtJPCHOe8IsYo6FQe
rqpJWzAa8pgrZoq4/CU8606vxFWwHYFSrX02cjej0GXwSRjcMJYvf5MsQkV/pmoDaVYexwZ13bvH
J6Uf4ANy8cvsSxccz4Oj+GIMk/SaMuvJIu7nRNNZbwka3J9yoVSE/jdbVRRjt30rPLo539KBAh/G
xcAGaJ0elVgcV8MfNcHg4RI6AnxSdyCxmVCcnbeDlPwm1i7Ay0WkPkTZPL5HnbsBRL0z9ffhKoad
mcF8OS/zI8Z8e2rQeEFuLjSzCqpsGAHnUXeI6w2me1dY39TTq3Fk6P4NRwpcT6cPZseZ6pBumPZ5
lFCh62vsFvb2hC88txnvaqv97aCUPQ4u2OeKdeC7VZB/HaytmefwL188yj5+TUdQXBwC3KXvXQO3
YWYXF1WaBWjIukoTGIYb7ONp67pI3uHnVizisG+a+XDcnG3VqkkOBDvBhcg5+ZkwK4iH9Ysotsi5
Lki5EyXLFSjbpXX34z6Glb643qccTCYic0YXBlaCissoB+z4lacmE3n+riai6yrzEg3k7uc5Ythl
W5ib+Tb0dGtSwE1inlWF4x3+C5Ir/NcCUobvu9mYEGhQRFBoi77bcB+JRe22XthpvWBZgTfy6Lv1
9T+BXWeadLnppwwbLNpMlkxyvpD+3TTxj87LE/MwMdCiQywJ8yDxHgONdzUeYrqd7dNTVe9+WWYE
MD3V9mAhrkHkp6GOrS2NoRRuyr3VzwXPBoBgWrWQiKEPtXQxYrNJwCe4wLrb0xJHpZtzfEF9rLVJ
/GLynEM7Eu2I03EWWzaEb3p5q1GHL9HF3fHFbyIW0xzdZhMReo399Aj+ZN7fnGpgRWce98j8PJ+a
vemQjtiATuxMsnR+9J9iqj1dwrVQkNQ+R0tUo/iyAROHQw9BfWbEi89keS/KmQBerg+yJQbivgIB
y9CNFVFE4tXhL4IjfLyfbuZMMm+8G8lTCJGT9g5UTnbZx7+tFwewAlh33NqANqXds53BZOWzPuel
3a++ObZsp74F25sNDPLRcaI06XRMBfpxppCoV4Xr1EAV+HqcdWlBYM1CK2wrFJNTkVdx+MCkeZcc
mnQo11IYPp2o42uxQfbX6yZk/02GRguyf374nfM+sb4q4bdJ77LRKS7/ICD28XUgG+o2Wk1Adeus
g4vN5Bf5LNSDjUIJI/MFjynYvbxsugwFKCUPb6x6IDprhWBchXI1sE7v/5UoyYZ+VqoqGzBKllfS
dnDujDmM1ZuQh49RTBjDNEywS2plB9uYkBc6wDV4KD5knygXAqR95QfCsWsg4tZDXkGZxr7x5iCP
87XoPH0zi9IEp5WhScKH8cO77UPjEeTM5+TxEs8Wz2LTE2uNsVVEpz0pOrdIDv6YZvwcw0It5YVh
sI/bueH5OtSkt4sKDj3vAwoUfmLS7drwlCy+xUFAsV8tDXFnBzVOkyELjxXvI+6GMUaY/Aak2Bcd
Nk932Y13ZkWWKGEp9Mjg0rhwLlJC0IturaAzQa/d1iSddp2DqGHfy8TeLdVZGUgXayfCKsbViq3c
8GS6FygFoNIw+PxPT6cwW3nU6AYg7ieNIV8p/T0Jby2/tHukaiebJchcGDb+UI0FRZ/I3hvuIepb
Z8gc5+41G69M+W3raVSjMjc9/vKBieLWiuQ/TAHjSTjxkAAqZHJre2NaY21q8rmKQ2kuvpJT0e24
K0D70QI/M/00GB6vnIgrgESY569vpBy2L/VVTrgyG9FzUAmHI6YeaaEMDCDOJru+02tBiOEfmtPD
yCYtO9ZA3OiDEbvBrJ2rywDURhkFaRg91tXjW+7AZz69pA4YOhtBtnlTF9cxaiuvuropYfNpq/uS
VpIk3zrmUhUo35IQ8oQHRhjP2z7H48esGTrVRVHtMJvWo+Vh81VoUXxyoioyak3lQP4TfMtF0o8S
xsGklu4znaVE2kp3FKqLzEE+PNp3VnkGHXDezLAHO8xetyXcXq2YtHG4T1wxz6ILAAkVtXmHuBQX
xWLGV9WWmiszG8VcTXjl1wShaKQaSIP5C1JsmS/BE2lSWJOFaCgL1TtvaFidf7Fd+WmBMvpCPItJ
Dca60hZ8QdaM6IfmBwAoqQsBqv1495GhA9z3qFkaMuVIkAXmCwe6sS2bpgRCxGVig2bR8uQ/fSPD
QAQxm9UdMphF+qG/Qb/0MCStmG/eXAwxZpF7YS1eAJoW/bViSKRMBTxyBU3P7ihHwDoiajTt5ziz
9t5menvGnFgo/G04USznctHM4688aCS8OlWyw2OOlT2JCWKQaWiPbxPHNZK7aSNxxqn1BMnsKYtA
F8CJoNhopUzFqS6J02n4yRYwWbdq8dV/n7GqpLgCz9EJM/7sirJSBGQK+5xCT5fLV3GhunpA2KIW
GKZt0HxDkZ39v9e1CaNmtMJrBMc9rAHqNb0hh+6LnISgPlRhhq0biEeXZonNkPH5n4jipS72mw2d
55capM1AlIA0T/8FQngPLBHaDdn4JPStV86T2NN+OuqbM9Hljwo5psPF1N03Rd/guTAt3Bdy2dKM
2cuUWTwgHVox7LGKxDzRkT/FyefXFZrUNKS4HVpZy6zcewbHTok7UUPiiAWitxPqFzM74u4pq78A
Aq9Y4vnkTX1SMt6Z0yehBZ3jVrJ4T+9iiJOVMDh2LvPRH596A4d8O8z6TghpUb7R60yV+whkRtwL
Vy0SGuIumWbaELcmq26D6N57rkgU74LE3tHgtx2IrwF+17pFtpWsVdESagftltJUvD5dVU9mqBoA
WyDPY+rzmTi85fP93HgMuZ4JYFyqTUK7O81vxxfv+GuVtsHtEnRfm9svDImgB/o1iT8Lg3VvRBUb
Ca6FTb/ecBXLvuisialcSOhQyPj0H/A/Ix3cE8uW84PLfv2WBqGfZ6rOUm7x7i9NhK4AByQHsWIw
C4BU926kaEvg6NsjXanYS3OAgAK44CxFyMtBIIiNmgqO81ngy9d2zWLTORs6YpB933jKjTva3FvI
KWlINID4Aso65jmaZMnRxt85TcZwDZV1B9uUMNC5S+8vV2FOSYilprUgD0SiRP43L62sfzNweCoo
xLYI72UR9fcG3TIEaMo4kUn38sK5WzYsELK8j9F3y8G7hUAcCPzp6a9NbAQcMgLP0PZk+U7vMQCT
a79V/UV0wZkda64J9x5Ij/Tzqv+r2DExcCRDgenZOuSclOUqMtg5u4Rptc1TmOVdi1oikHmAFnnd
Ta569SxipS4aX4UTjIwcr8yQGGJHuRvYldf8zzP1J1cEFqCbJ57Eu2ZVmh/PibRg6p30I+5fBQlj
WHgqsFQ4GxGarXZkBNcKf+8SDgyfEj6ayoqRQf9PvHc9bIgt61Yvku4Bs/9ejyVAIQPB8qWGR4B5
fp9fHjkwWmT18yG3IBE4x0yfvjHoxBTszA/YN6GAttiMLAzg+AqsyuA81QsBKmL1zaKzumZsPrl/
ifKq6XyRiTmEBmkjAa3dwDUDEYtpyQqJfkjTa52PM6g7flNQViFXTCLF3w3Yvz4YOiaVDKMpEOqn
EcTKf23mOvQcS8n3cPd6+3wiT+cWT4DO1fyEZt/x6BMDV1ElUUMbu0kTNJkRRfoT2V27jkVi54Kf
iuLXhZfotSNfcrd/l+MUhL8NPCDUwthxZAtoRMfgwffesxVjbn4Q7NBByJaH8uYw0wrGCsnTAE//
hhmTmqeHZOAjKERdAwDDz/I1dqkKGA37sB4gZQm4uQwR/1TPNWsmuDo6w/eGxz07whdDA5CKW0oj
WZAYNe5aFMpNTK9uYpVolNeOoyTpDlxZcm/iVbQPgl2lkTMBlGGEtk5liDYSyCLzAGo8cc/XXg4F
Km7mI8dzSD9kcv+jRlcRChMCCw1kvoci710nUxqhMx9ToJSQexSYaiHRk1bqKKMasnyxtrzTvgYy
i5N6NAA10WJ3PPSAB6RVYFcCoCtAKDa2JqnaHyCPOuF+zEkdQj5DFuaduj4W3sxhaoZ66McidMzz
xy4/1ooR95FTE54JRZian2D44LzA7JPI5kEVyThUvOyp8YiiH3i88b1GT+VkV/qmAILFlS6swSvW
ctDK6oKVnJXB7qGmkZ2b0n7BW0Kjhl5FiE5M5ck2JH4bV8IbRcmCbJzi83xvcXpdoyzA+FoWPy41
2cJEkgkEAvGGGuxTeGCgXe5oJGqwFEINjaMFGKx/4j07sCrkfoGD3IQNEPNcjvdIg9DSntShez/Z
2zZrYY0glMDYljxdUINRo2eLrKgUaBV3PhonZDUhPEHkW1GD/O6IKDUKL02bCPAjCPx6iZNIAD2y
ZTFoS2pLclQzvq1CmK0brJmHk83+bVJE0zppUoGg16ueGOvjzSpRYfFnahuZ8P+NSQbmwKsk3TUj
yoj+eOMaOHl1hizRbh4A4VuAP3+PlcsZ7ppY+ZmxRAeijSYuQqVQEueHyrmEiZjuwnqIkPM+am3O
miMrp1qYGYbdZfY+cihXfiYH0I1//GGc3Mr0aStyaeJ8cUW6/F2B21t6HO/NEoQVhxm0Q34ijLyt
Ug1mnezYi1QD4cVHvzrqmjjR4Ed6PEgsdfut+FtU8tRdSDjr0NrxyF8iae4j/Z1YaK2DbfFOAQZ+
NFBO+9Vm+Ooi6/rXFLzqKlbtslVZ3GvT+zUeuHJ9Y28SYc5PCV4ByvJNUhhjAilLrm2BvsQaHYPk
XpisRK6PDQKC2yPTOJ9PQT0M9sQEMM0k6NNYXEN5uVi4ZCS5VuPhHHUu3MsFrTupYRS/6tJJtTwN
fG1w3FVihw2ECNlTyikhGv15/iMmfo/VJUIrai7iwtZ+3jVHrgX8/OP4YA72vPcCWOGfEzNni11v
ODjq0Ijt8mUqu4pd4C9AFcecr1pZbfYS2zSrxqwE2cr8nGyj14syGdNC4x0tYyRtY8d1z0WdrfGl
AKdFZWp0t5Mtu8kK7kpI+kB3tyvKUghyGsK3c8KePF3KxC1Dyx+r03zqRClpiZ9SIDOIuMLY0vh1
tMkn9EUB/mFm9xAZraAGQr+g+FxKRE2QImYiQLjTI5DJha41Zg2voNclvCTz4dd57+0wWBzy9Q56
fX09VfJ6e845CuxKBNHr+H5yD2n704JWlMrYHcSYIhZ1jbfwhts1XgVDgdlTH8QdDjJzV3kK3XTD
0GbQoLX399qWaOtpkA8fX42bKG/s6+Ifk1+jUEAhym3Pj0og4uzjylnKrHLWsQMck3I/HLI4y318
07ny/5DGAzSDxsdXOSdIW0EFwjSJtIiJEkhptxhu4Hmkllx+W1GIRz0ts9AaCZOfBjK9jcY8/qaf
yHF97A1hsxba3LDp53H6qMGYx1pGmPr3cXEIrUtKZ+TBlHZslLSLGeTkrIuqMLnw3xLTZLfNqDL6
yayjeaHTgsFUAwJEyownVLcZNhtkyMi2lE2cV0waXhcu/SKfr39F88pBM3eaSrRGZYhyVfoy5Ekl
8IqFjb6hhivZwpfqcl99Db4Z3FUN7K7PjwAw1CUBNVYZ0i6HQAlWPZNhCQjLySTyrpFiFGHNaO5B
0AOUbsQ5ZBHt7hNMhac3M582W/Ogiy/Ei0s6RAiV6J4Cse5z95Bb2bHknCBGtEYSaThIFA/4rAH3
JPcp8XZD07XAb/cGaCLo7SJbRZcm+cWmtwzPvMd3Olw5S++9Ob15eYaSJN5N2C6iU024MGVnuqGQ
82r6nRbZnCxwxPi9SowgMBv8F7fLwozFV0t0RcJVIVgMOZMtZiyx9bFRfzC5nfII7jOj5yvUKPQt
l3kyv7RcXkKhTw1ooTWQlqQhAyDmzIStvf4iY3MVDOdPhcFTq0YubyZ2CAGBQAywIKCpQRz4muUK
/m8mKS5OiGCPji1mSA2sW+NCD7ahZKGE3D13LK2Fu7yFbTNDU1I94hQ8j1neX97GZ3n1cZDwjHDB
Kg3qTpwW+M9XgHQn/NsGQXlb4gd6V2Vy53xKP3zVjyMtnlSYdHDqKXKEY0U5/UHq0IN5hrPxjJ1/
THJy7tHwrqrH8rYfgZPXq8Hbtea9k5m+cOwqKNwKGE4l+Rj7Z2ALNDZXMbM4v/tYGWUUhGVQGLhR
7o94M+w+ecPLU/wuYBP2J+qWKrGBtubCdcEgAdKoYq/hcgcWK0YfJsLD2EclNU3Jt6HO6SToMEyp
EmXFAUqZLdHfzbO6xx3/lsrhJixNG+b16YDQBAoSEg2BrbbEOId9NySZ1bKOJOd1XYfhbDHjfIGn
9vdTwbX64kGZ5LpxsaWw+FoP95nmJ91xXfmNv7QtZx8PCccEgFjKew3YbXBV7uiKgfTETCPgnXfP
zveL0z1StQnHkHEKduXE9iR9d4w85SQ3lHxq83E+JFLZ7JaWiN6jgG0WcWk+HJvOi2wxHIqaebQo
U/9r/5XBvEr3QVkKb2Kw53fUQJgxo5RMpykCCRWaDNHwGul0IXFVHj7Uo5GMS20CWQw6q6lXydKE
U/K9ox25iaM5vIPz/Pdr2i5IP+3WPgBK51fd+9XSOHwlYngBqw1G594BKSQikY9p+tPfE35x7r3k
GyOOtLYBkpqcXs0gpaKWv/yBEnpk8qniL2JaBxNRnrfi+RNd768WUGvLHaqyGCtUBapF+eFykllY
PT3pCMMfJ1ZldSrMkd4+fLcvd2cocSSegx6LxT4c7UnFOAsX4pm2UkT6egeihb4l8mD3vqlOwRDj
JvW6asm3OOc80kaxigSYSfAlHjeejbiIfcM++kiYhyoqpdnK9Wgqvjfc/2H6BBZbYoKOtIQDvAA8
iKeU+WwFwU4W2zW6+KqDUIRUGMtJ2oB+WxOYxT3WUxml9aGA/Q2ElV8sdK99Fg1fvNaLko+9lK0Z
bXVubF6Gh0SWlSdkIPGA5xV8RoD10bqm3nDlUHyny4tv/KWfhR2MZfD82h0WNgGRakEqNszcP1Xm
8pkKYBpJ5Zs4+YumWwUNw05Oc81ohDa01ref1JW34Q21NGuPTSquHPZi9ig0NruXse808/Wt1qlQ
iuWn0Zo6ZoQavubQoXQ1fVu4WgzipBNmQtKw9eAoBL3rxZgHgmsrBZoRCcZHVhdIwE014uNTWBL7
ugx4/Hx5S9q+5Yq27oXBSBHrB4hVoa7Jm1aHhOazwoDWM57XXKsWpbovAh6y9WRRrmu1h5Kl/mkt
cAi5GJRLmlMxYPpxe6ycYOUFAF6xki4cHP3b4A+zgkABJMWWDG6Iac9Y5MiSLYXYuwrjy0kFwOkx
L5a4bZ4Ygii92crh3oditzswOa8HjX/i83Qk84QITwJptWSKBBV1w5MljXrxJYubUPYawXm/hInd
1qLNZS2SOC5saOz2MP7xx2Cq3CCzSoWO0Ig7EvqvoQO4Wt43LCnKb7F47vSJ7VwYVCm4OI+2XcPe
yw0wVzzYjdtsHe97fJZRcc/JHUoYttt2M6T73uhzd3eaIoZL+GWQQB0qD2QStmyuXZao/nBmPN8Y
rEcBhiFhABr5NNwpofoSmocUKTDDEVWS8da6TeEas4Gefhcddg66GMr80Flscl7ukUFCQX/Azzk6
Mb+JNo9dYd/svQt7OMTa00U3XCo2sc37cF5V82cLhkSBHIE8K7BlVko6oDMW0MWfivJ/vYyXncg0
W7gMB1yytCcQwQXXR1oDOh28vanPkJVmLrPcuOe8UUY/BlVOVlIMn0J/8Gj2lk740mU+2S31X9EQ
9+tL6Rm/tFs/eue3LzmnuQ+PfcaqIAbZLbqPvD/K19UVakJsQUwLi6aJ6DxLG3d9Eke+YXu3/Ppj
sLUFNJJ+FjqeAybZgcvwf/sKBhOTpGQ+4tvZbEQyWHgzGGdWyqNP0rJpllQyvgKzQ67CESvEuB98
a6AMxYXM6mAzZn74dC30jOh4SjtD7nJCAhs8l/4YejYOb2wDPkvfahqSlOEMjtL1OxP4d590D7CT
wOyBEISFX+yHQpEu/eoeWUGDKEjTXsBMTj3f+tkGVObW3MEev8ITHzE2+uNZxd0J706WzHA++4Gv
ldy/4uEgvvFwVWC6FlGUHSf65xwXhXw9+VtakRR/SKp+pZ1IU/CHxF5yIXLLxOCzH3BVKerVKGrC
TYBBkz7E6y8o+VvsYNA1KUCBokgag1omKNDSHLEbbuzFBVFAyqMzWsGbA+MtH+qkxCQBhOkGUwFj
DmD1SsPevnofVayozqBaFDfLSc3nstKmOl1OGtjTh1+7IdASEDjtxZ0ggX+bYjAUMWUmF/C2KnYT
cZuhF7m4EabRwD6WnwBAZ/93KQwFiN2vfR+Zt87dhXvJNUgwcHlrM315T+IbNldIgLCkL5PJFqAH
D9agqWWN1VmMDwC2w9ZJdCfkg1C/fAlIWs2vWzM0cOPmGk9BRaCq1SwYEzxMB5G/PGnZp2p5IuOP
57syy5ZdDBL1Qfe3a2a1SGlwZggj3R6pQ3sZBXLOl3/YbtLgam9aAP+BDA4Sq3IPTzrQO/oOAmpi
+irur++BRWP7oyuH+IfGInoiyFG9XXUqaAF8yGbeBsa0CK9g9Sa3mO/G9XcniQjHrKuN7etiZ+GE
BDjXW5wxkzCnciMli7sU7waspCeTahxzTFiYfsKitkAwx7+JH1fzC/mfTArPq3D040ZkgXt1OsBK
MREpIXPB7QZue9A7IgQAin16eNy7FQXrXEbC18LAAcKTJRnSVtbAvSCJAufhv/v1O949ggVtTMIp
ef93CtBID8+5XuptfTU3MG8eHZ6Wb6CFn+wXlDOZKcq+3Q3vbKHqdLVBBNT+OIuUVD2Xx2TV/LtF
ycfMb0A2QF7BaAADGRRSBZSGov96I8j4szt8oRuHU4EueuXAlDkSFXvQhIZyQgjKR2nG8uea/lGS
9wMc5QtS0ohtn4OdOSlGXyVLQoB/rvpxYJbrPNdZTad2+B+1G37dhfza6dMdGRvrpEzxXHH/M1ht
vbhWpZODsybZmxsYsH8l+UKvaM/xVlWuJG4q1CKG0v4fVcSNcqvXPaDHkR1jX88QOpnGLApvz+x8
rIh8VwIQbNuiwru6LByrC5hV1tcWtFtV6smnVNWze1576SxowRysVEx8RLQwaZkFUppoI+L1lkGP
v9GebmA2XMNV+7pxdr81IxOWkBdLYKkI3hwEeot7s3MA0KNsN+unzY38xk07DShJ84RPlCTsd9S9
IjQ3+b21O7XnpijElyQsuIQkzJI0IPnCk4YYKqOTR3LuHLYqCvUO1RK+jEv3D6Hok3g+CXpAQMeX
LtBwKEo11mgk0bSg3wuEOerxjNBYSbyPF6S17faansT3n9j3xwg1c6/zxPGTtFFZDQXbCCBgXa6n
RGuYzZzsfrspFQXVQ1hHwTxO39nshuClBNSu9e7jEjiCF+F53iFfV9HM5RLtMWmXkJgzx6NhBcUE
R8uyfa/CerMz8H9W2egUlg4nMYF7TkcQ7y+EnCM+53G9URlwpOxplP8wgcgR2MgRJtl115iMBn9J
DGU8OB75dRIuGBoxHtrtUtzmNofHNgfIF4uk7G9ZQ5XuokMVoAPnOgcGX6fWsIsUrpT5+hW+yzgn
vfq3gRAuSfMDm80FF7QDV1W1iRjHJGExNCtogTXLR+GJaoIKhXEXjRJMwthn0ZiiBTZhiN6H7iRB
IfreBFbNU1jza9dDITxoY1zlQKdzgboKyIhjwVt1dvB7QGlfeM2kPnxTRaNjsaBE1v2Lf4abp7R2
4NfFjVD60TShXCdfZFg3ydprsO/1eduJrXTK7xo/7aWrsRWvWX3PvZZbG5St1kYIk8RzmolfPs4a
MrrL9kEul0U5d5I+8w99eKmpzF/heU4u6lMGVc37EvvRVeOhYR6srEpOavXrB74ApPP2utZ3L9bV
oZy1SqZntoMG62SVzOyWFqYdqYjWHs7ng/Xim4rGqhM1hhLhmNPtqTD/fmTL5lPX1E1bDytl35Pz
qGIlbgmF/zVMK3p7f1byE61iX25N1pUZGF2oydE4ymwL0jYFsLplNQYnzwdFpW+cpiaO1llhBOb1
BxYI3mbQY8UD9DPZJkUDrTiQo6bBJG6joehENS1oHbqr6df2EIXI8yhLBJe6o8dPKSDHvbrIM/cn
r4fANdTANwwtl3GCg7B5ES1qef+hfatvMYN84QoBYnufbNEkXPstU8xg2TRXmrzZ7yJW0clxts8p
ehVwpJ0u2txn99pC9vllwwuLcmSntNkB99Cdvy0yrGJDozI3I/HETRk9VwqvgQ4RlB7eNBnmX+hm
DZm9GYXKVV3xnXuEWr3HFBF3lbxwrWqhpqaWfLgfCP+qO1XV3IFWBhd7HvoJ1DY6ZA9kh9REVIEQ
GWeA+243b7545055jQgvAMVCAbe/ixM5Bdc9JDJxmSZzp5ys5XJ4g+dzEe7gKrWC/ndtdMLwsr2U
P87dUCyzZO6hCNO/wMCD0wvd6DBmSzBlD3LMAncUeUPbBCufPaEt+nQarYIuZYjw4bnyFLM5ZvBJ
6TxtNIUfuvGF8DVyCpNXjp0v5Pp3oosYY2XC52Fj6gYMnTe+EFha9ZDvjf+y8toMFPOhFA79WnfA
wH2Hl1Xuoq+J+gWnMJglMUx57grxpOsalDqCEFPkx8/mX8NVQ2PXyOCZv4ozGA7YW1OLQxiT+NsU
CnmN1W0wMeSXZMCzKLSJ430Q4s0/gT6HOT2Qfd8UK33JRPEnzvdS7awJ01BMPw84Fs8NDf4Eafgj
hDvCmiB60owV71H7j3ydpu1uGjw6mMFFrQ285bLnsrDwTVKAyusnwZ8HV2D2B4uQgxcHfeFjBXQC
+bYmRbAjsXX+kNAm4OfEOvUo517vgImNUC3KfuIPM0JNA+C6l14dk8OSE5oXISb2apCOTZe+LAuu
njwBBUX/1oRLi1UguNwDzFjrIGEqQP3SwMDlyiBA9oe2TVI0A8ytQGFnOV80T+u4AqTfksGqWfm0
mT6Bj4nKcXYypBoV1WsYr2dyVyn3+AhVLgz/pdXKv+scCYxN9xLlzzJne7B6eeHrQ0bhoBudP8AD
xrC0gAx6W9Ys3bU9j6lrmSkKgGZSB+BdDv2Lw0H7pHUHWg4ytdXcxk/f7gkWizRLHgpxKM+qSLVA
oYrv4/iFqlapq7Zd3iaVc5Pku0/Bqj1CTSb/VWBs1oePFxOpfw5GMNhBrDEsUcLEU3rnkO01su8v
+STnzVnZYvVV47bM0ym1zxvN1l2hSaxdoeqeUNacKjHdvBY9kXYAtrUx9f9VzNTrak2PhDj2iJle
l2FY14zNNNpDGQQeWjGc4v0JFBlQDJbqbV2NHwD24MH4f1YFe+uflSs5X1zgUDuE9uQ6H2dL+bQA
CP/PcyLOMk7+8Gw4CXrStWeqihNs+UFlQ+CmDXYi8N4veLo32feoAyE3Ue896W+HQ4cZcIVNH9xy
O4Vkiduvn1pAV45NKUMq6QzsE5J/uUlt2KU3iFgnBd0Se6JRij1Urk95Xn6eSgTPmHvaerfsq7sG
2p5bn7NJal+u6PXuPRs68fn8G2Y594UyFmuSGuNVa/kUY/OZ0G164juz1Ut773KL5ddHBPXOXahg
XIjjMIQi744Br4xjBWJV9bPMc4zF208PDnguXyoImnuxRUOFNbdhEy2r70MhcNho/69gCMTEhEB0
mwR/jZt41phN9JETsBnmQ1L0YdU8MYsUUvt3/DgkwG1KGF4vlTFCDaMTn1+aemEGvNgPursCiXuk
ZLEq7fm5Nzj9+TRwCo1deeZdX5EJqam5Nt/c8xFeFWlhgGPMhac8hCUE9PGNUEJcyhkIVyMYeGN7
c9dTNHKFDohV/Zjq2Uuz6KuPhVNnlSNSZNNFM+jRMvMrNSyj7hXcr70gABUIXmn/9IHkB7X+QCKz
wYD4T/fPPwiLMqC12/2raU/eO68uFC+2onT50giRQqDZMb8vX9HDNn2Ad3shiXQO6zV7lAWiOwxx
XLa5WtewUQSyefFt1qXXeeIGb6U5BW8gcj+VkStp/mA8qq+Zi+5P/4MqMX4D3whyn1L6uA+MedXk
xHwTKW4wX2x7Duw5XSBAa+aoclLK/bxiP5nzFvXehVfw4st69LOrTC73ELF/VvhXQKYqhVTIefEK
7WtqbCu+8AGMH1+zU3j6+z9KYLwcMiibFbVAC0u2ixpN/acLakO5ZmdcDWqxYgg+WNcV3Kgl6acr
3jGEQEea/gOsK+Lrj57Yg7l8XdHfeYDvK0o2HfSBow29hfNDDD7G3nwar2KFs2qDvoQXYcUQB1lT
cvGIzpdWV8amimp+HkEmd0qLSpo6lBfgAKKhGEImrQjeH4cIGz9owvzkdVgOZHS2Xgf2FY9mZ9ie
E2QgRnsSAwcWOg34gNy9/UzqrfGWljpq3gdXWL6oqbIprLjI/5KwHN3PA2pcSSMf1ttaujb1do2L
NebUQ7VVpXRGQYcI2KPERKQsxm2ZKPFlsESk9Pdy2vfH1Mh44thV2WRFQgRHwQRhz/+BKQeiFuFI
zfXvrisxi3bd9HtffWFA/OjkE70DutiOUCUOLPYe3SPHhLbfiGIUU29yKdFn1rJBT/Uta7CyBxUA
EUUPGT2DEAZBSnJOsXqU4biZ0/2NZ9HtNHm8mevvcO22o9t5lPUygBKlPbSm5J7YmtoueyC6X5t6
7veWZtsdW13voDiM9tTQ0ZWvbB/ebJwEo77dfuWuMq9pntFkQD3RGG5petr34NflXugzOa/qvqyC
xfeiY+Xf+5GqQMSpJaKlKbG/YKkfJYktm0yiCSNlyEho3yDVwDJXbxoIog7YplAKutq9HFNYK6tl
4Y2B5efXSf2k3N37Np1G9za01MRCNtVleJ7134jon9vGyXvatverrGzh3kLorwyQ2NWJ9utp7YvC
LDYRY4RuA5bkdGcKhCf92QCn/Lm544L/D+OckbjuWh6WiQr3bs4haKeWH59CZ4GFzEmCDVTk1b+E
BOLF46AGaonS/WR6jzcigDNVcVQ1B4Y6L3qUvJ9HC/gv/wwqGBXEOp5NmRzvjPPvp5gsLI8hflXS
DpYQQ8iiiXhdyQpeT4yduQ788MZJ0NRNc/U663coTQLoQbSpGjmDI6dZGwwbrK+8E8oQPjjELWv9
3h7EEByr7c8IIA/AwrML91q4K2Nbh/efVxOwawtk5uaDeyXGNMMmGYdq+ZlprRyB/GGppXuv7eI5
Hpz0e1DtHtduDzZJsayan0AbsRxZ3Clvn8msKr3c/3m/YU7RNqormNaQbrHqFSOmLlERS8CKm9+D
z5dTcMpdu05GGBMgcpe5TJK96DTH9kJVqNFZOWlsH4EBgZmFIXiZiJorYmBpUCWcrivMOZ6iF6Mf
OQSkUBBrFemo9KS8KUAUvZ8RZxxHqwDaFX4cfXbSC8gNg4QA/mt2elKufQMqD2DUetspN5/Pw8zv
78etNYidNA3OYqVNcIaQB/Hod9+vipKR3F1zsLXDP8vWljmil82Sh9Yw8QQWGQWdMIrfKL2n/lYE
H/omruWVorgxO8CzHdr3oYWF05oBV1el0ZslD5Wh3cUmHAPIx2+79skGIWbn4oJMbdBI8pf9CM/n
jQcVMBHLKhgqqcEGqyBzwDk8ucO7hco8LOwW4LUOX0dNkcja5U8orv6x5N0ocwMUkWK6rAt5sn9Q
uH+JuliS5qGQpuWblmLPCp+LBHsDMXgueuJW77n1OuV0OsWnqjnf5z9m6Ck2mPboWakOYyMQJmBY
sefA+oyAZBZBo2+m+wh10LR80+jwaLQWGXHRbHR81Z/MAjvEXvyBmgpI4Tq/QdOzPx4GuE1Mfn9p
Vujkh7qf5fRL5iZeYLGUY47GQvs5GGdasRU97GViOzuvtDtomlZ67kc182TzqbSxg/nJh0YSLuPd
Su8NRrJ2sEnB7IdTk2gr2yhOTRNlnm2BvilCJk4jlQwTmKkG9Fb3NlmlJ2CDhzyYJ0RjqaDqtMjR
nOBxK+FPskQCjTJ1Clw3mgj6rLZy1saKCsGH4r0kEbkO2udYiT/vRIbtAQXuCPgFBjbNaUMOhviw
DYCxq9w7wMT4IMUdQ9/iW3+s+jP6JYlkM0lLGVhM52m1+M6olyV2aj0pB4TlNoXa3vFG+9d8ozRr
bKc2i38KOR5H8V9NQMHyyFvZ1EUC2Qj7x47DjfOtBdA3A6x7uox/Jg3y12cVmKJSYafTrLAe0iyM
yKZpwer+PKqUWAevkRfXXCj9UnAyD+2cDC2OandCd0WK4UPMkBSCNg+KRehfSEQBTH+vR5Ak1Go0
8qK4FFy0JeJ3kroQ16ruXSeLmWexd2LMDVKIDn6tqHTNewOyXXEJet6R+Mkj7OJZ4HUdN3IH5XX2
2OhM3RuC8a/Yf07sNzkTkz+YnYzCUk+3TlSnymiH5uIkDM0u4t2XCVD8sJOkLoU5UG0k2yFEb12u
wQYwVWX253/S2/8NXJW7sjdnOVdda/tib+bIA3ovqDVQ19Nj0Id+3Sd0A1wUk8GXsG684sjR0ieR
mc+I8mCTfKJtBu9+mPppNNzWNQLFWif6SaVYyBXZStKzsXt9lptBojkdYeNHL31Sbo5Sd/viSf0q
CJhzDwHnpRd7IQCme+oI+n0yFlkLv5cX7ZWdlU3czOD2Lqyo87sEa+yOjarGwNdqoyDdbLnImzgG
ZwxB/c8F78srpvoBLijZprOwvQ/3Z7xQuKMXfqR+b+M7XPaKPa2YSByLilUGdS8t9Exng/ItALm4
PhlTBH2Vc8uxjNLXOGO40mtEXfGOHqOyBCsM/c7lWYx9SnNHQ9ZHc78KRBJjLucQLUAYKYsuiNcS
xWMFG0XxkWeYueAKfF8l0GEaip9pdvy8GdQvCOdd8YCNOgyNfMYvhyRVz35+kjHKKG0Yae6HxRT6
T5dq00kDCNUr9atbvKH3R8QDXi/swy5qcDdqQFwyURGrm0y4Nr4HCW24/2aUyOmA2kXRjiGoWkkM
+y8j23uq+kbVDZtT8B8aNjACITCVUrpCQWNuvq8DEzTx+knzAP/Kn9foNPxOngN2vpeEnFB2EQwP
djQolD68MPSxaY7QIB70WTJf5eRsXvt8LDA7lGiqYvFQ8msooKmgf4SxQzMenIq/7X+htM+urPKC
3NnoCSKvcqk39x8edM9L4Z3srAcn+wmDr/mu6Nt6Ea40zs/rHTBjeXZdf5uIRiIaxCMRcnXBwL1W
4bVNzte4CeKSsgDqPcmFSY44GdQFJgir/CEq7wZgChAHxGnTW9z/gVkAd16z4s0PDqaXVvvwhmbb
AbiuffgK6WGZ5XK+LKDtSYdLklm3tw0EBYLJOkievySqZCkjbwFVyjWd7GXh6TKIvb1fLw+y5aZX
TJsQttl3tg3K3MtPCkY9nG+TRi0xWPPzJZi0ZJb+cYygxuzXKe1htCV1pk1Lwifh9SSdC9ZtqpSX
vuCMG+JJlqveH/g/tM4Xq/iBsgGsrAyw12GAUdfJd0KmbYjYSC0B4zCmOkyg0hsTD+Pypz/1rc8l
nU9py3fgGeidTc8uEa+8yfxkEdZXZvKhL+YDDm2xZVXMSd7we5B7/W1DxLSOw2ZBH794KCqS/pgA
0gK1v9BHTYlSxLjMCtpamJGM6FcpkPVmUw0EXhl6UAdF/u1dkmQ+OcNlFFuBzz71hbEJsWblq8IJ
e2tM/Z9ufWcq6PuQkszr95VREA5LzgIDy8/l7XEVX/vD5syD4OoEw7j64jiBB0Gz1NCzTId6l5V3
v5VY+tedXSIaqJB727Bxfnv3XoDpDP8lc1Ys54zdc9A7slcFa5VVBVLcVHv9TtN/zti5uejToVxS
8TzhTnUQlyo/w4pN8W2DFdFqCW0Re+Icr3YCdziScY+sRMvQyjfeW549wNpKhpe7NGj0y+Obbfc6
svNbN3ig4OF0u6n6CixaiMMxeAGVHSb4l+/KkSWohUq8Lu0IvOWO0LHkeX2jqdNQKeb5jE355eSR
HwqDaWl07m3Ezuz1Tj6OobqDAAurI2Ji9IFIqj5Vm+kumUXiUtP7pNk/nsrBgPnFDBjIbkCmDOXI
v8h2CeDRk+ywviSoImjSok2U9rSonwc12xk58dAD/in7aJ3wMdIChQ5/eF6fE3izbOvSaClUhKfW
p7PB+y6LfoEcbz/BIAyc5eAkv0X5IEJe9jW4bvCEC4qY2EjMKVEyraw+v6GEy2sPNxPKfVRW5O6g
78E79XAgxR8Cmgyr9Bop4cjw+XoiHbe5Lsp2yyQRHGmEAlzjUonIL8VC7t2mcwf40M2TCsRrF8s6
zdArgDtGfPb4lSKbkVOVapF8Iv+QKdNwp1SRX6llpF3ebTRYSVEAYXChI10yp695MCucKPj3ZoFw
qDePhJrp65Dlzc5hd3j3q6f9kXLV5ZzPqWoSwgEBs445lPperEzOBENXtgMi0c/276PiWfIGp9jp
bSq82ad/2sQLVJ6Lv/GBJnVOjxZJ3zksdLlg5vzJ7eTRaisiwzG+mLaIYRYPpyVKOlNjGha+Bpnx
8hcmMvTIefPpHj1PrkyZiShP0BEu3wY/FW0Vi6ZiIwLMjzYxkZYbRMp2CGYUvK1A1zh04VpxwHyG
aOqsGKIf8DBHnRmVQk5W+4eICRA31UEzqDllvPVPYGo1SDp53Kmu7y+8H9by9yKavLQA/V5jt2+B
cW6qAmmK/wlq5H9OKCPgRKv9F3NUmEAu62cxgCb1FdvzNWo0+I4AJecUSy5NLlL93vik3s62haPy
8eF5AjYEAsEw34IS+API36nZhi1k5z9SegDuvhIHA5+jiI0eOgDOnoE7n9/QdjgdgIP5prM6tdhS
no1aeacTUDAYno3KV/HhBW/AIBiROq/jcneYDcOxgXDy9nKfgv2J+9G9MffIzhq3jF/6MWwtiwHG
OgNqID9nfxdr8zPBsFeit27jV9voGiUz3uWSUf1/1SG14ku66obQiMl2RZcnYIoJr41feunN/SZH
msT3Ge+sWpua19yWSwLc8QjaP6Oo7xKOtNBGgMOv+T6Rv0bgalwhNisy1ZtK/x54tgBsWRkO0sje
LK/EanQ5WYpD63yzrUjzOuZpwN05P3MFx9PzKt9xLHDwK/+iMfevgtUpWIKuPD9mQtHk1jAb/Smx
Q1B/dyexhitjHF5zylCe91tEnDtXEIinyTfDO/1nvTVnRUXWHWgp1i+aazQeg+h4f/nGBYVdAvJI
4tSeqy4MUGiSDQozVAIhAJZeKYM0tHEjF5nWgibmE5Tz3PFqPmFlyYwDSJhemAlZJ33MpSQDqYQP
MbCWe0cTX4phIgPaJQjU2SWassxp1eyqhWmzpoFUJhLYfEHodzeUCP3Kviva/dR4Wmm4fr+3Q30x
/gi5DHmzIju5JZ2U6EfEIRQQAW3U/hdLqL/6nCzj4Eq3+AsIECggQRZXI9RHhbn180yBGjCLEZuv
xkGe4DlLPh2j0pCj0RNOVrTRXupXx98uRDbFpnOss+hf51C+39qb0xwg7cpBnW6fN+p4q5E3lSla
5ANL8bciINrdwOw/lVuuDPcHQkz/4aaQ4pMdktd3dw3uiqbAnbk4mtb5YJV4mEVYFZQmlJVPZmji
gdiMnzT+m5xYR6cH73KC0IndwXdFZabcSW/YxHedMDkP/L6o8F6gmbVBH1beRE+tbuplnLaPDpcn
OI9FyN8gyO05yfLxhkF3ZlLtqSKbOQ5Qz0Gu5MzjUunXqpT+uEyJNoLZ9v2Yr9VqmDTZ49Rmho+6
KDENt9B3IKR02E+UJWCUMFnHPsQEMPsU8WTStn+k+8hZ/rUeJJDBRGhvrntsyXOYntdnDAyhH7t6
9GzFGOpQUCiuUWHAK600JvrpRGgSC+dMTs3Oaqnl3ehpdktnxGzpGgEtx0/RQh3x85P7HXt6BmMN
sA/bTFh/BRlxNW1CWrj+SYNBMSXgIMYLaSddboorx3Yq8CqL5jFlwsebd2QGqR4pZN0kejiBk84T
54V5VI+XyYLD2YTn0gh30De9Yf0ePCKmQRXz1AW9AnEk+pM2gA9uJYJXSUuZD/GWw5yF5VK9q3cH
meN1Dkf47ItOZJ7ldo837SK9usN2/siaZ+YiieAv24WNT4L7hLUspNcephhju/cEWQZl6457PvXY
WMK0C71uIGEn7RPoWoyffjsmDuNiC59CjvdHpfx1Z7//4VXKDG33MK0HssK+efKs61ciBFU/ryRU
XZMsz4cgxDsXql8NKu+2zUAxn69c5Hgrp1nDv1u1dGtZjc16Ym1aqq3Az+9nrVmQQpLy6qP9MoMK
AeW08x21hA1nexUXBba0AjV3h3J5Fz4lpcXxGpAk3CMmL2Hj9xmStzzhy/H679aYCNaJqzdAGseT
MOG7eXC0eAVep6VGgGEclLWwPjM/++xcCHtDUmNPx3uk43z0hUnbPz4r/gKxQMPK1YPqsJSZM2si
7K1slBnFWhxbTVTA8QnlJCNZGYJzGVquB6eY9nxD7V2xBjqPX/sXT5D9dw6WD3s/IG1KFm3SJZPW
bNnGK4vDRFq0A4C3sZ2RcGgevEV2G5NB/Kg3nT9VxHdoIx6O/z96LaGD/Wb6uyfYpO6H14XxHsDD
vV38c3dvm9gP7CihO6isw4CFPU/6JTPJnD1d4p1d4VWYn/sJBOfW6iAlu3Zi2c1/XV4POY6hMDBq
5Hv4p7MWSAj2jJwEnyn3qGsKqYD5Rkx7D/jZEVo04aSZg/9lSqkvJhpinf4h63sZ+6edBC8TepTV
3kpKIExXZihedmB89n9RrHVRpMYtJCGpsD1/+v6yYaYE4jCdKI8Mnyvio0TA24dbrMDGL7kmWeYN
1qeJLDnmzQGSdD2gErqJR2IXVZe86aiO8j29lyxoJqdShHPk0oUAjUgZvB+i11Zz86BaniRXIS5u
/+EK3Q46wRz4DrD+7qysPqrO2n6QnbPFQV42YcJVy3Irz/tYhxfcTAgAGKbNRyhbrT1vFCAgimD5
++3A06cmmCd3jeqHfLT1CU7lMsZLb+Otjes4XEFQY0XAAM7g6+MUrAoDDaa05LKk2crZaPgTSPz8
ikAe53BGzqVAWJPhLvHY6HT/4f01c1LlxqXHczIgDA3DfzCexChqVqRKqzgcMcLFyxQIHQ4ub0jl
FlJQ1zromxdSvk1blcheKI5cC3nTtWLU2jc0iX2hjW+mbOm2pFdVwzsid5cTRvMsoEKyjjMdZKFB
QJwdAzFENM1AVyjfpr/nXqptu+MAHVJdRtvyERfKbDpoPYZGgrjx6YAM1LNtjfCffeR9aa65O6zV
rspu6vYqcwIeX0AVHUyAXebOvDWhb+9iS5rJ+FiQUWkWRFMe0k6QEf5gjWJi4+g5TTh8ms8pn6HP
oUbxUS0cdHB6AVN2SITTpVDni/D8DRi+wW3foLmCQEd34z6wYXY/KiOeE7eotBUY1NErEAIiBp86
vDh5yrpEcVoxth1EdCumSyO2oh9eG7EyysmIfbQLPxgSOtUaAF/FH9a0X+Qub8XQ2ftaGXsMktk5
f7F2z+fY/44VmSBn3d0WKHgZoPe+ycjdnPbcee3fUkbnQkEuchzxetJk3GPdv34pUecqA0kBULj/
VZ7A+lH29l9w4qXE9U8Z2GUJIGWM8ud4KIjQgfla+XGYdMtBKOXiL9/WdqqotQ2ap9T/6ET0Iwe0
h3CQUg0Wv6jMWx8LAQc0HkoqTmxeDB7t3zBs7+/b3D4OzLeGKbrj6qh5+CjoSKGM1r8EurSqMomH
h6T8kMZD9Sr8sMc/ItHsKxR9Ptcs1/PrQMHV8p6yau56Sn+2job/jV0W1Rx8GxPo7WWHzMKZHXBq
Va6cKyh2JmP4QdUDwkVLmEa6FWrKMGyi/5RSR+Og7JEtIxHT3BmK5XupMH/ZL63/hJMb98zAfW4q
xvQEMK+cbA6aIRGgBuCVp49H4tUcvdvyvtglDnWqt1FWnTbvCzY3zUN3+29EApHt2nr4d3zDq1yz
IlwveaXALpH2wW5ZP3BDuy4muf7/vgIVcSvpCghiz+OU9d7Mn0SRjgwakZ5K51JKzWyxafZy5yHI
eGumiGZ7DpcWb4CWS18fJfPczBbmSUVZok+ZsHF+gCbpv3X95LQWtKPDfSweJjFja6cSSAeImHMF
FZr+ON1GldgM1QeMryaGcPt0JgG/mQsxDmCXp/yHxv2r2CXOTCJLNb7Z3mr1JFSlUqo8vYyQ3ylY
1T+kVqKJshmgtFo/OtcqG2qh3ZcIS4asAQNoy7AeaD1I4pLCtF5UqraldWgHyztEUvX4nVZe9kgo
0ZhZw4BKRxgK3QWPxz2B+bfuIKqzdbwy93dS5Z9+vtBSGOu5fo/0QlUJlMPBYG1ZBgXmPYzdu1og
uKQ6Smnt8y2IEhQwmTGZMXTkZI2rJPlz/28GgG/1M74Yr7u7eefWIycky7XCcwxA3KZB6kujUY5t
hQLxzVqBktOVXpLZlvHQRceHMWiS75/YwxFlowFc5wGi9OhssW148imUrVkoedAhnQba32oBiYSe
I2Te6YPLdu1v+FGOUVOauzmwjAMB0QjUM+m64flj8BV7ml04S0yxIDFe0gWgsJ99nr8wBF3e5yBh
I1rhGdHTi33JP9vPo1YoWA5bI9VuEUHm46WISmdgy6Tk4ICGiem/i4oxj/BN4Sq5QUTTW3MPt6PZ
8D302M5lB5G86MmBeNJJw438DnQCxHx5/VBYAP/dofjB60n42UkIq86GMM1j5dODXoNyzYvChULN
Y/Q6ddbIdqmEG79aWsBvjeisO8qrJhZgOAjjShM352ENh3Gd0MhwLZNy9q6FJofHgSuPgzeTuFAg
KpcD4zhKNDfiUrtX/I+C/Nn00SZ4VOm8Bp+AnQx50EwCCf92Ob3SFhRfSqgPTpGK0yjw4PsFs0X7
fCqtOu0J+O44A9DTAipqFbiNXMylDEqdyR4VcDPBiZf1tAmICU/hxoO7iIE40SN3fDXQr79PTta+
3rl/VXxZNL15uckcp8Mz1ChmYAc2AVdpXK2l9Ts0yStdXxbRV7KipmmV7JvgzCw5SMynXvcHlNol
ENDtdBTRyrc7TggjSNqKn+sh1NkrocKT8HEoPpTuFNAmr/OuvObZK/h5WKmGM5iezUTXaRXtmWum
6IB5xERHPMkgKOxL2WuHB2RIVbOuKSAjJeYumx3st4Z5ildN11WpZaEjKxRgST0sWQ0n3memBiQ4
ebE5WnxqJFYTWOhPpheJvMYogOvIh39vEAT+4anJrlwiFrhHvpbE1YJL1PIbsCaKxigykhHYE9ei
I+rnVd+D4z5EuHVyT667pNW7GLt+RgRridEWiy4zBWwPqB/P2/1UrlJPdBeXVphV4cnbWbU1eHIG
VVgXTp7L6g6nHCWyjTIPHClSqg8mgZx12+QrEmYFyNOn4t96dWozVhXBQKkuPkpxDc/FWfM9/P/U
aCay6gIBI6YxF09o4Bj9hMgvkUWPI+xzMF1338wY7RcPFoI1nFdoRTw6Fmqf/d+tOcKb0JohIqGB
P7swlFcwunDdX81EXUoBZvT3s7M61wpoqe2549x+x30fbRmSpJ9YeVPEhGWGMJycgiW18ePqi/MA
L9mD9e7n8V0yXtrrFEowQf1f8lSMm8U4bMEjMgwAfpgOoQKyRfq+fl+VhZkvp4bEqrNIQ4lyHO/W
4t/2Him1ZLsrSiivdcjv7r+4eSOZXpTCIcC9IllWl/Z+h5JXzMKGwCXroCSK8s5ShRMcKItjFuSv
KIKr2zVuXRluEh84Xx1pvMXmtV3OzFTfDnUBcUvv7uCJ4hpzncXkYX1pypFaWcHCT3IwK8oOR5MZ
X2C/cpa6IhsvWm+YT0/Wea3BC/3R4Fu3SGQNfRV24jK365SuA7Ga3jFO3c0rziYjfSl+0auqMdo9
Io/AQFWH9HVdr5tTCWMceU2GbHc3W78VI8U5C88A0Nu3JAjp+gODhsKxnSBU/D233Tz6QuZ4kJ+G
K9wuJGqITvaRrxWy40K0rqhzuoIoa6Km7uvQATTeIc+LKfQd0y10EPYQWFtVqAhaXScW/4wN+rpC
kqXYuSbou/0tcQv3mhTdIXEziO9yNG/SgNDaYS4I3rjPe2DLdb0db+ajMNo8ZndYnc+HGQtKtf5T
Bk9NBVwNFAQhhl3o5n0owP+U0Nx9LgL406FXnde3N5X6tSp3ALOBF/WCv+OO/jCLLNTHlR6si05k
ZCc5viopOZoLSwbwspst8+r+Uzee404mCMokYPewL1bkGB4AFShEs2kO867z8s0iyX+usw2/tzZP
gJ8KpJWx6PkVvK3EBe0D8kScVl/+FtmLBLJqELRl74j2XH9YscUIekb8T6aHxSCm3rvWMFsJSt+G
bSayy72WMRYnByRl8r1Kp1Q1/4fwrh6xai28wl6YtgnirjYkIm50abUWkRGy7g4VwsLyvfhq03+Q
omrYrQwMP5JY8++gsSlWINEJRBVgo73deID/4g3mjrZgx+Zv1/U5JpccBw6JXKhEapRp+f4++pEV
56TZUu/74FScZOaUNXYx9eDS3lEADPJZCF3qSf5qroZakiUxSFH0rhAXbQtpDJybeV6T08ZyPy9h
/oaf8+etVA6X6j6OXiF4huX4kdbBTDQ3ZrHqLphjCGja0AXdpnINSVVMu80zI0FyTiPDqbogMMRS
FHpNsLHJfj7hUNgEd46Fd130N9/KXJ6MTs50fURGO2YXkS/aG8heBded35elwDycUIwfM0DIlatx
Jk3yBySdVk6asbKUhMtzCWPuUui808B1x3efuABRjOGefGN/OkLMld2Fqen14q2D64v9cK786AOb
+AyFujyeROish1s2oBO3OD3OTl2kn7CvkO/hiNMVMcVHyAqhepn2xrB6S6dMmDpHVMv6zbWxRIdE
Q8BXpqaQ+LGCSiIPLMV+v51JWqHdYXHJilh8g382wDP3kdR92c1ODThhcASMjL+lr9ldaR+d6sd4
zaVAuDeXfbVCqpqyTHp0ApIDoYDnzELvimAW44sWCI/vPfNnhjL4gddmb0Wl6qthBaa8zQFd/b/z
leeAz95PJrW9AvtWBBFtcqHUUnv9uGYtCLHvIMpAcBssIxsmbFOsdMDSdTgFcZVVQvvbkuYB7l0Q
gxeBLGIdsvBvbS09NCP8PcDPx2qjBq0mv7BVr+ov26oQ+EW5p3goqBAicxTpaM46lu8O2ucUt7Zo
93K4NvKi4eU+g6QB75sKvF9GSfFYvQtDjrcYwtIvQWlhRAYEcKdsUhaUM1oC4PzuWGgdTuMgxwZF
KztPh8DjFi6STi8kKOi3CDVYEPunmhO6dFImToSMFQaG1PVmvhs6wkg8HqWPWjNGUd49fi1Ofcsx
qk3bHCKfQqtiVbN7owNba9jBWU0bGB6fcn8gagzGP4jQTExXOWiF/mpLS8BoukYrh87tl5LtcY/R
AlK3Xhra9SEMxfvtDn+VuGh29+3w/7x8fTnIV2Dj+dc3FEAg9unfXd3UhLCRJeb9hTzlx15J19hl
aoQEs07+O46TwFH3ItdPcDVcGcUDgsz/GWvbozArmEuzL84WuZFle3HSzYGxaIbWlIUaIuz/SCAP
EQCKzzT5cMYZVYiUOPXg1LydQKK9S6yhwp5DiKL2TlmuJGzJLajRicz7NpJ1OhQ/W55JzgcGTPbA
IvI0WGuiJVBIq8WNtvFkYblzeeh6wx5nKAPk8fnWO3FiOaYWB5DmU0e+86R6+qNGlzKDzta0fo67
UxkyyL0J4/WdPtFolocJesNYMOSiWqVcnSTWMq7iVy54AvV/CuMvhkMYKzxskyDTcGb7FCLXUl8p
0vbUfsCq7Xr5J3E6yG9Vsv6BmIPVKG3NQiLRr4IqHKF2PMe9K78vSyaYZP8LXlZa5NQZGg723Qve
hNxkrl0Y1Q8f7dmEQLYnQ/4vzAzziI1WpLve/uVeU3yLBTE6boShGF2x9xAZ+f/i/L4+fOFf0gSp
a3FRONa9rvDwMifkV6JVCizzpo29G3mx2AodwXSwBB06HT7rg89cIU2y06gr61U2hYBrxLcZsFtX
eBs4BTZsa4TDYrue+LtD0HYFu+AKSUXtH2UKNQILl98yXcTFtyw91xl1cEtfutLYQfXrio4nC3Bu
JJRJoJIWF4BlRBpJVAG8csshRQ0/DV4ssPQRFOODAd2rP5ChyaW+GXIFy08vq/zHGtFUhRW2FNR9
GKUznNBJbPYIF1ZvSli/nJJ9AD/32s6+FtSwkqDGwLwUE+RtSRTQbqiQ8L1K1FByfPuMfHI6qWSc
8Wxa/07SxNQgGeaJcbZPmQ2AbKC47nP+HGanNYTVMK431uEQawyj3eRL5rUhUJg3ghJb5mxsn7+o
aMn5ypra6pVNC5tFb9Iq0DRiObP+3ba7Fu4wIhHbJ/OVd5VI/27srYSvs2iSASusYlfWQ5Y3ZeSo
sw9foqfmnlWTK39D3s0fX6r0mR1bwTuVYfnzqoytazptZCPaeHn+IkYMr0ebvGCZ7v789Rqr/dbD
aLVkyiQsx3wutulA7+BBXSmttaM6l82mnN1bUg0rLPP+7+moJGnj10r9+D7uJGndbsXBa8tYr4Mj
N8KVo8F4ZReR03f4fUrQLMDgDthrWMExb8pHqIEAsQYEBwBU3wXXkSllYgpiP52qCg/MP5yd2a1a
wSGjT7eZEQ1XrFQz1e/FoJf0AZjgLi0BfD8+XlH2eFfcEs2cZJ133lFwswSe6Redqqz7tEzesazC
Cv50Uy5q7LTUmGTTxJZb0Ir2/tVJUi4pLg9/RiIcGAI4aMVPf8SuEj8utvAM8vPjwalx3geODdhr
+k3fVYCjLevLfxu+B94PPH9Dz4deF15r2Dgvjx4hFghpDd6TiDrOg4CjdVJuaKngcRxst36HOqeU
FNWqPqdwqqAIkAeWpJXbRnMHZtEBMpnfmqmKJwNH+BBCFMQCz5ddez4W+xSgaPXxYowLbI48M9df
P3fDTCZO3nbsybstKhZaEnL6/Z0ZgKQ3ikD2U5qkknFfLnOubBrNx1vaiqCAbr+4FgS0RSzqAc0r
wHnByURjQaGJGVsTMgl5T4aijqbN2sCLEB3fYcyKjP5UfdqHLktkwNz0PC5DYimSwMlxr1fxSYYh
uU49bJ3SWwHcpDDpvfefM3Fy3ntAf8GcugPxyVNTt2Ztx3EFDud0xg+Cp87E3yxvnw00WF5PuBSQ
QlduMITarxw8xGowaz65xGIRWtDMycfdoJa8VbxxmXjCPNtOODmbvJZq8CkBaYLdZZoXQLDFiQ46
A/cmkAqAGV+Xynw7pfwloYKdVUWeRjghgbvZOCpvdi5BHPXDeQYq31UXNqB0vX4oYFzRK6OQHtMS
cxIVVTDs5mhhKsP8DaJtW4bTNJG4k5o4gzAhcFPfjZdXKSBRNJ+7ixduz3kh0hYrmKG995gZjTXM
3ETivMyOEK7DOOhfF6Anm2eHfoQMnb6GXbZq5kW6QjjnydLKgMHwiUuFDDimb7V8dx2mQpHPNgW+
mja3OV8yEX0PNr8iCy5ecC8zRxK/dn6VmLozu96wSk8omKJXS3QVPKn9le7slXHqTjHfstkr3PVc
cR4NnNQC3G0cBzVkt4Ky9wWmnxR1iGYZ6Vqu2SIAcLkBZNyafpiz0NTTq81NtcTHNWOJ27uxPC3b
be1CtlRuGYaiV8XvVPCkQZDelfD7aTlLOQwUwoVw0klM+uShFYMS52aawC43cA+si9Em0tG/92mU
IFkx0TjvlYFHGa7XJf4SUFUTdZseTw93DeEcKI0o0Xnq9ILv5cCKRcZdK0TlHkm1Oxq/YSaVNlIK
EzJSHcSETsfzmi9BdtGgJUHE+bot4co1TRMhiGyc+ua0CJu5MTPon3zidfGUSKTefARqCCQL1nr4
DykNF9cnTU74X6hLNGK+sFtwUgPgg4Yu4yFnbL3etGUsZXBRsYr7a6S7BN49emGEzO4ml30yIsxY
UwaM+vuC1H6xN/AIMTmANhCpdEmMnjh3dLIMXAJtxMjPPSxMPE+CDSoboSY7nKKTAG+9kTejCX2H
vSzEIzgaHGCQrPa2dTrM21Yts7kOoxOx3/uTceFdl58WdUnUx1ph4ZPGeLIDMZCGNA8va9mOr8Pn
26N4yHiz8buslJ0S3MKUdBdvsbItraIV3ra85oF/cpbtjmhWlANjpAwB8TdKZdzQ3OMgWxWGbx3L
EecJ2S+Ehpf1fdAHfzkdj/IATJmQAh8Vfk9G7XwD1tjd7NQ6CM95f5RcS/kBUBzPWtpZmwVA1cyJ
Z6a3TeMbVccqKVtZ0xyYcG317yuc/GI964zt5Cnzz2QJXlvkvQH+uGAV0/z90qGtFH2F5yVwAhtG
3P1SdZ/I1zUnq0787M7ulHAjB0MJchI6iqxbmm6D8qOd7owJOlas80E81mjgjFJremp+KAYImdm1
NI61D5kdEzBcBVf2UOOm6RrPjxlItGLx+Kl3L5MBojww20emTrcpFIj79AW67rKDOJnBha4RdfAK
Q0ONV+ANtsUo1NSMGrXk0gpMJ8VYSAtZnD9sYK0kHWexMGD5ZdF712Bk7A/y8zCZ0kL7i/RJvJjT
uDHaboTDfd0L3xWFT59nj93k+6MSjwDB7wEKmVWrzpm9iVIlBiGHqdcneNeiq2w2LXE/xjzhpEOa
kzDesYH0C92yzrlLWSpv/p2vYlcuYlKSpyv7umnaoflSBxANPCr8KZ35aknt6cTOSFcXYESFpjZG
0rVZdwDTmFC3+zHcu1fbT62xb4+e/gifBClVUQOIFwaU+8hqJG5ixMzyF6C13sQSB7r5G+o12p9V
9c7hdCIO11InlZhsspRB6WUNV6fwJNmnVn6Hg9+QTPRqpV/nUXadyrb7oskMx7XgGibga4MIfr1v
tFs4fSnjn37wJHs7aMweZa9PVMpteg8FdEdwU8wBNOJ+y4y9OtnQgdgAj7ZSEc2td9WbZryzIHUo
+uBggAne9CYmpBL1QmJh7GKrhLxphERcwkQhU3hLYfN8gV4Y5nLx8qQHXFCJPHCqLpSIABc1uJUJ
Yc2+wqHDgjY6vgdqRlJcpDyTT3IVJ5ISGVoUm8Dk1gp/n1wY7+D2GWe2hGsXvLoMNhK+qunF2Rjt
/W9gnky14TbtkFwRwbie8XEnRYGwIdjGyGQ0ZsoQeivyaWNFSlJjBxuvv2tucS9mPbXEcx//PZK4
F8wgRSy2lCwBSFxGdZpNfZYozSoVzvhZzHRh51RQIcCEjvvvD9U04eB7UUMcOHcnOsE6ShWvPEu3
1dsXQ3cKm08/GpdJm8glEBGb83YGTLb2de8AoJUHb4tHGX1SewLhXeQ3sWwPWD9xOzaw8btB70ze
Bju2KOZbNmgVNN8gpKXzF6cdm/UvPQ2/AvPgxi4JY2MMwWB9jyzIGC4DThrjm9CZOnZYFoDaoD2H
eCewRNIwGqKWaTmjt0izLimb41OFWFPS34da4jAUT1IdYVaIXoYCbzGXlYYmO3t6uZYZTJfJuh5I
8FQFZO95AeB1h8a3Cq5FReYhtPeYBEbYND0ayZccDZMtQSYXgHQ4SH24YmdGf5iInfweCZ8swf0o
IEl4gWwsLRZGPVMWVac1yvyi614inyTiJVFR6iZiMyRWsF18TyhoTHOso/xhYZrsk8WZD0H+qd5w
Ffx5zZgvV+OOloAlZ+n9kKv/zkc1E/OqYh5W+mRn4WQPbHLfTGEwsono4qr6ECVWUyDbJgK0It12
9qFqORsgFFEPDcTE0pLiKUDqsb3c5MuXPxpavPN25AprIpMST+I+EO6P74VARizdBGauC4rRpc20
Wz4X1mrkGbIzT0bvDJMOGpMUOUOC5IXmzxPFp7bCrr2PqLWRvgFGRODTHdpTjOIguzQhAujFF579
2Su6wipqBQE6eHNS3/C/E3RwcdLZk3K0Hw6HoB8ReTGGfoSLrbWFQURjRL2CAxX+NJSGjWs+3YL0
kS///Brt0furUmsrMFcbEvD8JFm+huqOqwVj7YkzO44r5WnSfsCirHAsAqMgMLx1QlbNFYOHj8pQ
xCAB7QLDeXYil62y6Oss7LkXww4eDTSByY0lDRq836IDpMjS8yHMeRVHt7b2pcnUJmqac/5OAGoa
vZ2rSL3sKDDMut9BM1Gkz/px5x3DhRu0yTAX9DJKXl0YYssLRJDwoGEKPMb62Ez5QRgeEFdiwx1m
yFTDsTtYShy3CfxRewewBYGfvmHPLp2960CEjxKyU6NtR1a/6oYPkTpKEy+Uc0YtFqptVq/8nIhs
ybloU4oXVHU1EToVa2YFCFePJ622DOP4kG4MviZz27nuN14Rmk63YX1DqbVsDB6jaLhzUKwVaws1
x5GvRno8LDe6sS1dpxgVfVNMoKXdHWnJsZKvnCBaSd4rf8YNCZoxSBAdU1mzoG1uGfY0EERSdyKt
hv0vD/iA715HRR7LagergS6bAxAml63jUUJfFNwrpsxd9hX6ZPxLxC4gscZK6eYzb2Co4/GvJOXD
+fjfX16ezsrY99BLyUOicX3O8/G77k2VLmkvB9QYiy46XQDguUPALZvVklMXcyiEak1A6igXiReJ
EUXxwQfK/2WEquxhimREtkgVykUnDxaLWBuS94D2RGqL+vVgdzBdcXtDuom/vOX7b4XjChjT648o
Nsii0N5rwp8TgQM8Pc0vlQhIWdhbQCuT3QBs3mugvrKSWYHL31v+BNxqxy/Zce/0AwSh5bB5PGCZ
O8ozkOsVWYTUcDx+1lpTnJuQqZxtLzOOTNqczbrIZPCvQwpnJHqUK7N4nmq4epIxmpaTfNmhYf10
4hyX676y0A8HQpKBY8Al0ZkJUR8jpOpWz+/4ESRfQN5BOfsOvMiKygqF+7H7PZMCw+sQywhy4lqJ
kBmPlwpFIzO4tSphaLxTF41E67XLSlQnCpZucFmEB21ulaCtLVCuyDNf2U2DJOnMbGu0rMqNMQvI
FknBoFk2GzQUJf5Mxm8e8QeaMiOtSu5iqBfqk6TmopMKGXgsbUefBUouerzeYRKkSHN5rCfOCmyw
qJ94C+zd7sH9y/wbKMAgYtd+0PMwC8nIRH1G42lNWrjw26PjDmXCEgvefuBULb8jEQnsdllTyhir
+fPepRmZsz7TDsyBoIXfKtdBkRszxGI0EAXSRB3ri78wvdg+emyn15zSXC1SmOqRxelcRDNhuEDh
LRyw10OEOT6G8QENHjOzb1I64tAmDn4+UcjYOfOFlyf0XF5m5hv1AdsxwB3jm4lLM6sXyjugr1q6
pRX3JtwClC3sDUW8mEorY/P23iQEt3UG4wUz4Clldo8wZ8T4J5vcRc1XE+hCvJtyKYTcrdu89uPv
o2u1rU+5q8kTSBb3RbDGn2lfOhuEnCc/TDnYPJdnlLfQ+59OjSVTz1upIqLpY8b8v9qc9g3rphPG
wELxAFoAMGJPmQLZO9X3dBTfamwr0R2pS9+kueLthKiyzocEpxlVGDSjDjMJnMQocCIMZwTfNhZl
6DvvM9cr2Qp9npuaIVgIBUJkHFjqVp1NgTYfKLwFiC9oQJ/pagkbcRMkl0f9CIeYSp4GQgbOApE9
ehrBgTTPMNSf2pdG9BmMYv05iDZy6B4rqT2FEFwjOoHvIC4UKciCv+tZJYhmjXEhsYYIE+VHQr4e
IKitlNAyuFAtu2r6hjYG3iFb/X+Qm0UbiSEAqKtMYJ3bKwjJ7DPrXrSwhXhk02o4Z4Qc82uX/bZx
SNq0KaFR8jUb1tt7M3pqykLTodyw8DhzZblFhY7CLjk1RG8uVMZ/3pqGqm7Av4rDA08SjPbGPyE4
ySXvoF0AIOVSekoH5TUbt8WSMB7Sx77YvVYu9skzMAnRyVo+fS7TjF+bgJCf8S0Ob8o6IQaZoaul
IEROrWCZsMJiJu/uYr5ZSRXsNsvq7DcJaxShkc7Cy7ePf3DgPuFU3f+Cw8rm/9bUiuUgHNNNXeqo
n5PKhqFULCuxtgIDgsKQf0nnN5LeGHERbNF1TYGwGN03vIWFgNKCqlNfAHeNs/hnVtV97yGwlfC/
5DyZONRf5lj0ZMnSoHZ9vf4UtZZ7cfh5zFQexhKtNEaMDoFsv8gfd9h5gZaNuiTE5TbTh7NqPLtX
gbGXvjbk9v2L5UVO+A6D3APu0w9+6ZakgpH0UoSnqSwqHj+hkcIiczmbyrqHTdqJEqLm1QOkcfjh
yOC3eLoSkU8452e2aEjn8vKrg7JfpVa/Tq7Rh0edA3YdsQH+0YqTWn3Lx05S6jUMiZmw/CfG3ERi
ZHNeAEBLowZaBpOEO0u/8OBx7C6b+Y+URkg4gWyx+ciu3YVZnW8ZKBylyZSYRNSPo+UoRO4QBjCq
GQhyKUGTBkO8hMJI1AvoKJ8K/jW+RMV5L75g+H7/UXqXzEBL0OMKRo5Szq6Sape7Vtd59k2s1fC3
vAXLqoIDr/3fer4hzPkpzEz2hpcbdzhvH4/J1JHlmqUTrdYQ/mJOqiZytC8pCcFXcIPgi2x54s2c
qHvMXUlopdNPTFoWarsOu3sv7fWtwa7WEFHoJ5eNS6f9hzCNV/iaUNJDsRogyDp7wH4i70tXw88s
mXWb/b7JBZvaehyg87GdwXU4VXBxt1SfNPrMUbiuY4jQsudUMmbzOkI0qbOj5orwiStVyHgNVQ8F
m2+9yiwoI14KRmHYpfFNPJygK8Yx4McBZndVtUGMe+wXd+8A20w/TuhNEuep/akaGDF5eCZRBC/X
U0KkEvr806cXXukKncrctKmqEyfA6igENb91URsuD5SnXjdEI5DCgYA5uLCUsZAQqY7rpsbV4EDx
0LnnA/+0O6AHaKoLN34pBkhrF9q01ffuVYwMLiOEFosvHCHrSzpbDzlEk5ii/0zOvSbKrBV/gTlr
auZOb9oUINOiK7p4cHkFXZKWGOZVAVM8nD+WOZhHZ5CPHChRClKgelcLsCC5YbZrgk0AL5AkRnBf
WdHzJnvr00QljEFJmecF7BCTajn7WUr3iozKsymZ7TLAmtofiDNM5amKIZOhI9sTrTfJLlIYqxuV
DdLj4qEapMvv7MRIQdSGLYUJjtQcKsV0tKm8AWymyiA5gFgRVIdOf7P6PFTy9h8hQb6+/0pQ1pGw
FDOUepRbooLOFMFmpxa2o8Y6VUTXSPF5OGbWKHiIk1SQ+gdIHAk6ktVK16LFZQFpwQ1z86Hpgcd4
fMAgpLW1DEXyQj5MeKxk0vb9J+HH6+56Wn49aDvZY1O+4Y1dXIh+Lmeb9UPMthAEU/GofNWgw3J3
jOwIr9fedysQ4MrNYxmOwMgq+tpvdK5eDFkG5eo2v9XQlIVZc906glcIQ5Ws7dkazP31lu9TKfMr
bIL10dXI/hK9O6cZTcfYhFpHRr/1C7Q6yIP9D8YVNsFKhwTkut6sSbTarmhbrGghVUTqHtV6jj54
nyPSL/RUOlN+ZUAkUIsV0zPnPB0eEaaU/8yHn+rYZMkdqok57+FDD63EoHOgs5Orwkgfk9l6oAzk
fn+VbTwV5QpU0pJvDvNMHqNKRETjNubJEPMpnxY3AivCmHCs1k3TdThj5309EA41uQMgUhPZaOdv
PQNVf6YNLpELYHF/RS8Z1aDkIae22rs2trWEVjhJaI+zF23MlN5f/MrMfBZFvMyCN3pcJPg9frr4
KRn8s/OqVPNATRKYFuB7pX1Ws10EUMYzyX4YmJM30BguZ8iQZfHgZVX79h6+eTXnHpvrzUA1ZfKb
z12euLEEx3AOXRUjkhoyJM+FO9F7ay/bocJw5wYBSyMBYol4eMkEHEw2INrgmcnQ7ab1SwzA2DQ3
BIqRRnTiMBp/qmz4YKBAp5dfQ/Unvkag1Gu9lo9tX+V1RGY9Qv7Au3apw6gn2Whkk4JpsaqkTj04
coyGMeMV6VulBKCxsqLW6TV5izvZ57LdI2Fw4L1aAMEDMYbvE0bdZW3p/AtqyGV3XFJM2mzguhB+
AV57n8Wg3QzQdsmdb7241Jrcz12kUL2kGh+aRvdAlRHrpLuFaIShohw6n/SiOSEFPLEOLbDfcwiW
17zcJSOtrWYvR3e2Nnl4+XwkdzodsmuDQ2Gygo6NqK2MNOq1vRoGi1j1KNVtEGSMqqksXOAuqLb1
F9smfLeciza1b7722sZqwPoJEWGSfcqd6fFw5dWiW4mzUpSUqbaxJIlOcjgwQO4rddlD/1z7CpM0
l8ALPNLN6UkG9NZD6ipLDxFlU5sDzSThPHsvRZltXRQF1FP7dxhoyDzWXGAstUroRDz5gn2Z7QK0
Rb+XMIaNjhXxFp+DN3fWKxZGzVeDnuiF9qvtP1xO4uPmWUHApxGInz3kG2L31FnFZc9saG6eyK29
wZhHwtJpS9gyYMFGdq5U/OTuMiaPSsxuAgaLoBJ0JbpDhkfTtxtgyo26xI5XY7cQYOgMl6WZxPr6
FWJg0irQBr94rrN2mmqnN1cak5MIxETh6IDhNxG4CmYwN0medDIyhYgrKR2nnS3eJHHDwxcm70ni
eQawLRe7RmE0SkS7KsY/I4Tw3+SDP1MufUe0jH3zX1hAKCXXcd6F3OwYUHCt5sz4XfBum61A7Jr0
AZpfwbxsscRp05z+eXgWtgJ7l4Fz0b6ZpJzJbKBYvMcbutXSwdoQHCXpbFR2wH4J25zGmX97JYEF
Z5jNvHRqce/Fr8zoILY3KlJggwtLy3yWMatya968P6+xsNhWCx9YASrr/He1xjNHtucmxE+vcOT7
Iaiz0RTCzNzn7AD/Dz8lzdA4lJa8ecyW/yc3BWYbJ9CwDtlHY4KkcGOmOorpn85XGXGmFOEHWTqR
bRf+npxvvm4vUIv15mIfnfVlWD+ANxMs5IB/eUVM1zpRCWJ02/iSV1TeF7ZdKEsxCgFKdfPCLd/D
GLWEeLRVtAOPTtCUIIt/GKPPy17yQcJbOLsAUk1GmcHQLrDoxqqVtiq3pxyJW8y/vbOcaH+iJq9y
SUpbuNWpAKaH7dWQcy9/mzwyRe6B+rwPXKcWE+QR2A6abjpIYMZBv3WaC1bq5SATLaQtsPxaiamG
JvlV/OPRum0c6CYX7qkZr8+vKzrqzGFggWTOW5pJhvh+i6/hpaZta8lXvBE3DokdrZR4IARR5QQk
I0OQKDv3dRrq76DhNQT/X3PzQSeh5Sa3p+1ng4htEG7QOsT1bzcij2T+ax7ykGgEpxAbdqGzYxrw
ka8k4RhWbmrXPxVNdgysioP0OUZ9BnSDOyjR2GC2hx10ENUQR3w1BfcShW6QQnkWV+O+ctk5i+6b
1wZoyYITvyVOoLTArRk01mZ0jWCehC74Fovz5SgS9zw3sB90fvF8HQoRVLFlsmK/oP4LdmTRGcql
BA1enJK+LzGichY8Pa/FNTLHkgSXkKoOss57dLFhYHR7KmAyg3cQ9SUWaMwNGVPXRtxw6bv6IGMX
uRa0llfKdBi/jzpolekaZTNUdIhOM4+QRj7F3fgfAAt3a96QwWBpOcWqZeyO4GyOG2rq8uKrWVKE
tVhxas4/uuiu9vVT2JJ3pg8oxucWPmSQ+ZkTjjL0kR9EqwJek1M6t0HEgvhaCxyhkDT2uIzlLGCH
4r94MXbS1LeYdOaAhWviurcrbDctAByODZe7jmDxpqXVOXPwkVR4KM7sVRkF/lMUYrjNv6ex0lDZ
pZOFiJStfB/PXFbOdmv9gHdtyJ2U8+qS7OaxYBV58jlJDaRKDPKywUkEoTgnBIP57e+DPeweh3Fc
fRyKcAXn6ixh5lrAJEH/HfEQIftOfh6nrr9jkLSQ3pqvDjYw1wlLDH6gcNe2wLD+wvMkYUOjM9Le
fM7dHzpaIva2yYQtsnL7da3PknCxAHIph5E3AW/mXWKS4tWL7aN2cb2fEbTVtEtgR7LYRNuy5fua
DHbYSDchTBcdZlFuI6nyW84HftuY4fQACXwxgYpE95iBmPeqy5n42d+3dF9jErhilRfCGzNQvIpf
IqKQ4+nYJc+R1Aq5XqvXRtBPwKE3VqJeH7Omm70RgMNQok5iudywJ0wmIHTySBfGY5oj+2v6kUey
jlbg+xHuscnBgZrgTl1PlHsFwQ5MTb6S8cg/dF09gMOE+S8ty2/JfPcfl7qndBxqlYLMTukGMP47
vLGTtM5Yf/jPg1LZ5lUZOJD53Kjvi0Zseonq4Gmi253xGY6/pTjLFMWTyC68D3fXG4+ja3F7sB2J
VbsjtT/DslgSNiIujwHYffsWWisNR/3DGK2y/9rLTdkk8t20w9SArce9RjfXYGjKIOd+a0kNTr42
Fb/IIpvhH38mdznkStaGUOhe1mXG98F5swRp/fiwQLRcdSBChVWp3ZojGsYHiv7FgyYztgawswb1
/scxF1hBN+iaHm6unxNwNOdNJRdM8U7+Kz5eP5SeDTt/N0tja9EVWjs6I5orbYQVIQgW1aHHlkAR
rzU51NXv/PUYUwsfHYxnJF4RmYRGfIUqat+8Tqm9WRiwuoHacYDhyUHGdmzdgtYqfS8mtr+2eF2E
ucUf/zuoNCn0uve6yXal1lZosBP1iIq26FK0ntr5/6fdh6ibsaRoBgc0nVbOT7vXRkNZNJKoyhA/
psE84yX3WmNINqH+Rs4e85tvP22BEz11sr2s0xuHHL5avuiOaadLCwKEqm8HQb3jxrZoHY2/P+FG
CC5f0vxTVK6RfVO/uxKukSPkC4N3eSkg6OESzBVLS6rK1YNDXW4RwAP+UQZKmlVIHBk3UfIUm97E
ndYz7goRoNrQLcKLl43P4S3uDMCmfDwTQY/4Jh8MvIJLX1woUxzcDqGT2WPhqCOkpenRBMTtjKVU
c0vtl0gel9hRKehlc/+jzlQGVCxntPP+MPTrJwXCnI4NI0sIafA6SF4nwgXjRtpCBr9qe3iAqhZx
WXU9qMCJ47L9ZqcNL08eVLhdDXr9Fk0W5r5LyhJylLZITD/FkwRpjZQyGoirlhcsOn/SrlagrtZG
9105HFQJeMiXcK7NtQWY7vDblNSlGrG+r5HmoF6G+3c4ZiofDXismi/KnoHzLVGy0HT693Sj9rXR
Y6olXnuF90GO69PT+YOg9z/rv7yUpdQ4Iv27if1xx56Wa1QfRHnQbTPeEXN6EXrWr1Zjubyqlwdp
s9IA5Ycyx1ILuY9sdM9yy8Ah18A9Kt/d03P9uldwNQ/iza1Du97wkzKZM6tTctGf49wY62s6s0fh
8CYN4OCgmt0bAqJTSOR+RToI1TCmExjVIUNl7mw/8wRDeXq+pxmZSdOUhSMfSVpmG5MrUts0NMpl
1RQV49x73i+MJTBteaePf7p+f24DyOaOtOQCaOCsRFI5GZiZj6ZOwP8nF4kxGKjSeQCo2FCzUsVK
PQ0AeeWQORL2Is+RZMpGEk3rmMie0l1la3v979mTuURGTvZI3+5FIkMe/GFrfYuTBFI4PGLL6sRD
XgZN4YXwd12hmPvNqUR1VZ0FVinem2jupa4wIh/cL5NtI/b9cy7bPho/OpxYeulio7j270ooJuGV
HWH11GOlmVIEwDmo7NVYz27dO4w93ozuv3ZmZLiBStCy0ni5gPCDWGf4GnEh/3kuhIEoF8kjRGt4
p9gYT++L0WdwvTZbj39rz4f9PH1uJbzYRzTkUhZfoWBLhWz4M/M5Irhd3dIe6SvZ2BKkEJrInwtT
1oIk1GZKiFZg43l8r5H36mV6bjMUPezLAfspG+WCOtBsFtph9gK++V8JlbuRKmX65z2dPy/Sw7XS
pIB3sac79aBwwWbMbgBMndQ4zuj9AzWTg1v/7mI1yuXmlMkohkkkSyHZq2uDnmpjRVR53/CBvs7H
BfoxRfGIazk0iMlBM5qF9UtwcGQvafjK7LDZZyNrQWjDmN4Qn3uI3oTaX7nonX9VQYlcqtfWpWq8
+i8zGc6e7KPwWT9PCg21dvocW3dMNBcRG0elAA56sa+c+rhwDCjShU8zfNqBJpAnLWTv9b9KsyW4
Yswhol36T/TA+83Az/R6prUouVy4ZR9CX//KPM8bkzwcdreQDaQCENMLTBrIv0eCAW1AkA3JH/E3
LeOYVkrcWMT5b2eYPAHVOnQ7fxD4V8TznapUYQvXXg2X/nwUm55hoiaU4hduLVwVT2U0a9tDxioZ
xlnKvqr942yxZPbHHLA7m/3LZn78aB27W5K5baxnBJqt4l5x8QDTS6hpjZY9VsorajpAQEL7/iqX
jA7rSWjSZZ0X13WQsCK1CMBL/KdgCq8spIJDJ3uyvKGb2FaJvbjiH80mjFYkvwstPtQBJuCP0kU2
hoBedskQatW7JqQbdpzrS0r/91Ro8ewiGtfkzJJW6B/TqZp2u0Yj1mnwUsHlCFPhpaWSXKePGpCW
6MlWPn4TfAimeKReRnQZ8vDd5X6aNR1SrlySIhyzQGfbCB16ns74YVwaLCbL/1uVODwASZVza9Rj
BGPFfanKFjB1z+Pqi/KZsz1IFNFNmHZ406RLevyqvTJ+bR7Khe5J/eGV7VLy+DnE3rCdqyWD1r2j
CU+sFLlxOAvUsb2LqZOJPYWOAzYxDzdKUVTXKb6tYHpmY8FHwg91JqhCMm7NC/Z4FluCBSkeZrF/
ToGUv2gudlqm8HdViEyt1H+9rV8Ts7tw1v6uD0Op54MDyzqRhrQg7rjwLLkR5HUy5PjvY7/+1Dns
6XFeYYtEws6e8BABBzQ7TzYg7yzNIGGsDKzmhv+HEqtmGOImj95Z0rwdYjWd5HwzE/rrbf3PA2IC
j3pWobWve/IaUdhEbo0JnjrBOi0O9BJ9G1QQPR2TvXo/FVzpyN3RgErZR+xeUTMax3PvhSequDA6
H1usBSukUrpGuWf2iDdW0BYk1ybUby+N/oWZokuvBY3Jg5+KqWRgwDHnkKgFnnNXVe5NDcWk0BOT
dVFyK7TAm3eW0oQd5BErX5ReijpLsLrOuzOuNWzSkKmKhjGIQe1Ts0U0JMyDBHXfWMSVpucoQPKR
CCZfQYjtaaiIFOHth/V9PNnBf/QoB+gSfaCMXsk9lZb/DevhQ8wlFuecfIPwOxX1IxW1yK/mjg1H
9uzC67iOblUTMUbrSOazOXZZBPEoW59yN/nZzhaPE9uNZ3fjp7w4797hhoU4I3cfCLr/YB9pFAHa
r961sCRtQY+Vskvv8LXdgGLjiN+ezI5sT+7/LlFP7qNTRvpyQMSmgxfQ1WgImKGon0Xm06lxhhDW
q8syPCxkQjsXlMGxYCbJCBGKvIH7bANn5ZcSJ9TaEd8drgdehxx6oHr0VkqVk3Njgt2YZh0y0u36
VbisUjOLoHTcZKrngWJuopUeMV1IMONI8ZvdcoApesP/x0IZLXIGqs/e1b9rWziMgKZrycFnnIrL
Bz/tgel56OLJUbdmhkWQqd0aCqZvSB9OnVQulEwOQS9FNkCvwjP7CQvSU6f49Xl5NXg/6QBZ/mYa
NLf01IwzqnXwbR1qJJQ9BdGmcUAruJqinUUyoSJax34IWjVM7k9PE6Vpd5kWyyejjoqag/PN6OeA
et/9nmgXx20i3ThG3OH29Kj9l/PKaMeYc6XCDF1dOY1GrD+4VCEWtD9knDJT+g3RhlWRK1KKvda1
yyovwzqPCRgIs4ksc4C1l2NkpOv8p4HH50uvwr7X1HozezXqn2GO42Gork/srt9fCKNAEICyPTlB
SfbBYNXaxnawWp0jaqQXCQ+bpzKRESdGjPJ/IEzsuqvs/kf9uL9XQr+aU+9ZaMxeVonPmVh+WgrU
e+btoj8i2870nRcP6Wpp8hBc3CvRYDTRnKRpKFMwjWS1TrMA/8pQDu4dOEb4OlGkfyeLeiYSWIY8
0yYhXk5f8o8g6B9tNvNghUIfFPjpSqQRifbCzNzm+fD5ZOTLf2rMcKlKxPv13DYF0HwBV3xUdoKY
55MsgsKgexLgI/VtFZc9NDua1NzBAYgMGReZVs/IJ/fC1oH6AHS5IxKcYctbUDuTREtooZ67WxgA
C7I75H5pUahVnppQo76EeHhWO7kFwSWuxpIFvnEnoQpTlaxjwn6WTfIDHuFo7dLx36ZX2Eq0BoMK
LdVoKKIY9WJ8Wy+HmzFVI0yGqdfXYynmBFgmdjsVyJGqhGt6vG8FYC1qZbZNvUPT+DYCnu4luqj1
pRcB5MdadOrc+4dYP+qu6fS7EgIz4O05tHtdUayODFCVym5Zc4k3Ea2I6NooafyJ6FpIgXO85UWO
T/VKwgkfdCR725kmlPsgB4+zso5TMDD9oBv0ofCJ/0K4hKd3eNoqLl1H8N3BzR4crWN8UUlcRaI0
wl/kbiH3njbaXsCEl5s/YP5MTbK1PppTvc2JvwuegCFOoTW4umUVczQNgdYAzfVdceJFunVQH7yJ
wBC7hWfoIQ8rzri+HgSz7Xn7DvOZ7OOLzv50TuKaqyEH/FjNeSp7m7x45w3HdiuB0ut3814qd3v7
W21vp5xQo5cwszVd5iaxgRxPLBQs7pHO45FKIBVCtLg3objGtUhCiep74awvFCadCPGza5z7URgO
6nrDLDxSBNELdYVWNN4WFPRYMnY4NIHRwD6HvQK/pA9psacSBreeBZbnWZZzi7W4OOD/spYPd8hA
K+veOYx3sU8p6NgVI+TqVADXOMO20N2ntQ2rTtVg92wgGmD/5oFE1gMAgcelQSzy9UIGSGfogig0
KTkQ9uiNOZd4nnCfcsmA36wM0eFfup+7A8RVucZYejOCmnA2zK8yVM6WNfWLbN4QTR/ezTWT+2Rd
h4H2OwPPgmjgh4zVQCpV6oUh4K104jVk2VMp0l53spD8SPvFhrFVjvdYjYyIc5qg7tPYnSH1FDis
tiVtf3FI8t5Kg8YiYDZr3ZAtZl/I3BFxj7SC0evyKaec59jZ4Fshh+cO3Twcs9AHLltXOIzvCHTI
pqxdQpGYdgygL8V4mGw0QWY/zJjvguz5EOL8yRdxo5/Mg8N5IvKWHlVSLI8MdWLnHTqL/Aov10eu
rAT3Uuc87pMiqfSy1jS8dmRurnPqOlG+6Txz1K4JXEWePqca8SrceG0H55ECQLotpeIP9gA4v2L2
d+FHIevloGOCkKlPrv3eSGt585zt9cD2TrgsdCzdHCyquU4jg4daBjJzqFa7e4+uUxPIijXp++os
zGI9wZvUlY0HDls1qJ3oPMI/vXq+myvT2HzFILA4vNmBtg10nQv/T9LTF4+k4k+DwSGp17piLab1
U8gmIGWw95JucjEHmHwgtyUI3ESyjNtDU221zaJHnRQUeBe70Rrgzf8fJ1s6l5Hky+rPEkZX460f
rAJ2oWwDRtsOxbjrFUX66bEy2TSbA9tu1yckvBoEUJRzKcadiJpUNH7mPRVp1P/0CS/NqnNL8tcC
Id8N/jvaX1Q+2Gsz4kId4hme1TBQNhevGvMtH/y06XvgAACNrJGOokbeJU8n6ltp1PgWjWbD2Gq/
/qhd4eGNM8BBvrjYmDf5jMl3jfk/tJuNd0R9axmzu2h8Xy9ITCMTj+qij9gkspsTojk9/MmurVB0
JDDVd8y727Ws41ehyDshjIlYZ9WC3SJCmKZAv4alienfZrQfAfZ7wnmsREB1R3rNHxIc9FmUKUvz
O/iQeczBcQfWFuxq+W/+15NdpBedozBQM6WcsuEu6KRmyNP01/0ua0u58l7Y3i+WnPFEHPOXeeLu
9jdepUqc85uR0JHY5S0msa84c/AWlnt8MoPsZ4Qkbf7Am1AQrf0mH624/RnAaEfdXFfvarOyZGqR
9iBGjsLBQrgt228Z49Bdj1kqyfPQAXII1OlX4h1y1pCyPVitnyqu0MXe87c11zvMgPx1ZyOCSgYQ
nm5xOKZGzxYSX+f4vV2bQkCqAFPj69izQugFj4O2JUNV0/KCrW09R4OO2WB/FiNasnKOFIXn7mmo
HTltCnHEF1uGFgCzSUVUQRM4VTG/qlImw7ztdFgEhgmqVC3Q9h8Hp43voE7PxqgNCPzWRU39GZal
5FXliI/tY7OQmPVPnBt+psFuwCL+sMoLZbSzCmhpMmJcU0KPN/4qxp9Y0NUa/2lHMUGaHBx+m3BQ
7Ay6fepEyZkV+VmTWAphQ2z/267Al5FWEHI7+Pz1faV+FSLWAQKcqJ/jEHSzVCFdlWeehNApHzoH
7rFnoxUhrUv/5GOJ5zaFiq/aXzgZplBS7h2Ob+tjUzPq9OYHcg0O9dDR+htbAvfnZd68Xy3TZYip
JQkJgIKCuwbucBfDQd6a78gRPnc+yDet3NaFymmL3dAVOH5Hg932V8cv5Ld8mSN3myTlnziolelX
EE1TO/Xrsl2lpmxJbDMl3QLDTGWMEYeLRJco6IgqucHxCFACTvRfEEkE8F6TX3xzTp1yeI0h755t
pTEhpmh6FeEelecKvOtNOHM+SASdngMT/EE+CoUihc/3cnaDIRNaPslrQsl/VOjGgzeUwFV/pIVI
BT4bGrk9tY4cBKogRf4Ngad6UaBprE2QThvLb3N0XhxR/lulufRhmUg73jwUim1GTtR3AoT2k65r
jak2/Jt5mlts6LgZqIEadcHgrZzpiFho0lZ3RS+vbk4skMUemtoMje6cdYxWXqTnPDfGALrEPAfr
ulNU9sMMOYQd1LWLXoX8ORW0YOecIi/HSP3WKk8pq4VZSe/IxQWAkEnZpdQQtNx0HucMWOeSASTf
NCixCakdpt1BGNRkz/n7OZOwXSLZtgc5kzfBWjhc0WkUQd2YzQIcGmyxnQUz8Z7yAq1VOy5tKufQ
kDkbkFlcjt8pVhwDbMLQp7X1WQTZ/uBDtQZ0F+NtgyxTp1r6nmaZJjlgOQ6J6hCeCRow59Hg3pYt
blX5/t5QcOSvk3/uA5A+U87cJp0qUD3CwVTm3WLE/SYq8OhKXFuJrw3hjDUw+Vwhmhnd67Fpm+pp
KhhJ6E0NmA+0Lug1kw0PLvrKJNYDoNg+w7Vvlu+TVF+1EoEsW4DilHkIRXTYoncE6Xn74KobYUBQ
uQ8gn7mxVGdeR5iGhpYIaJaEpRHsrgm7d0ibYE9pTaft5QBNyisGohNFtjZU21hsTpq5kBi5bVS2
4cAlyWkClA9wFSGrTY6NJbzm3fydP+FQotVAoS6e44ldXHGiPJH4l1x1MXSwuSCZvVUJG69Cbzz9
XqZWDkWoQmrfkSBOcmuzF7ELNtn6vrJuMqdj9C2vYrUdIhhCK4HMH2IoPRIK6TeeCn43mtHDRj4A
VHbqzybL4tArUWLIZrtEYH0+2jFnPTSUR0I68ojvc5qkHBDpWYVJgRsZJwq7xrT8CZx3p7MLwlFY
/RLI2qDtXomccEkQYIEFvjSNaW6gsd6Pq5Dp4zboYaRC2z4FUpWGfRE4EdM47fEOnwMsI7TO/tfC
2eG2jUGUoozeofZYKZ0S0Jd7K1Dn4rhCbQgOXQjgzHKK6nFBn0ysRrq91atlpiQ7fN0GEMUiTDq3
90TJ0dclnypAhnbN8IJzjnZykS4phFhLFh+m1Q0g2K6AzVo2DQrsjv9SxkeKCCTRBtplKyyRQijM
HhbAZh7AW5qe6Fx0LyiOCi4WePplrSox4QD4JPPL/p5vR+8Kf02CFanOojAdeC1WBUMs3z3HZ/DS
rs+BfrLdMUgsa9sUf4xnuxOYcZkBKv7n0AoLtQsG9DNWx9kqeW0UDKL7A5i6NhfL3W8DJuX+6dbI
RxtUSORuvXoK3rHN4I2bZrelei7G8Y81WASVoi9vd3R5MPQ2+ZwIu9doua7tz7Xza8mkI1PduWBL
MU+lB/BfTItREcUvANxczFBmry+dR1IKVKLT6kjTWrWt9AGGk+dooDk1o+sP+UWenYFn2osMeN7m
+vSd6L4JC5QN7qm1UjtLyPyT4bzbpjo/26qoNkRlgTjTruPr80DCeIaPz4S1H6GJRBPqFJfrviEC
47XQ+eliXFptODLFueCHNyhYR8Gx4rWnavhbrL8Af2VIe7CTe85+DR7pwksPmLGTyVRHAE34hTNr
HMGRDp9PBzYkD9hEQR/OfE+/uYtki1NVJfjHTb4V2I71Url9RHqW3Xf4yo0SfkzLZsxXRLhn5pRU
Sub53UOCFAVMxmprmrIojZssXqwxgL/HeQlZIVnxtW9j+5RIQgbkJHvShLpfbjjR9PMSSUkqaMog
t6IGMHGz3mrztbKq6q0ANSENke0H+l4YqgRXAyd0idDS/HqucPIqksNk8THdMPjZycmfSj0O5tKH
WsBZ40kzZJ6KWSRCyV398os8d5YR4mMIFWpIx1K8SxqZIpb7OdQBbGU3VtXV3T03DFw/FeH8MCB3
o71nRM7so7uJDq93tnfVq/+OhlLSNUKruoE0RM8GUyBQyViFuumk5uKxTrKq4dN6PpjVdFw+z163
APN3BtX5OZ0gQOfnxMBzLJm4tokAKj6+t+u2CFUJgREGMwszPduYWTEGyrmUFlnV28NZY4ZlvTRu
pgiLXn9xH++9y5Bvs9qxHjEWSauqmosE9MV3dnND7LA5FHAL8GWFY23ItHabYlahP7r2WnOrqu/c
dU2pEuojPrnWps9lpjEY5KPZ5vmUi8A1wubreN4J2MNlRan0HUXkLFGq8aOV/G/E3LwPHlekQ2Jp
BmHzN1hKYamNYU5HY16L8vrr3hOcAmlsaT2jFkEM08dkwBqFMAb7kRlHq/dW+IZYYnlrYS2isHtX
zv36aZL16zGQEeuzDPoTgF2b64Y5ziEzju46Q2ICO9Vv7a3koFBjSx5O8NeVE0Mg7zeAqH5+rgA+
m7zcNZriw4Rm51RBiuTEA40u/7E65SQk9zdchsfQwP076CBtrLx8ockUklHtNiAXwOpAavXVvzT6
bbok41sUiqhOVaTiotPMW27auUA1Y4lWYaRFpwDt5GjZ7LncV1y3ZlGz4cTpqZeVFEyueG3NTxWE
JAmJPkyn/im5f0d0vFZNzQnMD8xUMYTA/U+DFtqQOjHz6Mbk9PMfu07hIJ/ms22tnUOR1YBo4hzb
SPAuYWpOD5ghBgkSYOtL79lLKMQcfRL57qLWCjjWk/OMcRXxGOqVWU8si4AtCTpwxz6zVJadrrNv
2HDZZPiBrWr04kdN2/UkPZNOGr+a9gZLzh/gr5jPuXwxR7y0JfbP7ekTwBZvAa1FFqGQj/sdFh3e
m6+y9bH8F6neVxh60rzR7DnV7g69M2poxn+loG2SjAWC1fveYykY9SuLtI224R3HcG/wJeFsGwga
ClrkhzgFYeeCNif/0FXAMXUvaup6unteahc1h+8wZ407VGIaMJ23BLQ9UmmP7OBeg4377ZMWDI+I
wa8tLSCmfQHHw/B43eexp4WHB1FXd35N5wQEv48ljkgBhbDwB833i8Ug4W9C4R+GgbVhOCWzndpv
4Fu1UZ2GA5cDzMffxWSIz3Wj7lkImhPYCbIdjzrC0uvkStYYFFwSb77akeRp6ObetNAjeDYKwvmJ
z2xCMHEDlKcfBj/i7SxusNsZrZeJkG7+Rrfr4utAlJPz/uM1y4ZPglNDByKfRVUbYxNUCA3LGiag
rFobfJaVLhK6o3E849R7c4wlrMJv9pX5cHfg7fqOXw/FceXZUZvIe+aHBAciLnxOSfeXF7nYQwpx
m8z8JA2LqXLdgkmQuchQfNfMoO+sC0yZc5IBBMK2zemlpwIbfg9dGGwa0rgvEU6tvvC5pM4GWh5W
482kz5augGJdmxhlUQn2I6aDINEEnAt4aP/i7gVd55p6EZUepMn2YMoaFNNBatLXMjRFzi3/bo99
OZNasy0wuBLH2mS3dZ5iI7Hm1h6WOc+/Kh4cITmTuv3JvfLBcHNd43tLOr2L8eERFbLZx876ckjq
Rd9klBWwK/2K5aRd+DGuDFdRRg+rqpkF5z1UqmbvgYviNQKbqLZg3POkyXW6pWzsWz35+GIhtIkM
qrWEmDSCANwuh0exT7R/moH1nAEjkQvMLZ9Uxn3KOEf30YPpArJr+5PGK0bKXUtrrJpqGKzbJnM0
4C7xwGgUJ0WH30Fjb1S+m//JSc3GX1ZhSN9YdwzDlwmzPUFKB0FfXRC0DzHAeQlUobaFUeEIbK7y
t9ii7ygMevvQ2odmGm7NlI6VmWPyeVk+qGQBXk2QjI1YvKrc5dZuVmeVVXmy6fIlsjqmMqvZPMum
9gf/TsRE2KWk6WBGvC2poYPCCIz0ZFIx65aFYw7aZ8S+lZqTGvBJwmnUeIDr73c1HPCk8GMIpd1o
h+RO/ipkii2XZz0r+VToqBv8CBV7KAoYtma5ILzuvJpUcHGscDKhlpgzwZjqMfwvyY5VekBbcS/4
OfFw0FeSh98barRaUizUpETKp+jID64rdU1JS0l5HxDVxmIId0EJeI5s8Fj5ayMmsJ0S10qyg3Wc
yn/tXbDz1P5xlCjH2cgY2hzgAzJ+4UJFwXwha2V+0edZ2OJXCPYLS56AS6B9LhiSK85mMJzE99Nr
yZOnD3+eENh0nzlHkpZuoMYg4Xl/gqT/MQV0SQZz7uyP3rOEnsrE4qa4r0eCRmnFg46YGZKwsg9a
arS7iZmOeb4F3dg+aA2xD+BojST/QkmFcqhzNO5kpHxrbLg42XZoij/iUh7F9Ew+nqzmojm3cDcG
cu3VwHHJ1JyOl+B5NA/CCWLUkWWDDVtq5XW3UxfHZXJS/P2GDCaPV5fGSL7q9QK3+HVWX1HYEQAd
oawbuuCCvyYVU0FzfoR66TlgA9TzHvy+YjwI1DhuJjhDAa6OoDGCPUxduOuyjTuRH4slXowJuu4a
f9bEOfM2NwudKR0AD5kpWimD5f08/YnKMT2e3CqN8+oMLHa/gkrNBs6V+RpZYrcWhewwYdkyxD+4
MF14wPXm/T+Hc2Ytx/x57y0dTf5/IUUypMCEQczarnNGMgNY9/RmzATpEbalj4JbhOzKFCgkbaVp
j5B2fosgypwkGDeJuz5bIHcq5mLG0fhgOWhXG6rT0bQGdDdZabX2S9+F3vXxHuM0mUKvBQztQWpJ
OmD8j8f1DXFlmUQRLvrgEhcpvRaRA4bS2k1ZhEjcVBEfCmbxHrFTxl5DwASBIw39DSNbKaYBXUtY
a9dCpjhn6N6FGQc6hYha9AEosE0nUxWB1dK/tZiTJp/sVB06tB6KhlHvosgkaF964/JOh/LMbw+C
3hmUnvIH32zsMkiMDhcmatb+yXA3LZ/cw+JmhvquDC+iNLK5HaZpKfvtarieBGIeyXRX1b9QWQN7
sx0Go41UdaURrdIyer/GajASLNCjlS6zNfBGpQSzNMD6JbM4axWarXo1nZglnVUHKgo8yFZ8LvXF
KWXRgVa1zWJJ5eISwxVVH5opZWVVuWfS4j1DxWvL1ySSslfNKKfBXi1/HBYjGSFQawFgPzZiew/e
eZBylrRxb1qKyLi8LeZ21LAK0vu0SN79IB3gfIDu2rCTDuNljeGcbxzqDJ+Gp3MirRgqWFLE4AnX
z7DSpil5/PwNO2jFq9v57bMz0OmO2w2YSuRyb7ACse/8DcIVpf+xkEtv65bK+K4WFQ0R/GQJXvsb
XEbCeZiTNrjGbstzbZHCkz9qcCbq5poct/8pot7o1fRknIZ6O5blMvy/DL/IAEyaGXJLXowBaYVI
yZZ5mLlSi/TnrDBdvbMfd80cW68gKhOfUhrAwSJm2NqjDdWLLrNjPZ+iO3nbqXpo47bA1PT6US/R
rRMzMq7jDE+CxGALxko6yOrbf7P3GSkx0usz8/kWqj73Lv79u5r83iNa/WPQHq5YGVG4B9qLCHtc
Wf14wJ03LVEPhJmv1ZxMlPD1z0/H7Hx/wI6eG7M9W8UrI2ywye0z/gdZy0XXh7nX7XbGyutXBfag
FEORP3PaA+EAQryezBWqicJFMgjvyZUKptXF2+adgtJWSFoikohlEBSuVV8srMHJl6Fazvy0lUTA
65+GyUXJ4AVGJLtWY6ux6pD8aG4fgJ1GXmDw7OFbz3Za4xYKY1RC0lcc5x1azvnwVnQC6rmDbYal
qRSw3kcBYD+ImbAIO5mV2ZPnvAqtna9NoTV0lKzG8VNzEpMyIO7knAWymUDh6rXyyHE4zvekFV9z
1yOmbnPEDjVdCmQlgki46Ghrba6Zk6Vx+WEDHt7VDSmaUn08vSUT0vc4A97g40rBpVO7AN/uzfGW
mEJrK8dqgDW/I4eVhLtKIARxCeqWeKRndbl0AZkUL5cOr2jjkxNvqABvlBfy10TSqf0+c9parheK
rIRPjhoOIG9QyjuCSUTHnGoGD22dZDmLWLHAh9dY4J0HEnMZPCqjBSaoD4yUtrT0VVc7Akzpj+AQ
vpXJQoAT9PNKb/tIABPyuoFtxTGUDhyTLrX4Jbo4hHRZU783fc6rBurk4eoh2rCT45PEPlmMeRHA
uWn14IX4gPZwGuPnZaAAb6an8s2T5jHcs9mLBBPJDOplwkdiEt3cjSTk3RRXZFj+0VZJRulrLcNn
KJ1wgOYL4JmISfYU7grkGnsOIdDHAoS61k57Lw+ze5vVAFct0cyGJbsfhp9vVkF+oMT5FB8qQmw+
pfSursYbxQuzX1jeaNerEHxd0jX/LW0hOhm7H4uQ/gNIVIzE2VMaSwfzZT+jsdkYvx7QDDE675PU
wUR3alVvUQ4j3PmhZqr6V4OqR/d9/z0mqFHvOOJPtwqbNaIzx9FPj+NRWJ0I4CS1d3G6FmujdOl/
vuhopYX2VHAYBRX4mtVXkQ/wGZLPU9c7dtbtmoQ6GcmCBLalyvSBqZn7HJG5Y/HWFCfLb2zmEc0B
/A+Ddw3eDaNDGSdxDsi4SeBGyw5qXCvhTYZbnEPHudtfhbkjEJwN7Pm+gM5oPYr9Rby7cJfeEMKy
Yy70J6JWV9EcHWFd8brG106yAxs84M6pRfliViuLEDgdHh93O+JaLxZ/Pwsg8/XfyyVFrUBC8C19
pC34KE6DnQCgXK9beF1FIkhXq5CoIk/CwOc56TiZDfX9f49S9YZe64m53lEm+ou4wHU+74shV8xD
RLxyL8xWKroucpZwSqfOk2ZmmGivca0vj81+1mMP/eXiSvptfnfQHbp+Uus1KKhK/btidKXu7RDL
PO+OtSdx16yfcDeM2CV2Bf0B4EYX8zEID0xAuygugRHso0t31/1VVhPCxnUA2gYmal99XVn4IkOL
mtl3zdAzqw1JEj3Qm7flsKC5fv7IeLHmaKbP9rKlyY1oOahayeRuAPyLjOXL+eQYldHPB9RskN26
rvT1q+Nz2/p3TLe75wKdq989+bIeVtRH1tI66gliStF3oNM6wmpstkMF2mzTwivYyEwZxeQCpLL0
9cNsbCij5uxUjSqkRDFnK51nGS4rF1vrm2JQL0T4gio1lX9gBNosDh7WfGJ0PY2ARc0Yu5xxnj3h
R48BZQw0fvSc2v5NG4Z8iuyay914pzwhYzfisQ01ugIndmgchgJHKTY4PnrdygASkybO1zbAfCeX
bq8jiRFjK8vaiNdtWxB40kyTw3mc3Kixw7YAFUosai6CgkqCe0WskX+oFa++tpLR5fKmpGG4LRDO
U/4KmkDA+P7LSDcM4ik/Vh5NvO2UJFzB+hO13qHnEmDcTvo628/XflVCYEVfcbqjrHRX3bUv5ZGt
9nEwdJQkGET4LtD6L7eBarcWZ2Fh0S6SPqPB9DVZeJa1oHE4vPAc4ITDevg9OzfK8gj2SoZqpS+0
dUtQRQeDwLxXyr/bZhiY0xt5sFBlTPPZ+RC1KyS2iK4N4PQjJSyoj7v4PDHQ9NVe8TEjSRJ9qRA3
b/87k4uYZnCSzck2VCn2oyTlKuTSQs1zReyMVZlVnlv2J9H2HElKSg754QK0SnOUbvPOV+KHD+1t
MIHF6o2NjzdA3tsXJHJF8oc1Qn6kUVk72Scwc+QeHeWtnq24qA0qxWQSTXSQVLQ1OknbBv+3QNwu
gEi7lbbesLv1SSHjfYJjQZRm3jbrowOU0j0aDLBE/W3ieIqz+HsjJJ5gUSbtOLH7BmgQyre+dC+X
9RV4gYQ0WXvvlRSXnTxnf2yFBoujxOUaq/ncGIGABvWu8dpwwEZg37kpWQhNchlf+FfQYLpab1QP
cm+2Ud6f+gNbiHnHzFe8fBMuOfj0fyhcpJ6D9brt6wQlFfrLTQj5iR4WOa45dapH/oVToa+LvqWk
IJYqNKbjLopdf8XSzpDfyzub0KJlBLVS2Ncg28fH0zieB1Olt9w+vvq93JHYJEvHDf3wV/l8sE6a
N5qSJa4DlAEqjNFOBEwHnw0Ip39HYoB1n3Ix643S+x5PMT0a0fb1w3rDvsPEu9anmdSfoiIviAne
tkm0FD0ptgH7Ad4JRqnuAZofQ3kh66WjDh7oXwBx+NKGGymPZ4IeHzdEmcefBsLNAp2eQjyovhen
cHaZkukLjywI/FSh7+9mWLvV32SzBfiFWYeXHtnoYmoP8AWjOHaHuu7rQMr5lpHEpDpFqkw8ShyG
Jjc6+6DOpio9CXJn56lgniE9HTzXO+2JgD3LjxB3GSU4+3+J3f6ZhJ8i2sJMvI1m0cb3DRE/3CNl
gPvazvro35y5zXB8PqzydL2i3rAE5TMVzimmToQJI2fOozKW701ok5hseDbuq3ma4TXA4VqWHfUL
xvWH7YUmKvES8EngCfpVUBc9EkKcCXS5GO2+n6N8b86CdZ1PSGdsbY6tQAy2rUI7Qsr80Fr0DGmk
lCECfqDe2ilw4HdO8lf5BoK0KPrZdKKcYR4X+/JaAmgQl3sFKh73EVHofCaNl3yoirfLgFC3j9ng
ln8nYpZLNq0IInDUh1Z90fRMYCr6pYOds8m/74soqZcLwadYnIDngfpvrhd8oobY1Y5XAc0uA4Jz
FURcDDHTYYnnu5iXCckdQSZpRaBRvWLP7wbCNsQcd/hILBhUxpXV603ATi4cRYk+mltmhSN2q4m2
HKOzlnJS/u63SlOHOPuHMMw2/chP72A/UBAKjfpDguJFsPQ3ozr9LawgAN/9KvIwVg/EJCxfuIQV
q6uJvjajv4njaVMxrCnNNQIPZQxZj9XQtKOI9jrC2UJCAP6+dNtp3CxAIofwXUzbVUu0FNpgl21j
WGlehD/7hXguRNWFvt+tozpuewFqz2g6NH4l0HD4FqkOIW8yHVa7WmsnAWB9wLVx6XmpmdUv73+c
Lz2mR9T2iD2c8u2Jus9aDzaH3/1lExjcG7J7AEhKmYK+9cTwpS3MbdSCIMyKLP3riRGqVlC5pBUD
vR2iF5FLdhl3tzDTpJAE7vX/kFJJnEnviHt+GspKBqEfyd0DlBvTBgBOosH9uvI5iKKc4RZ31ycz
Fni63MYndthq6AUxh2sUgPtt9iFmjq/AVSWDGjPdmaIZMB1t2XjV0SBp9E6ppl0fi3GQiWXIF+At
tigwzrbqZU1wuoZ9kA2GVbTUMy6LxM1rXzVKGrGdUD/9MrZ67F/use08KpW5KzoXmvwruTsLYbTb
0Qr0azr+dgLnCK0fNhRlaIx/KyysszyoJhS91ZYS96htm+nfwl4c0tmzwtgw6GB68kT75HEF1mEk
h9ile3svJgg6l50KVivSxI647kLBKfkeEc2tOKg42byneky6gyBkcChga9+wJL0h3NYWWEEhcrFa
2bh8G6IIk32JdpAH9819IfnlWiZSPlIGPsipzkTaTqICL4ekp5QIIhD6S1RR35N9sCAo6WhrJ9MA
Iz0gAOB7fxHFN4ueAeT/d1CtepC09D6I1tUdx28amBf38GNwKZgybweAOLpdi+CgTkIpXxT/f1F2
LQMqQ0qQ4rEPvsoPbaxn0LWBEzVLQ0LcExwrqUSY1doxqiRVkr5yoDdEeSKf0RioCNhPnQjyUeFW
a0T2i/r65mi6wocQGrUlnCp25j08XZbBRxWQLnQwLGTxQgYLdYgrwSDZ7th96Np2aprIu1PYOnq2
VWB1kK8u1O/nTdTbSI7erw+5s9iUwbq94vfwB4rexZKJ4NyO7uFGugmUHhrMr5SndiaMLe6VvJ3S
CRExURntxxMu91iWVYervt5j+8LBpk44iT18FoTfeJQJPyXiI7LX3e2EWwA2NOoh4/Sa9x3pNrqo
cuAmqRBhQwZoM7jgtx1K/ZyNprNj7RmqzLBH7lkQwf274w5O0NhNATXJcA9AkvD+zG7aS66wcyiE
Z8b3w7s2Jz9KuApmb6i0IWRw6r3VVSbLopj8tPN3x1Pfu8JL6zFsYDRQtfvDVcNSQJWdDwPydsMx
fGTZYzgjqIKVgIe4sB8HqyRzs+2iTuih7MQdAHOIgOt2LoqOjgXL3AQ9v3AFIDwa/g9oatDJkW5R
Pdv4T+5XAAJMHYOEL4ItLULQRA+3NIGS/k5Tji3f7pYiSpjiJc+j67ksj5JgxuT5PU6bMm94U2qn
YveEX7iZ/ti8fWe9DLVrEamk3WN0+l2io8avT01M653+HS5oCPmgQn76PNbtOPuyhGN7lrqBvT/C
W7OHt6lbvhS6fJE3oDMomuS/qv6p9O8dVycKkzi8fvNNAElN+b2GXQRFbZ6PN8AQf2nvQLPCbNfQ
j+3/UJWX1HvTx56gBCHAjCkIltt+c8Zi9I+FqiEbu+fhXx9q/qtONIEhcoOYN02bWpH/DqtKjP9W
gN94u3c9FVrM0aj0vP2TtMy90f/VBXQd2uq0AkZRh2cjwSO824Fa5GnSy32WJpsKgv1Y3Tq+3Id+
HP8mH6Ya32VWkMLuZDQsvbDeprwNhnRDddvYFG4K/BXHFHlDtDHJNsnIpgirW/cIlrIBW/t+9dAD
VjMhXQ0X6iZNlVleOmKmZwMAdRxzC33Hbyw+w/RAY5XgQAcx0ukDbbEB6MwIK04HaSt7X2extR53
uALsXRlQZKQMy4VpdEreT4wlgMBmTAJX4v/WrRgruDkjfE//nNBxGJRn8mXUptwxAyC3VDaArUPY
3mwKZ24UfXnGSwF03tyyvydmzxpE9O9f6Mx36/KkZQw4JcjunVngkrjbw8Gpcms5YkW60EpPdvsD
MC9zVT+DVheuAsK2ECpLIFCA+xGQF3iN52mLHiEvn4vdv2MGKb4wahyrBDn2y56Xo0ZzqAHhIRJh
26lCdXYBYK8ZJRBonUhlBCOLtQt1APQVmqBJeRZxpSG3dBCeEcD8n6ZwZk3IjS6iNXW2TFKOswk6
7ik3r07seCTbcugCizDELjUdDEyDxcR1WiLynbTYNaHivps0ghACcacQXnKrONZPK8D9ZoCaPQfs
MfhFfN69Q5ojb0/7gRqfTO5DQLrZrFZKCeI2Jdy5W3DZkTOVlvzRjta4QvybnDTPgFRod5H0BnTE
5q2oNfI+U2xvM2FMLXveSb4Uk/YLrjmYmmPI7vy1n8HXN2Znw5vJAszROg12pydQMvTMSoIsK+eA
QiYu8RK8SwbpQtEyvd8aWW/l+r69W2lYePAp/lyXFj3H/qLPEBJOehbg1FThSK/fMj8eruv/Daa5
dHlAD2L6zcAnPsYhp2X57S+b7CUfOGnKouMXo4PuwlRHtPxwyVrctgPIdZD661gH6m2ms/bDucqq
sBfUGH1OzzIxbVbzol7tMBebPtEdc+UdePsteW/nlrgrWe7RKvJm3BTqwutQh6m7BAhG8sTBpe6g
RkiIgTOB8WL/C8z4v4OgzRB0EQFkk7dmRa5Vrjh4bZYftrhBT/EIy7ncWG7hmm+gcz5vlCiZI00x
gEe8TT59wAXQhpye1g7x8APtN1jZbZMWoh957UoSNL0rgNLByLxKb2wGoRLG3xRnlAswyuzWNfJ5
zN2CpxRsICDJx7Ps72DRYMO3A7CdLBJECBbnmQH7BQb/p9HJlR3/wWQ02CCWxpMuycfdZKrLMBXp
P5F+a2KcVg7GDPobRc/XDa7G5Yz8my/gGp+ptlsSJnaYjUnR2nAK/bE59EljAR+mUyvQzHCv9H0z
g06hz32rH5cI+cEKXJMGO6CxtZDhsAqBTzqpO7x2tSkv5hTUQhfSMxsMo+UihJHkQhTcJcEsv0Ou
oGFZamQmPIkZEe2sXY/9Xqj6a5ghExTuoZ2Zvrc1yXiGUXbWbsiny+geYQVgZ5X0HYScG2ePluKo
cwZsbhxsB3vzdqh99OhWEjtD2scoJO9qU2d5dmge8pALdvkKfe4ab/j2zrlhmJZR9/K9uvaua1iC
1PJHRsRd/GK/11JV37N6ufOPkwS4e5Lnh3d1sIQ+IVMQEiRll50BJC8kMk75Dj1CPg3UQV4fd08b
2n9JJKbKITH28+8AuE4NIa2QJS+EW7bv2B8m69jC9OSJqmc0//nnL2qJkzTnWcyyo5uWehY4PU4l
WWXs+WIVBX8Cpln9QD8EhmOJfpQ8WdE1zj7uVi0ovb/fYIqtqwD3ZVPtBcKeqIfvQmxfw+UjM1GT
FR3cAI8o09ClqlokWT6fWJtLXEHTYjcgnm26QNJMVu++lzPtL4b6ul2ZFwxP4tNltMido8vTm5Wb
YPjdsQ/YFVlbw4A0FwCQLqLo0M9clCMdynbm99Jz/USR9NxpYAOqZK1m95zPDsCkEmUybVcn5Zud
p87jZ0VUeUekDDFGKXjkVcEbnqIxOIR8EFPelLy3t+7+ow3xwmjbJdnkKeuplaWxP3FgRaY3+/Wg
aN/+hSuJJBGCFXj1Sm61gZA+feutq3GTf5tLX9uYS7usOLPphR/+7zpzeXIbnc0mqH8VrVOTRJws
UaItCoWZA7dO2MeX+qTWgAnOzW1Wpy5bWKBMs2uEYZW0WS0r3CAufA7ziyZNy5TIAja0jDW1Q5Tr
2SVTA+t4dpP0+xASoHp2EjofVKBopc6TN5LLp66bQUUT6Gy3GJ1J1xnZFhGpxxeml9xptW/7Ys5T
5AwtHuMGPOKEoWGorgFGardle73/R6WPMP/lgS7Nt+KpfxLf8Hpn/w5hevoElHl+TbSorCX2WJ5E
oYPb065mmI8zBz3bZWYMcHgl4zynLJd7f7Br6RQwn6CwqagwWG7OTeagu9j0RmWLfAfv5cbahD7l
48bd1OjgZsJGRllOwaA2PYlZLA3s2iAuxStctoRCgHNfGNp+tGO6fDRL5rDxlQpLBIu8Dz2fTVlx
sUBRmF8gNXRjujhNayicCdw2B99S25SioywnTcT2hjwWNgB15qLewRHj5UEqYn+1937g7hmITrRq
dyo+EUhCRomj7gyDhziWFgeo2+TCiOCIJQkC6hNFxrXjOKCw3MVsx8kzrM7AALVB7QgFDXV4wyTo
EhfVHY+qqH3pvbJ+D68AP/ryvOrU0R7RhtXMhx1y5IxJu4n+AuxqamswRn82RxdmckNgQ3ArUWj0
UB+UWumoajV2eq235lviiPbU88ZkiGnVxAAKYMjpbab9il7f+yEkM7X7VVuTjj7pYgEh+CfGoFQS
ELZ802qmF5TG/BjDpnnrFCNzuzl1R7Z8BgoR0tszGa7PAsHVEuZoNGBQTHaFuW8/AgBBDiVPpBz7
mSED+1v48U/Akg+aYzUA/KF1fxGXuJXGVxJOjRkTvde7eAMOrCqHiarUZsh52NsInKglis1LGzM6
PFj54IrbkjOnilf6r/itYP8fP7QH2mw9qz+y6WAYGLebiouOrbQfha14RAOvAVqv9XEJToIselXg
cr9kxzL93HCcWcrvYJ+UsCLsviwgX1lLi/eZxEwlhdgipqah1O8J5Omi+6UOeygtELkerpFqQ/AQ
wJDygQrHnvOSGjIDFGFn7PXRwEGdpGsZ41GoLROqV3X0C1623sK6JghfPpe02Wt1AAWf6JwATEvR
nTpVVVj6C3e61U1zGTTzcPebJsYg84gcUTQfRyqS04+NrC8yReghXR+DAQKxwnDcWErxb9IReMvS
4A3fmRWsTpEkwrugUa+BrH9QEWQv+JjYFD+SuDr8Eyuv76mXzrF2fS5leazUciq3sIDeZe1qmxNU
gzQVln0jpGlkV0UgWJR7vDgnmA8sViMZ5VWhkNRrkCS0yYB4SRGjvqmqaffoTzRFwr/8IZvlCNXw
YHtMRWE1MSR1TRnAKjVhCWVxWdD1LFICbJEePwRDio1PhgrI+LUamFuWewpD/HbiYQuCNkuUqFlk
wkmvqtvSAOfIw9GyUTk0xunmqB1yafm8ryafPL33Lq4CgJfTGzn4qYlFqG2LleO40dZPcpM/11ek
PZE+JAGe66CQpglGdJ/QXbxnn/k8X3zAsRV6Bw2EJdWCCY5XSujTIDuDXNeZ+25ufJUZu/t6RPHr
SybRwkiAhCRHiVv50L16sHRrguebWovGBmfTaDDLOdqMQNciKvVNJFTTvfN5SbN4uOEoG2a7QlDT
OCulNfEZdUVmPCPGvQDDirif1uHwxMq2jA+8H6asdMNpD1mVCqZlSRZKqOiIZDf9EpkbkcfheGDK
nIRzVlCjLE8xoZlzSPwrQH0T8NasIBCn6KxZRzgoPxBXqjTPtRqNe3sUdFyPV3TV1Ibywdxt0CIB
LcrpFQ7ceb49O+JLfSC7La646pQZD1CsMBpw9rA/cQ18Eq9DIS9atx4k4SULgQmvGLzAZkHtNErV
ILX8CpIUoggm6dGA7j58SpRCprs/c2NlQgiGjhXWYTBvThXsNuLMjGflpUT+jWLUbo7f+RiRVD+d
OtCkSZG7EyBbkLh+tXfHJXRTKdPLDPRw28ArFp0QJDXAS6zVXajaox7y+7wrLLM9nnrNYAugaQrZ
kTV32VtsmvmxeE2E2dwHcKSFCLutDVa2/Y7xPHRWMWr5JPUVx+bnEL8GPZM+/QNqvaqpIhwyOCKR
Iw1Xlt25GuN81uK/njkNUhP3SG755XgE2kEBtjqsXAofSDY15Hm4T4tv6hu/OOoYzkTDGscW+0Xp
9CxX9YcBE4sc8Mg8BgQyVOYqJgfP0DKlzhLZg49+rCEmbqsIYzF0gErb+Pi8jqf8hy0Lq1yt+VTD
3RGbQEhK7V7Q1xeU92HcO1bGNQrCgmoKtTWj0AmdJ9fOcunhD0y6kVzLYfceBZV76nfUlY20dWEo
WjNVaHqUgTxaPq/JZGgAhC1UErX2egl/d2P5SLWUrxQZEioW8n/U6GT82mg3n7lKI8HmxjlFGkfU
Z/4h1SovyS1V+haGebUMMse3uQMGL7bMl9X2HKjYlM57XpPuGe8N+ha0bL5ZC34TH3nnVl181IU5
+S6Nfv1oQXPrYFhHgDJwm4MXkWVuJnoGgnUsLYxHiONcWbPFUQYOSPMx3MTRFsmS5/hsFgxYzlTh
rFSSjzAUUvyBEzTyLlX+u/mYpGeQqnMLSU4vb4Xv28KnrQ9TxjjNxYUHUJ7ZXhY+hsFZm/azryy2
4xjyK/pYHeDQXGi7V++pk0tWq49DvFo4BzcPuGyzOjhEv3J+jxFCDohwSz8xgz2+gjTzvix+byz1
M2kWeQexq+ARXV0XLQlNZ2rTOP6HTVeRJ9bsERVcGl+r21vkd+984DFyPiT3jOmDtYIH4pUJ8tWc
wq3VKLF7oU5lrn0RCbU7VkbtAgaV0wrE34wBBd33PrjsJyzRNq5oGZARK16sztPhjX6L3cxNCjK7
LDpAyHXlp2+m8x7q+l2+blwhkIZd0aPFfF2PscXAu2zS7ta694X3AilftGgQ3ty37t5uCNY9/L+k
C8maCNEY5aPcXJehDHEeWJoQYdeFf4JX4f7p15ZmAsc7Uw7f7Cf8+c+cbMwwK+7jXhiXh6/qfRNF
3HJqBfDo06VaVH9iFHLECBYwWPBMfG0bq1Sql64iDCN0s5mHoK56Buo6DKbWKo2eks/XOiukc0ZQ
k+kvLe1i3GjHDZ+sWTDlna0XGTU+YHl2mqayT09XJPErQg+7o8gw/AnzbXA8U92eptNyXvQEz5bR
E7ovoWWkh++3sLuluODoJBGYO8KK/XHCLc9Oywh6p7etK7HjFkro11nV/uBLNVsQ17o6FX1ifYGQ
AgS9bPH824XQtRHKEa3LrhAkzIruQ0D9tpIzeh1jdPTY5MXkugpd/GAyGGkfr3Ixm9wz72qnABDy
I28oLq9QtV6DqZK1IBOJK4YrPm+8wZi/GUDaBbQpu1FVUx8qFBV6v0JvTY1Teh+wZMF3lBxpQ9SU
RkUfLzHC0mHIfKqzIV1ml6r3rBjWXxmf5mwgIseIsYNCr9AcfjFJsw3rE1LmZ6BP6X007mFfNhTe
6wRZD2OOsfDbc+E0kInV2Zqb35Dv3kuG21MHQL8D37r3sf99ijMdj0wgw7GR5jRvPXNIX2j9oBrl
+XBLgJyVSZxplojxtbKPe8wp+sMF0/OSZ1lUXDncI5CAgMtdeZOmXjgCfvXCd5mP8P7kvPtS2cyR
BZFam7PJAuriogMCVTBWc2bACdQ+nfLfu7+kFlu0oN5H6McbD3CAKGsgu7lPNwGMcYx9V8IjiO2K
oSLs+om38oY0Z4f+BDoBQnlnlGMSpGS/CTCkxpv5VknT0Hiin7ypnTUXRgyTVpBtdvU6c9iGRGfd
bvnXSdEL/1xPgRE4GbnbG/c9HKfs0Oy5Y9K1SZGK5POAd1LiQhriEE7uvuSvMiCHulQZitUrY2DW
yo5P/HkfS7oztMn7agZ32qwRvwgFCUGwoBEBOQhi3Prm0ZdVusc1iVUDVsGik/zT4A00VkTBsLsg
aRnqfnXR1SxMXYMfQN9N2yhezlnMeQ5dVynNw6uOOA7QT5oGmWV4kEDKz1IGjRIqxKGNCK4VS2V8
TT7pb4AxonGQaPnFVKQvHUIMNKGZlONdad8Oa2pSjK34AMgQS8JfdZOhbd4HxDEjFPwBnckdNIQ5
JooruHZVGD73qmcSC6S9nYYN0717XNrAHuotvLCqfcns7r8Hxcqwev9+Ylu2emF7ZhRb3E0z8DHZ
kSoYBHpLFRk51cNWca2/YSo0A+96rrmedzJuIBo50+OzL0vqkkMPDH6Y1TGC7GctOoNSzu9GFAoH
1AMpVG+62U6oVfeZGykpwa14x6Mg+KBQDmGFAQF4ibTa5Nq0NbwoYfmguHrKMOKOn99oj9q5Cpj9
7/7sT1xB/h1Cm2ZHrU5b3F8avAq4P2VUoU/ydfCtLO65mIsp4rHTTwrEUrHOo7VhONTMOCPZYNsr
cyeQ6Oz633xomi4aKO/0HXkhAL/pFk6ahRaX3OLCs8i7kdG6MGOajBD8Ix5f1WR+wgnzJ+Bnlbn5
s6fUvgpg/Bs33tZv1L32PJdZO9fIxI9sKldQv6kbtXeBfmRMsBuGiY7yHuMpdCjV5SUfKzpCSV7P
MIVLdLCPMkXX7eHlAbxbe08vUsRM9qtrr/kcXHQMOdfRl986GZZl400PcEU6t722aHhmm7dV2iAx
NT3zhjplls3+HhfKlxm3gKYWUDLkrBNZB62adIfRLZx9QKzX2njxkd+np59q/uG3qF+U8YO2dUsx
X0fZVF/zdzq5FwikjayhCGURdBhVGzuDYCCmH3T/b0yyss0ChrWQ8Fc2KTFs8T+uJHWL1WE/lian
OurwEUr1sgH+76qrJ1uGZUP0nasl+NXk1w2A6e6TKKU7EFOTUD2lQBXh3jy2S20AMr6ZDLyLwzvo
MYcNWLvcBjn57t1YlLcwiAZiZm5S29bhkI8RgqfPzEgE3EK+mEJIGqz8W+3BG0IHFcuGntF4Ayc0
LSZvXgtCZ+olu93YCFBvHliEV3zPpaV1tHUPw1LCxwehbQkiuAFBqzdKLHm4uYLi0mGM+dFH1QPs
X1fBPSrrKbjmuDUDrCV3bCk6UBXlTvYpp6EZ17oQHk3k18pbX8zMlBt7w2vc9XC3tG/wnesiy5p/
OvxeA6P6Vi/jJnVqhXO8oqjBVWiLQCpjLh0zjuHPwvTWxLRTmP/5GxoWBcmITa9pfjfc4rh258Aj
zgTXplA3Uz/nQC2d4VaMzOYOth9EV8S5wRdcNVeNhSyUIhHz6GrO+FPB8dGGDnRmD8r9rUu1S+Bx
FQTWsVGpkBnFA9pRl2qx7WSB/5gia64HqeD+YMynLHyyltCdtQXndbrkKDZZUY6xVgyr7CCmKVxF
xn2kKB8q7xlp2vHbQZYuSn/YPfFtkyufXp2Mu4xtWQM9M6JGMCN3sDwMHPGTDE+PVVcPrjXf67HT
zo3i+yhGyp3POiNT5ImLko6nubg6Sejo5h9sf7iXH4U930j0K8I6KB1pEib/RQab8JXiFMvKtqvv
2CJl9RnwlOCh4UlvuVKZ5iCEbZLAYIOULqRy+N/2oTgtbe4xr/P8BLG40yuw5q5qmY62OklIzRkk
6cvKPPRblG0a7vLUGq0Un7RuCpqxD7FToeRmBLQK0vljEpAHK2XkvO7DTryyC3/CvlP/xqWJ7nrs
E+yGzEOpMmF9nlNAJA2ZDM51e/QCTZCqvydC9KvQnq4PYVCNsAdE3Ive/z7p+8c5eE1TphE4+JfL
shR1SOIsF0mnv+u1jU59Mc8h/es3nSxQl7e4UsCb3dw//WyQ5pvzmy9IBtD4luokjwwiJon/B0+x
673yl1gLcIn8JeJFffWyHZRzndLdWwjCU6C/oHw8DAZGu4TwXBXNPhMv78LvmHbDQPwYQM+YBEII
S6QMVQqwkJTBDXLqAKpR0t/FOFBGNkCCvi8Q/lNay0P6rJqPMeKc4kcFf4fkDv9QJ5i47M8ffR5H
FYUa0CMtKQh5ot8T9fhT1IWesrGUPGz0/YuGbGcI1hzyjcxs/bpXNOeNY8kqI0+Q4fZFqZJol8CK
49YYFDKV1cMMbr4M1xQ7wbMoYyrdSAcOPEdKAyYQUHSXy9JGK9jLcdy+8OPchGirN8xoXA+ZZVfO
9KH0mv8SC2a30FhZbbih6SfUM0hpGBQ8/Aalcsi4MNIckFOpc0gTqGeXrg3aYVArypKp76pMun8L
1XY/vGVMDC588Pw4QWgXgW1ziwG0LF95R1iYdd7rR9mOOVXtpXctdA1W6PL5izKDiCkEFWyDXcUP
XFRoGQLVW1+AZYpCSqO+ZFBWjNWRyJCu/Ua1P1BCpNTbJ07CTgxArwTzUjP2zYQhuI2ikC9GpTuk
UiDq5BYylfRsEwSPWaq8ROIMBJLhZx3zeS+IAol/Zrni4UprmN4EoTR3Gmkqx5Fek4Rdt/3vEg3i
aeCeo1Rlbf/w5QzIPQniMDp33ePewDBVXSIUi0gJy2HdZMyQRSX64CJNQ80BjCK3QP8tQsXcQ5pl
nvGtJlgcm8UUNRjghKL2YIowbhApRVEIFfQox+DzeYJbJpQNI0VF4VSb9DSkIvzVVcxmjUf7eakr
FZN1YvTW40wmg086xAL5h4Kx+IGvw0CFainqzwKX277KDpJt49UfUD2cpKNDJnm3FEKGJmNt2nHo
lAzKLS5n5d6osylvpTwgBqx6NCshM8An79M3xrWgwxjbEkZOmWSczZjgOVfir4XmEI2EIc60J5+J
mXkjPHMlegSH02kzhp5AGGAl77Ws+NXACFm9t9/8amDgVyxjUt1HT7PTJvZxXJBJUWWY0TeWeafc
+El1Rb38xhObYAx+nhOYUutNmE/EkUcK5JH8PWkr1bKV6eQwrKyd0BO9KETtX0sAj1hhuGq8vkS9
zOmJZJlOpiHjlEBJkDnuOra/ahL7EJjMpMMok+XcgGV877zd7gPH2KAk3ydxRIY/oyxeQl6+q59I
SetFf47cz72Kma5a0lZ2QPsiiNqDwQibJi7w5G7VCUrCJfZNG2QxIVdQMMWTQXCP4xnTS6ZeqZVl
afqXpI1jhN/xajabPT4go9gZxHYaBC7GBWdwCitpP41FAudoJfrVu+qd5cgZlOs00XeabTX7HBU/
TDIdL1/M860qCX71zt3zaqRA/YI7/HmtvoDoH1QgeDQ+V7IyYWoiFkAHZ0IUrk2KeeL+vEwuHZtK
EwEiuIozTu/gpNDv8el8MtLFxgba9KY8l+iE6x82/YXETq9FBGVY62GGpbXeHAcqa2XLt9+z4SKa
viaDC6Sg+GvehV27vMAVA1TUikmYhYWGGlf0aKn7KtIAYsAclBgns0JMvMHsmQvHgKNhutncFleF
+SBl43hgfLnGc07dwpZScnvl1CJtVo8nTSGqaUwzhWbZyDf0/rMxsBFlCftJa/4fJuGTOCFsBXbl
hGohz05pFK43M3X6RrJlv8EyjJT+2ZM5+jJks5p8OWig1nkgqZGgCcqDz+ln1xnxhHeT8zyr4JTk
ypaop5qBXQgF3dvvVSU0WrTHk9Z3vG8XDDIpHI+f8vm1G2kJLoRwTKy5MocZgCcu1Pf2RsjDQ5BR
cCUR/v5b9du8oYR7KbUk3bQ/GUrKaByA3NbfRGQ7HXy9eWb1pQVyxBne+70uDSNrjsAxsEkO6T//
IA8fHK8Pc3V3h0fXQX6IP2P+o7hECCYJdMs0Aa/FHC5gKmy+5HAw4gN0HhiN1u6M+HeDImn/7npO
SkOfhYsVYyfMBm1dxjwry5BY+vpTFY/CeL1lkJZjO9ql3G38b6mkOn7zJFXJ3ZtjzbpC0ghaHKdb
2C9hyudBU4GMv1dx5FEUzRm/H56ix4Lvcw2RtTKcbbhiep3NdfeqRc1MS44eAQo3AgF7zu8ksZKG
m3UTN35v0NwprEmdE8Vu6DKh8xCF1BVFPXm/cjiD0QWoi8Cx/W1QJJK9haqWqXzeoMKM4GGqTwBF
jIfMgL3tUkqyJh0EP6irlQtKBj+3EiqP9Fiey4cAQFqWOAYIrun0CT94xCddcbryruBTHjk5566+
oKkDe+mYgtYIyod6cUwpo4rx+hyJ/ll1Z8XewJd5PCou5mOsQjLNbO11z5nJ7daX0LaARcuI4Bn1
j1BYHNMZq/SG3ou9pokfpCJMfPqFLoco/rXPLr1DfVygExS7AE7q8hBzYp4yk8/E3MkFcgO4V8kr
bH1EEQOWZb/aj4TBk4wkvbYVSQ2IGF+C9NQsSc2vETKbHpnRiZXElwt+HzU6Svkx2zTEGEOFIwdZ
G4gBs3aLx2n6t9scuuJb6XERQH7Z5JWhv4EpQQoZ9LJJOZjEtQyq+S/bartO+AfLOJ13nJKUnYq3
TCbptylr/7+jwkUaF8NVU9N1leCla9f0yQfASOnJriPgh5sa+iuiok7sTmDYV95w9pnPyC7H6Kos
LBHnOQ5tx+YZrOFdMdWjBdFQ4TRMhbQ2Up9UuXeMkQZx5YUXoNTiRfofp14FWlUgEyE8mCa9h4Xm
hr8AVRf2qPmDa/DR+89+aQkzIaYxV2UdMf3lmyc9csUhIPQnPMUigSZuWQPpfHRkIJG9ysBgbGeO
t9ZF93+SZk7Ou4o9I3Nqtxn8tFiJymK+xdFP1jUY5xTEGi5u8n4uxPsiOtNx+AwLoPWa67z5V9tx
pvuNbsyWMUIPLT8tWiXLRdksvmiaxpkjzGSgEgbR1LBzbci4Lm7SnF9Bj4TX/kCzdw3G8+NRb5b4
iw8dqeyd/7PmVrHISx8iedGehsYiQP9okLkIa3BwJFEzc3ZBxcqVR6aM9/A2TaClxfNRQy9TKt3a
irKqnSDiG8LeGeOXNqoCOKHaezQ0Xq4vtOazOGIJ68uh+Vf0YQ6XALzLXJ4YkBKrtbWTWcEZH1lx
PXaHcRMsyal+t/kZzY8WExECmY2KPqobHDuzH0ablpZ6k/Cpl6FegHWIuNUvx6CzzcHEq2QRmuCM
iwAFU9ljA/1XweYAkcDy2U+qOhmiPv92h/FDBqCAfBj2XZVTmPBgpmuuZ75Wb8JdpBC7vLf1XRvp
uRvVpc4bhSPsOS+3Ns7GzuVLXeGc3Fz1p0+BhMJfVAA+MqMpCs9nP0rIHn7mfZh4sikk2dazanGQ
3XvOjdq8w7wgp54vXbKIzzVu8Xrr7nx0yfS5hVeSKqVinI9uahYDbspQ7EEH4w5pTQbnsU7ouNXy
M9PWn4eTig+oCFuXwAea/TDTrZ10uQaB7cwmQxrDTkna9/ozGKdv8VfAkidO5s8e79gMtnlHbCdR
/PN/U97Yw9NKLMuW+BNy7wbsB1A9nstVhG2MUxNBX6PlCkAnpWKI4s1JCDitIrqjG9njznOdhfHH
12/vDUCnGnUby4mdfLBfw0Gj3EAXmc2IapXgQCRvtsMdI/DiqAoJd0wQctU3yPiVdiV1fLwA0jN1
BrlPw1lY2++fEd2hXYfFT1kG46olohrL0v1DCuW/8EnYQ0MzV3NOdLCWJr3GkoCMgmY9IWsVdK5i
eNWCQFZvbHR+YDrOULGn6G4Upw723zzihFyFfN2y/0ykcOps2OCiP45sNiBoOsYxq2vAZg+roQVx
yqHLxRp4MDSBHnkyqFbILDdwbLLeAhV1oxSKVLSpti2zCe92xkfUE1O0ApDgyOBKJvXoZGj+HUjv
ck/6rbzM3eBaenUe8eT8zMSTBeJd7XSQ2q2R+Xa6Mt7gnNNjwA7sAhuPG8XI8la4vEeDPYo7/Arq
S2OWG4sfEmtPfaZPq3FUgAWbgT9b1BeiSaT8xUytnLFWKtqPR3QmNgRGPaS6WuilXMxtJUdA1RXf
xec9v3Uws4v1dLBEZ6+N/l41IS9oNJF8IUhB/HCoN5z3DmPSmdeVptXD/CK7fq90AdqGd4HGcxFX
0lQG14MiSlnTJ+6+ZXVYUdMS0dLX/ULQFw1cgigO4yk96O2UiDqVO7gDAw3zR7dZRDvWFXV218Uw
1NBillWlxyO+BuTjloIln2CTPPK7Ba2zaMdnAa9FEK3L92NVDGV8PYBhDpV5Bl4TsdEL1WJJFqo8
QV4x1Q/eY/1fVQxIAT1XT/4GA7WA29BsTlrzii/9sR5RepugeGnBjCpZD2j8OnHpbUsC6+ST5vFj
3yM62szXxyRmzxjg+Oze1P+f07UlBsF808XaEdj8I47epK6KLPdT3xQjwy3FqZCxwz5GppNqfy9f
4xufzvR3AZb5pcdz3mqsReDPPf6hBiNpt+VWN23LJN86ghJ2OXuaGzKnGmjnZYgh7vVV2FJAq378
+qIZFZ/xAEZlQ75xbNhp8NV7f4sxEaTNc2D4KGPngZYaY0uJ5L5MbhvQvdkg/WwvNCQsijbZGMCr
jLSitCtwTNC7pCjMp7F923go0/AOBzNEOww9LrqIeSGLAF1G1Lf8MnYqGSGSEBPDD0avJoae2Tne
PGWvkiK22FPPZrHf1kK4eCvoI76Pa98UzVkHLaQihaLJ2FGgWHpIutTMQRwezoCciB9QD16aWiLK
2xLNxxuQm3rgd+QdvFEzeGFr2Y131/6AE1M92zwMaIDYzBD4YGtzqjKHEc0OyC6ontvj24Cyho5p
MMx5SGvUAXjNOA3Sv7V8bWr2HzEkV/HkBGQU+GmFIx7CIfsMxkV7gTEoDN1btx5lLJV4WFK7zv70
B/nMxUA1vnrpf8W7bnyuuVf6tWHAWI26svHT8BpHxcnT4gKPFz8U0X9kAXH2kKj68au8fe6daebi
sWATkgUzlL8RJadVUhX0Kw3ez3RdsQqvQweCxwcethPXgQ5BBOSfCeRDLQIgm0EQp0E8yR+RucV/
wtUB6Fg2os2C0Bvsy1RB+d17/E4RmB49/YxozopJ5ManUugKtivCMmmV86KQNqAgfWoZ3bEFv2y8
VZ99BFV2ezfFsHUHJJ4ivMWw59HnbHP/h76jdylms5niM7OlHqYxn/n1ZKqknhoKMmQ4lsTf2qUs
U8vuNzBQJQDgLar62jD4maM6AWHKFFEEIMsxSNJ6kmQnBpezU/xPTdoVHE/z1Y/3Li8ICNIcTRLM
dEUaUYuzJg/5E/PD8Z+i2G6p1BzVexKFaUnjfkk2CbfgOH0YuQxyYHVl8FyH8V1tvh2kzc/wuP+8
MMZd9uto5QldcvcEIMaErYDnJWmd+n/H53/8erns5N28YQi8G8t8tKo7InIVgmrO9iOVR4sWnZ/v
IsRaZzL4NsLFC2dK7QtGLuuqP5CDVzbGkRlnQk5mwz1nuM3emgtin/Y2pXKHO8cRNSraSlYO0pbm
4IN676JhZjmdMMH+OqALTBxfc9Cf8q1xLHTeqxmcT9Y+eTLXp2WnbMh7ueflhgY26tZ1m/FDPRmM
UR0Gbaxk1rdsRG+czAOP0DDCAfVlFoHXPf4EZsLtXLsR8Z3GwZH2Lr1z1JlZwTeG8/3cgbdvMxOX
DuVZ0vLF1+2AfNY7Ua+hSMHLrNfL4FBwy6eBIPyTryTViq7+uqCfqZXGHrhn6hn2+c4p31xZpdE3
OJ12dcpNnwFr/SmpXZXD80c8mHxq1BwNe2k5YCa7Uhn4uhPIiGUeTt7YJUjP4l2XNqV6JSsDJ8Cr
5uz8XVHwKurx0HJoTcIkSH99CsAqE3jVn5g8fIj/vLvX7hWxeCtV6zDkA6KOlLcDLef92Zb7wvly
q1Mp91dVeQNPAP9dFZ04F3eg/dK3tX4RDd5Jw1+hQVnU4hgDk72sD0GuxHXd/N/vSE3bB+5E4E0V
r6LdKxSfZf789Op7kVfXBW4yKE+rejCGrZuqQ5CvD5+ih9Mg18AdDCy39VNQUqD4cGeK8kKFYKEU
hP5Aqa2wnbzmStwckYnsjX+UyXFUbZNlqt6fpUu8746WVcmpZknpdb/CLGxS8d/DFz3SSYxjjgl6
VCDsyFygj0wCZ0iZk1SE8azlaxxzoa6xGFUFDTRzPxekgKciU061mbwsFuqZP8pmqVLYeFjNzgN+
xBOwQf5dG/ICwsQyF+uY1ZrICNr098z0dvgmzbjFV2Bwq+niUr8fjazCWht7R3ohEb3ye3roTRbB
bE1vQcVE52Tc1gvQzR09tAq7hSOxkaT9ck2HYZOmvx6ATf0qSEaphl8dW150JXc+T1eRWEQ2Z3XR
zdOVCG3eQgBCaCIlPIQi9cRPxwb12A66m8nWhWINGM4SyKfINvuY7kVjk6iGerpow4mqk1e/UyiA
HB5nOokkkuNbk65FWFINTn2GMAy2+MLq3xhs8aRloZtkvwJLDHSIih9bBlNHCFokN1BzHvZRc+yn
QwvjcHw+0PL3MtlhxfE9YaMZDEswzotzlsnNbae6cNK2U9hH56T8q2RDjL86Mci/17UooIqxr1vM
uaDY9qtfNaJStq2/LekSNGmDFnqjn5PYFfU1smsMnxA4qC0IZb8V8OnLoouMj6TYsJPdCqnjZP/s
WCzRvMWsVQu0D5NOMSet9oe5LFxah+qgk/m8K63nB5tzqFj7jAxyoiU+MIGavAvXm5BJ6ox6qMAd
ke4Gi100Z/324/t9B/aTlh8anTmtcp/n3vgPOQSIcOCTvjxZwpWJvpqHUJyRAcSwE6GDPATeeudL
hijoqBRI64kzQxcWM1c9NJvwBQ4lb9+YkNawKK+IOXJU+F1AUUVpFSmDqFiQeWIkvfNsghQbKDZX
WzSmBiSda52e+YmyRMXgo7z1+HTkik8pAp48hVYosEIvZ34rK9nLxmQSVhTbZbDEnjIb0iQpeH/x
APr3AMRrENQndzBwJA5rltWwXt2uOvJsfhO3701eszT8Te1vzWrN3vWXlSz38I9mqqx8Ua31RJCL
p+EpAkcAm/NoGC97q4WUI1Uke67qx3geaboMZ978sY9g9HH3eViTyX9qxc4BsoLaNxs7BvV9Sduq
YCapvh0EeMbapygzCtMTagRvNXYFREGLB2ii/C166AMZ8Gs5L7aq5E2epfe0jYIdVRYkEVNE0yf7
qMeTO94HzWRQLsySQTGY43w83KY3kG09ORG9FsrKcKktXUgHTLGz5j7IYnsZyFgizm5QBCW4hbjn
dyyPaB0tsig91TF1ORNfAzawgWod1GjdoUQBMRxkj5HPI8xM6kaT7UUlDIf3lyyxUpw4hgTgnH4V
CbMubs92ixJj4KZgXhlHHbVY1p51InGjNw0RbiyNCQUL7VqLj64fuqg/67D8LjMY5O3/uvwE79db
ossQSUUNJfMbIGWTNFkhhPOFnYUYliqZ0YwYfeWgYF47AIMUHeDqQG9yXU6oAuFjds9ibd91m/9J
73/3XWnSW3KYTEpGOXAEiBLbj28U6r8wW25evHpY1i3MxXfyb41hBSHo99iZL9veLR4i1r+kUNg5
l5SBPQKSaITJLi/0nMjDfR0ugJE+H86+4i8zJttk3sq1GZsTkbj4E1gZkOQIkGFSgb+VHtjYdwI7
S7m7bUVrThSRmQdU/jKBjeRViG9kC7vG6uy1McTplMkYaILy2c0i9tdJ04izYGoc/SZzFWeP6FVM
FiIz4q0DeX4V2qwsTP3kkvxNus21jr56hDOQgP8+setUeTWxfdhLVAuGPDxEU3qFlT7TVV/0A1w2
VMkfacUuTx06g10AiCVh8KcCiXXNNEYrd1xXboYg10PuA17aPXmyxtcFZE1LKjjpTOnxyMCnAlOG
ubzI5eDFRCOwQZx6DFwncCeYsnfZaO/ZsXEP06rbM6pXf1j4pG/tBjIeVdKLmYNArkPXPz3Nq1CK
746577oBtoDFFYSKqnMIvHVKQIoGxLGeiqqrYM47dsx7WfJbWXcIBAoLofxUn0LnkWZRyyML0UGp
kTy27nN0iyBabxK9W5cAKUZbSP330xdIggtkObeQ7xNiygPEwUXtpmOB6ARYpFT7Ln0vvPTPdTnS
ZpQct0a62mqS+R9jXzb41qvybbQnuRh4SFKVfTLR0PKh3rGGmIEmGS8ay3xR6kYCqcyMnhdMZHLK
p727IKpAHAn0LF2HcqhKNX4EGYkukJtVjCl32MQBpT/93T8u9jPXiaJdPyU1DTXm0cyjCiaSS+NP
tmfj7dqy+xXnGC+ocSjVzSPCgF9/tG6I52kiwbP/TyUerWiVTC7jzNe7hN5JSYBTmQebZ2oiQjp/
o9lfz+VkO/CGxqZF2lyr5VLXZB1svX+sXdSjxeV1OLE8JojklLNkg4+DrVtZzw3Lmz3dMgVAFljN
miX6qVtqbeBbAbDpADavPzjvKbRJarB4dppmdXWR9vjZzwF9TVm/mGORBUWyQC4MpTrXaBKRhapq
G739oeJ+plyKIG2M68RIfPTiZgc1VklCOYTp4trOQHv3aI9faHou2RbAUtR+eWWznO9Mam+Phf1Y
g0uUff/3nU34MTZhtXvdbxW4bEIO4XFSwXacbZstVR6YXvHpBX7mTjwqycohGt4t0zL6jnPr9k7J
ZaSoLzBqWUzCLuElYgDyAfh3bq8oLvVOhamQo0ce27isNFToEFIjGQNMSx07QN2p8V313RrTOPe9
zdzYlWnfNHyn7ua+xc/lnU1Ck63CamEPCm1lcQ301AN+7Yef4n5S1WaXTBbtUbTQzuiyhoZ7fP8Y
sUlSqGmg5xFbk0M8TrQ5OLawda/+s+v+f2KgLurH2eYzB9Pu1VHWJrQLx/GyXKD9pzVZpC3feKdg
cddt6kxyAEjTOtWwsVKIVdPduWVGozdt2mcsmArKQJt7vvoRma2kV7UNvtiZ915j95Nhjx6pEa+5
rmKcz38UclfjZ+U7VPEVqkwVO1qlVs7KJiRoW/BehITETwcaa7FR6uo+x7BtXPauYimpw4Omia8N
3NGl+uwaKW8UP9jDb2TlNWM1reA2wv51kZ//osvgxsrJpz4K5nG4TOq8GWkFnfqWhPkOwC2UYNtI
xugT8V0p0AQV0EVcHUJWX/0QrBUI8OzSoPiYn9HIoDA7cMunkmH86M3LTIeHIj9IENezJtMuIcSV
Qeza0wbKOR9IflxfSUGqbKgiQ2ZFrmYtyV7D0NbPMKkILx1A5EXocMr+sAw1ldluKgbxkCadihZ9
BgDISEPW2ZvAqOO0Xc3jx+x/N8ejGjyJp+pZoS9AxFRZBGxBdINLOz6Whyn5Vikij6wz5SIitQrd
uBOPrrmPghkANeNjMhcr+ed0VDg5hXXOdyWH9Wwied8xzYS1B0WuLkeQT2kRAbBbOkUt2TgdC+KW
P4NqXijIC4NM6Axlbg1kIlnMH7GFmVsIrDHm/6Me6IVrpSRTrR4OXmy24+nXzL3s7z5q8K//OdTC
c3JAKu4tdAtUWWkTS9OyaCWZELpFk+zAFmU95YP9hVy3HgVOXAJ+d7BCUNPyWGlef/w+Apqwj685
7mW9sxGLvX54gC6Xqg07r8dDInCzoJJIXKH3azLe6EeI1z4nEZUTjvgRWpd3d7xwTe1MC0bHytoH
20BpKInI3BfKfkJRC47v3tsy85Ji28StOYpI/mDbhVWNet5BYGAtcXDQwb7gyFQYCx4BJ3L2lrUr
7VrkbgwxedcZ08dK/HeSI6v4SmS7vihXGNNyAMtwWNx+fmHF7T9OWHclmowHMIrVe16xz287FBRz
OQjBFcigLpS9HBw4zD0ZSqyfjYUNCl1F+afiTfOCv6ZTwDHqtuWXXyU1lITgfeiyephmAZmcsw0i
POZpJh7uaQiA1p8myjlsVCJBGZ5tyhgfCeizNIA65PrGGq282rGxJ4X5Q7p2Pb6Om3rbtt0QUsWj
V8VJLKv+g4ZcCSqOl/+khayf9jHOx7+/PS6wDiEMhDZtodX0uN2KA7K8MtmospxVnBSFJOQTKIyy
msm60Sp0uSUiJe1fVvda+uXF/lSIayTfauyBOYGEHlHg85o4X7pab8T8jzIkVLiGRu77eHgOfUNj
uL0ewCOvN+0RGx5JpHNEVDI67BnrRQXwhIc4QTywLm4BbYJ873xf/olL6bIdESMDg9JxqZSYyt0X
AYDd9psOWye/rcqdnraHJPs3T01+AyJ7K/J/FENVg5Id1eP9SS8Q8EJehX4FViynqU42IlLtosLl
xsF0JnBBHkpQ9aVKMRZ+s2palAq10bM+P64P6eWfjcKO+Bj893ib/48wttSWcX1szuDNPRUDz9NX
39KZgcNvsq42j6ePeY3DOUo505JCU9R2JCEMiH6mM0OxPC7VW24cRSK1b7ED3a4Knpys12nxsN2J
REjZ9/cNQ15Smn3O/M0GOZFsjpMo+oWmp80SYUSA/Y3N27vIOf85XU69IS8DlJiUTZXQlY+feD+X
A9ejnIovfuK6LajR3hruUBo7+dg3Rd2MEmNo5kszRIx28g6yc99Xy9Dkm+wufhCFR5BqjX3kskOW
i+AF0mFYhQ4tf8RwRFEQ13ykHpxW2Bm7brCFrcrRK+cniEQnGHbyAPNCEj5zpFkzrY0qwwZiUc/G
OgGmCXQn1OpG12xMCMPXta6GiOsSm1kOssdbP+Nvm3x2pWtdXKz/fsWJZTMFU0BD7yIht4DI0hxc
QI2zdQHGXGNidRXUZGVfETzMoLRnuaxLlnhhAgh3chZ6MVxEOnR6jCqvlLJacd8M32A/evjAW5tN
7vB1f5thLNQg7Ho3+FthmL93T49y4OrgEirsoKLHzT/ULCD/M/sB4alXLT8kFPuGMDTAr1Xqx0dI
8DQE6ED7D/rUQQUzSsemFuBZCv/BdnIFPndQspb+ikvF2ZE9mQ79+OkLr3R+XxAnZIRAiCcwCMt5
edsam+ba078Yn7XbTRujD6sds7aLvTe6C6NZfVjUVsfU40N3e40f7ZF8/cpo+txCabjJiEHujO/+
JkpjC8irH2llWR7k+nJRGzU1OSlHZ2HAQ5FibI3A+nwhPbLTmD6KUru1CTM7tAedRh2biP4ODZim
bRJwpAAllvyjtr3aNbKBzy4ya1iFr5+92Sj2rLg+umwWHRkfpmo2mpqn4zKlTv5VY/4vxgE67F2M
Nm8tZvTh/APt7Le3nwGW2gDk5UwK0jnlAEWaxbh4FWIXb5aDNghWyXaGwNge3XUdlxC6MMvBSQJO
jWrN0KCWOIxx+ekspd3bma3zvlV8Kjmq/beBGg/p/MOOoLhPLmoC0xza0ima25ppzrgYmno12h+m
xKJWZpv7GXq0VumKIWJ7ydSRdKCSl9Oe+x8o2IhyUMQWbuRbOIcO8sezGoU40rB5fHWHEx/SF0lD
CHfXD1NMDNZYC5+UyVeRKpf8B3FLqQMyex3M8j5c89U/GpxHaEPKZU93LK9/8IRrzXodDv1w+7n4
GKrvP96wr5HHhj7iycnAZz6lA0De+8wEmmAqdLTSD65g7IlNHsOK7U3LFWdo56R45THTpk7QHdwp
qO//B+DtDNVlZwSFRIJKxzzZowpCSvCP2AGTzOZ5AI1jDLCrxuBXO8wcIIVMWXYcQufgTG20KB88
g0K0uQ0x4m5m6NpQjLrhSNf+JrS9xX0MpRDf6Xa6kgE9z0N05rCQ6KKH1LAKQE5CHFzkdHGUVMMw
tmaa4pArOLfaJX9TSR5lZqKj+J0KqEce1a6CTll6rAmLImV03aIkwsJyWtflo2CcQOb602t5nnbK
Vj0zTQeTrhxdm1Q5gOPxynJHanDVGl5tZYsiEdEfwCVeVAGJUlJjvpNdG/C09UBSJ6ZAuPoBswI9
pf0bdEEbreGylZ6Ozle1M+8dOFe4pUcFERQ3gKm+u12ISVQrCSA12ywVo1QyWqT4Sx0X3hrMA6+o
2wUlJj8tLQvAxmwP9DsFWaztLVd9PfaKWJNmoGhXVPO17S2Egy8zfOVZKOjnlWJMQ4HRoy/ZNG0P
ChVg66pY3Rc+mhX9QFiUBJKHLxrk8VPmdCbA0EMAGnTbjUFPIbpCvZ7LMZE1Fqb8efCtmz7Oek2L
BC7Nk0uwOAX/6eaBdq0ar+N2tKLrnnehhWfH9LTQiocCf0RvTBmooISqzSrk4wTrxbCfjdg8Qga5
qW/3a6EaFHF5/Nqj9kTz8/31bEbKUI/KgAxvN0M/pNdlyBr3tAzsjdkdFzRAzWHFF/pcBEQvXXRi
T7PG3VeBYE/mfCwawPS0vY0dWu4ngVezmg2RF/b+x38Fqf8pjYcTz1x/0adtBz7kHt903EM/vGNa
lKZJYQFDRKDrVhNOcJxAPMYkUbGh6YO4yoZI+dFmQ/Q6flrULrtYJshrKw2xXx5JmanHOORsObSa
uCZwi1/m9BlcuvBk1ehUjsf3Ev60tB2NL+988uAOJQl6CXm2FiL0VjJB9OfbcwiOvNn51Bxh+S4T
ucV4J15MH2nIV/H0OxSik98Atsn3N2CrbadGbSHGmE6gDNhX9MkqIVsNeiC+VA4FHVLlWY79fegh
T1uNL6X0s/AoUi11vfPXkGwvXi+iF16MSuFmR7UzTZ3pRyVh/szOI9baml7aKf7JL16fX1AUPleI
wuAhu951gQWURmhbts9zAoKseC6KxRSqetmnKsDID10h4CxVpq0PdrJQFTaPDW5fIS10Ay4IlEY9
wPedP6Ncm2A9HWWF1wZW/sQViC4vu6238IRyTL2BI21ohsHAkA3vYfGkne4TGJQLOR1MUMFGOuyG
60bA7vY6cn18548pFeEDIdIYq2eG3DwLWekDP16NVOxFJ5luseNq+u7n0QjYKgGEvmghcdlG501W
mp2zrC6rrtFumVLHCDEFhG0b7OTpHitBOieNIwMz06b9yLcCqVsptAK9ZgoNvHiNCAfBeq/yrpVN
W2btzI7F3dcQkd1Zju992OLF9oLVXbcmcrkBWyEkKQNOQX5OSyvUTSdK3hP5TEpdjN+1VMj98pDV
N2/aJq0DL3ez9ThszU6VbU+cgoeYgVaY9ABkwcNRKmBm9f5J+0Iynqk19A9/UZcJvoR802ztLQAz
a2DBt0QKF6ZZGEOd5i2dmV00vXXAbxc2/bxkSsF1vlR8xleh7yvV+fMc8ftqHXclaM+VoJhp3Fsu
InPtwGToSONUY9kuhjPStxEoh5XuDF9xkqQBV7TiPR3wJdl0ZcECHZWnEmo6QaS9jbKX+EOhFJ0H
MYfKW8RJzR46pj1LJWfGRSkRcvIfLvVlBM/Z28idqlPiGaTHPlrSTV6EtoNStLgAQ/JkcOKTdTMM
v5TeBMCz06+BZD2i+450trYVV5i63u2IZTyZDk0ZfU3fX7YqZwNHBxEJHulwuiRoDSw2JpGAlM7g
Qv9+3qLwmJLF8V3Sy4e69CLgmahDIbsIk9ZEOCdb809zCW+JFlsah90S6MQLDY8rDFYBL4AwcfhO
XJgtJIqZQMZiD8wTn2w1dUz6wV0yhCwN6rsidWYMZvX4SbH7v6Mmu6YYSK7nXUWke/mVJafeCuKo
lVXwnbnWumUTy03wM6rD4yRdfAdMRs4CGtwLeKYr61XJGOI7olp3P4GQeeGcjVgFxJ/bbGuv7ta8
Ux3QKLMhfLtu0sPCy5c4+8AB1YKslytSAsK23gv8r0dkwFKxubAFrSOKNkEDwh0yLqj9XF4XAHup
qlzB0J4yOs9DBv+oK8IfBEVEjGUDp0j7zUDBwpKOjsAV3sfFQFrmIgqqxkKvvIP9L16N8pwveduf
VvNL9Jol6WJqsEkmSk93noIWjRlCvN2u6Wiivixw9IjqHAAvUabkmWpdIwMyNGfwxVSnQQUSDbUl
9ATOW9vHIsnIivpG2X9BDOqIWhH1T5KerK/C4tl06O+T0FIhZ4slNvg73jvjMJBBDLLtHGobFA6m
GchpcT8BcGIsXx3BX5L+jajjnYGp4fsh2Ir2Z9oxzF3s4+H4ema4Cx20mxoewmOyqGeympmxgLRg
UJOSv751Bt6pfsLMGTu2Y0aSGJCP0ZiH6iPx+otkjYfhibi58GMif/bCHBJ/L+9ZRvH5+tbkXzUG
yzZw//KFBYvBJHY3ikjCd2P7/AzBbAggoujre0o+d6rFFu0dXZ4nWheIHZJnn/Zuxrhs4nAx0b9W
D3vyASllct/P4rl5JhmtkgsYTkWreckghScqESVN2tLXp3FrNn7i3tjbu8yUH/SaOBfFQ8ZtJxHF
uBXh4qt3o2mBQknRwuh87AlDoYoCw4B5KxOjrloyVbLyIHmoivclWl3BE7Kr9RSi7OsbEbf/jfWI
AKg4assYPBRRyKaOGhW/6xjBodc9jA7rYMiql74y8Zr5R4XK4VMFW0RbjKQcpQRt6zLlomcupxs/
FmihESHwlgYwHG2iRTym1QiUNIa+PrnjeUyB951L96dQ9maLPVmjwf53Pm/YGts3ajb4KaMiTopT
iSjuxs3Z/WyYiB93g4wLnqHlNgrunAQlckTdI8qMo0FBuM3wPWEcs/hCY3AcnZ/mz8o7ePPFJ/Te
pH3DoTji3CagyMPphwc5d3Zax2VAHCMuxpiZp9quexFNSNQM2VTsKIcswlXaB4h7BeSsO8NSHzSV
FIQW1hcLr6QGMeXxog/T7/XWtmq8JLG0DiNfxpFC0x4IAZnmRkBd/nlkzinnB8nMdpIeq/5Wlg8Z
P1p64I3P1iIXCzmLJzZ5CkZWAEfOx3l2AGSjEOroyXotw6phoAW4EHRuLDexSGJ5KV4BlHWx1gi0
9PJndKMOPprJFSukv2nmRnp67V3zDutYM0TvtTZXW2w9icUA/FyKdiAC+LeMaDoLNWuXzmBAVLAN
i43d23eJQglTIk/we7yK9jBC7dBRJwVWGjUsdT/3t7mVJjSEKq1cSjQ3pSu9bpK03pBiJXqe3h8q
v0b3K3yLuFmG2mNSG0en6kTFy0mMAdlF+YC+1lxUdxkrSVsbbKZbT1pEBVL3WnVxv/MGQ9ttrLhd
8KOJtvtVu1481J3nUu4c1R1A2+Lg6BXD0hSR/etcwsiiefYjnbZyPQnhY5YX2WQI/j1GD9SXgcrN
j9CzFIyp2ig+clXmtrbXnVE6jszCDFOZTDfdg3tnydr6Fwlo8UM6FhgN/S0z2vALL0ydG3b+7bV6
mtf/bKT447CvwwTCTaJhQBpRs3BGtNzYP28XOA+nQTZQqCErIC4tkMn7BtfOW6CZZqrH5qd53ZUQ
IyxHNQmZ6nv+wpTIelSEw5wloq4xHCnyrbu/a6DdDDvI3cgqX+6zmU6bgdLhTdwkMGBTiIIX1q7y
w+UqMRR6IMZIrXHbxbzxoqSJ3xc0r+Jw4CCjjAQa3qcQls4TgU+GmFW7sJ0JII9AoRWL/tu6+CzF
vDR5vzVcSHr+OiRpczDNoJKbuMGInqTJ83L3HkFW+nCWR4+JnhtzGOH8Ab84xs7Rit9AEnU/PeNd
jxJjdtIsiMZ3I8fVVkGCal318ezFNKiyTqFTbZhlAFTjL+/pO0+Pgvv28q0vRUYe39DJcS108j2n
uQapbilwWIUn4z2ESoJSgOAZmbaJnki8iIKOCowb58IVzI6J6A+nkN3K23iz69Va33sFdP760XbJ
cwaGIc3Gn7WhuGDxBjvVrO0/PV3JAXhHC6agrQCKkGwTjVsryu5tFbBdsPPzeRmMMzluJsGaKAp9
Nww8JpHZZYHhEsecVHfzxedJjRKcIcLlNbB3zm7ZEodDmFQfACTXkSVNPlbC9NBtCTwtb5htAUQH
l4F03inA+BpzsZBjlSN+UhcQxD3EZ2Fm7+v0UknnOfkJZJaC9ef9djGsJ58Az28pDSiNXh52yj8C
3AWdPiIrIP6Ces4COQqMsEbCSF6Tn8BR7xQKb3iehJNjR+YEaNVhgUKDKM1Oaj5k1gZJ+NOg5HbP
fjdNUTAsb8J3rmWJ/JjgS+4KeBtrTEzLS29Mw5+AQknTdcq+1NBM41kX+IyeVwk09PVYDgvi+16x
WS6zle7BiPLVsjVGO9gvfxC33M1T8QoWDthLoU1OwG6pXxuGMIINsj2j1lB3Vg5HDRIa/1KL4mq8
Im9g/ywmfkW1fJ++Ff41mOpzTZycKUYQxekkMEC4E97uBDWZywl1Vwf607Hx+G1c4XhRd7v3/ToQ
UPgO91qUZP586E1UgVEVOre52E1r/XeSjYh3t9h3fVcfTFSxGjA6mdwabYYLgqx13rKKA+TeJayV
bXl8C2PiL7GHE3nvgqgHqaMvObaxOdETmI0liToL+4JiuNxaDkjZgrR1e2k5fwjuZy5WZ92eZPC0
uhEFxhzxedH0KpKb5jfmoT+G7zzAfOkQbEVUMMpZiKD7wxW7z4U24Bo2VbBzPwQqsedzL7BQSpxD
txRMLTba3XthIXn+o3sfBKicYfQn7i4undYkPttn5GK5AhD08ZDQbGrdLX+1mz6ckJY6qzF9KyHN
JK0hTc/19hViT2Ha29kG4GAq26F/7OdFEoQn7NhokDUXFVJEKNkhDYB8BHCehY2ZsxvenVWSwm2R
XTfLTUW8Le35S2cgi47d4VB/y6apx0Ux6YdXQscfNI9rC5q9CWpdZemuJKRYHYJ7ndrPUQH0LAe1
10IGb6MARWRv/FZ0YuiTplH653RYQB1ZozLrsRR47gTK7i5gbGOy7LPkygb3ZKL/qSgjEvEXJZLE
eC0rbutSlMy3DedkiqAzd7HbHkxbit7CriWvkb1k9vPv0eC523D5WEjVEgsPr/GQq3Us/0zU0aIw
jy8rwND5yaAszCx+pWx5rwQjqveyPNdAIw3hdI6SLHVaBBMXg1YXY1aSeBfpIing0y/XV3TNUOY3
fNoARuCWsaXKw5D154vlZj9LspMN2RtUc7S9G6uSc99VPe68YNW8bJhyTTECY9pJa7bXQ8IJxACX
Tbkyo60CzhRQDQ/KMRHGM21xsU3CwpmqV8QMjOpG9r6hYlsY9srlYm0WLjlqjvNHu2akVyra27jD
1fBQNoxj1TWrxDJRa2aUbizlM9qslt7DznGwv9PbXV4mFL+Q+bwZn3BNree+iNgzgP+CSNjGmnjC
8gspdI58Ppbebfh4cWq8+UGW6uDc9YpZxk9rQ0OHBpXog4H8QAVtFIsAL92PcvxHDHtX8ouF0J/h
HQhPKTlM2B7l2NYtwIpaxc3NrXx8IBteDzWsyhh2DAubn1ia3JTKIdsVed7gofdtyEmrrf37Mah0
NQ5kcej3/VQjrGNxJMM16jOOh8Z0EO1yp2YofsdKIrsqTiaVVGcmkn0HcKmETjmRBj1m4bcoF/UJ
cCM/7cbAnwmHVQW5Dbhuw7euySlRU0SM88v1Xt4yeQbS9jCl+N6T3ThNk8267P3LI5FNCSO/lapa
2UEXZ+zoQyuP/KhVjYwwMELa31xp6fjDZVhE4ZFX6VpFWo4mGxhmw96kO6jtne9WxVA8ll/bR00e
LfijGFgs5Wacm6MekBWB892l8mRZh5tslj/fwV67KxgT7h4qJfGsZa1QyBiVttDfn+pyOO5nJHGN
G+qrZueBq1nDAVV3tV401FU6be3rpsnZX7o5LtA7v5r98+PVYQJUEfk2cOC1Ozl9BCvWA8A2LGga
guwD8YIxHAf//nA3VZlVcaQkn06okqdsBTETHjHRAuYi7NYhoL6K+DBeoRyunAW+Ena9HldVV0gO
0Q5fw0YKKDHkpZD5PsQGGLI4wEolfSFQbh3Q7N3Vz55HXe/Qc8EReygthvSenSYzUOgPUJA7CZkA
uGUZDHl0cHAFa3lP8NBmOHwmT7cIDVHN0Pi+2LC3f4wQMzqR1t3n67dvxmTvPjsKygV25OpjDUUl
WZZ1ijwBu4YT/kIvyn3FUMrZ0+krBeISV5D+Ut/WKzK4+FgBMWWniEEq5bn3Na0wEwgTN76szE/4
bN4OROhBKBjhPEwlCyd0qrjIn6xn3xwff/ven4/7KY+KlF5i8EOzU6WkNgRBLcYyJb8IgQLFt5Wr
Cjy0wYbkjzynkccascCdiCYKIL/TJ8w0SlCOIqh0FapJURuAwSdoG4+k37Y9Mnp+NKkKMzXlcvyh
tpP4qw112xjGMEQEY2n4IW757VRP127KBKG3p0TyxXtMAG2aQlZnA6PAAFysXXBuou5fjGOI+7kA
t8zAww6VU+NDvIzfsLajkte9nuJAc0qslKjeTErX43IF9k+N2kxW/4QEcp30Uthbb9R5njh1cRD6
UhvJiCHtjxc9z06pfLsSMso9viWDN/KmPIj6j8kD2KaNJDNr8DIKH4D37/9F5W4dzjj+XizWpPgL
n4aiFZ40IZus05pPI6FRS53VoOTvHbcGaZswE9KlT1Eo3Kyjnr8R46OQPLs+z4UfWY1vMDTWGbGE
3cL1g5QnvJYkEiZrGFBP+C0t8EzaNiHX/euO82tuttK4+Jk7+yJd0qNNTOQ7x4R1Sq1qFNpezBc2
8dQkZjUY19RMJuFqsOlAyQ7GPp/1FpfSmCWc14NYTV20DJo+s5fxonpsx8khOxgiN9E/dPJgk8kQ
tdJpR0SBskSzWCZVPcy/HYwNBrxUo+HuNvAO/p9SLaGEGLqvGZMDJeIuRz7feEVG0JCTAEU/zO9k
YE8y+IPBnJtrJP8qj1ZxLbspT25suW4rOUuwaA/jMosOayIvj8/1wtyeQ/dO6afICXRbzAYZAr/f
/KV5ioA+VSe0n3bXZEsYNKfmcriVBc88jyIVpM4XqnlqAP4unpnUaq6ym7f/NsgTw/iBhYv8oaum
poexYCfDF2Ef2OW8M2GkHQUQ8hHeKyGx68cWH2KmtWT4Xm/U46pSlBz8XNLK5h+RtdVflTqbCxc2
nuanFSrhRLEkpHeCGG/uG2DYL5d6rAVSpRXNP6u/8bowkRRqGl6ByBW/2nrq8+VQ7GPxriGE21cP
1Sn7rR49r4Irri2fVqKuJd57vpD+Ov+CRVcyrDaVCP1tc3Tw1tfHgXlu/T+tEgTX0rGKgsQj58Bd
jN21osZAz5TMMMGBrVChCmlwFI2KvwGbpna928xnvhHIHgsY9IUW5juEOLiOLcGkRGU7oABtPp5+
KGGJJ36dFCGXdxpoCsDEaA+RRNuHgDvdOjscd3VkG5/sz9NeebMoglG7IiFTm9pWR/BtknIOawOA
OgjGopmb21L2wkvnUUjfndHzOHMuBDfMlzGG3O8Wv3bOSjrgxcgWr8hRmo3MMei+wuTxkICM+KF3
dIQ5DPETDV7xxx4tefr92Goer2wWRhONJV0R7BfrqmeriPUYoEEtcGkoJJX/SlBTf9L1Ko2j9X3J
AiRUnp74EG6o1YkCCYabD1VO1D2F9DIKzeSINHBLiwyf/QxCc555SSj8ofvjpbEw2zcRjtyyNllr
9eBn0+ZMkwaZEcVtal8fs+KiNYO/Q/MNPc8tXXQcmmhUUeP+gQj2qaMG0cBZS6WrZfInvocgwd6f
SOh4oKozWwIrFft2NT6zPY/i+2jiMtA6JNHjj/bw5EBqZjQynp+FUxxROzvmmqd5qHn10hnEk09p
ZHVCqjA4ihzHoBKNsumbwiKmLP/96xXysa+DWKQUoY8Mt6kR2sIbTSZUwCj0s1FiPGp6uqQDEdsZ
WwkJJhbXlpC/4phqkY30XtqsDpIdhLb7O1+Mfg1xmuA1wdChv3Dxl1D/p1WI4a3ge0ZxumaMhYyA
frl6l7Y4f9CKGElY74XSgrj0KF+DwffupYKlWS4kQlVW5vpgtNf0ZkeB1g9k7PLTQJ8ivWVmVNyJ
/5DWDatdihllA3pN41q4t7tnr8sL6IiDV2ydbywWejWlolRncYRtYFiLQ5rXjJQaTs0rK1VhbNtA
V3It1FFPJYw04Sh6UOWwWtgAcbqqDsBTltmbubTv1dd52rKNx5G5US0W6R3LYAi/zxOgm4DD4IoV
G0RpHdfwWSBSC4XI21wlJBs8An7X4c8Mw/lDU5S5hUDzvyWieFUx4oL3ZZPSm+b8XlhrAKtNuswE
d5pxx9hAyfax4OOLf3l6YFjXkYYSj++MHsdWzTCpwIgiOvZboPGA68bwvUxeE22Zz4nfbml1M6Uy
ZFGstPwG0MNgGDnaYSL2teAfahDs+8dKaxxxyt+KfWAMHW9s1r+zeIFMZWVrpw6p/a+PwC2I4cZR
GUX1yHgqeLsfPSP5N78FmMI4cCQB5ObFFGzFqtfDZyNAeuYgCudVI4Cc7zDcvsLzfEQt2lMhrOS+
0qZuoLjqdf7Px0deQK+QZbF/asfSpyyIpRbNwH/0CQORn0vSQXGJW8DDz3YF0SpVtW7rYQ+T2Chi
u6I+GuuUuJj5ioJ3bvy82LNcUrXYE5VumVACTUjkCn6cC80GJ5fvCUZyX4zGiY3fStkWvYOP+B7P
Ps5PFKOhUu3uSPewMZn3pZM2M6nErxNf5e4Em93dZwErZ3jBO0P9R6pzMSsC7OJasm0BpTQy82VF
QtqMoY3MvAwRPZ/h79t+gFbL9+BOwZ94QX4+rcxNi3PjLfODEQEsFnnFJxOc2WVI406kHjgkFt7b
FGbP03mp+CRjCz3hySmAvGg/5spEknWzN54/5EI1C2U2MWpuQQ8mvBPIArmtbPtcsNFgh4Cc9CdT
FgQH/KA4gkcRukWsMJHXXFZBdtZ56xuLFlGLebeLEeoW2JS25Yj6/1xJ94ztkfIrK951F+RaWJ0G
F/hk7tXsLdq+eKOz8tLnMTLxvUtdeG53AOCpT6Uv9kk6vDP9wQgjW67dXNp/touK5yl/pM6+i9A6
ov3uXAJCy3E3CjhxBXpQiS+Ls4AxXzCS6xZEEVVqtGHc2WCSa98IK5e0mZSizrs5x6jxWZ8/+bif
ii+WOocVYnOZKJfUTIDvsqEr9I6GEvaEOd/14kfJj0mMIhxnBIrvY3tu4Croz8yUZ4Be3CMqmOrl
RX1oFnopZ40Otz+4pvlPfQ0EaMeYrtyJI3qpJP9JF2fmLU3JgkFxTn25ofJf9e/a9E4+nfHQ50tR
7KNgBAWlsk1rDTfcvEhQWmWfycRpth4gNVhYlxjTRQO2812EW6xMN2n1NmaGJNfJRjq0bBe+vQe6
jGUKWhY4htb/kj0r0+F/FDN2mE8yEKHZzgjkfbCyMrnUZ7n4/ySvZ9HE5UpKqVMcRsuEMJlV7EzM
nSt0h/RsDhpLqEhZl356qu2vWfPr/kXEmG7wV2/B8W02JR20RsS4/uVZs87h1+6qFFUSW3iGVYFt
knNdEDOBrtoFLbDXRiLt5aMJ4Etgdn13JLM7ni2iNgnXNOiS6LOGa5UXHidE6mrp3pqkX5xrE6ov
/rgSgbXSzedth+ptEdquY91ifjwrrQ4PKt6uEBZT4u9biieZgVpNQfKkS+XR9N03YLxd2tBDExKP
1Whfn/n/+jdRQobJBzO0FoNXREcm0th+KMuceQeILRoZxEe6KsPk8BejEDsvoJ4bl+G3bDKiSl6p
DCe6ahwvvVG2x999nm87dToOxWjL8T3tN4sBcbQasNzSaOc2AouSCHDVPlBd7jZg361tOSRuoTxw
I37qXhe7nzDlG39QO89sV6X34hrYgkN3mdafOKXNnjSCaO9LF4GjEEXfadx0VYKOBcLJHJsXnMc/
4Irjbxb3jgp20LNFkGJ47zdVnUK5BcheuWSj0yY27nhXRjZF+/MSmHWg92JDKJOhxnnFPq+cKSI+
gxOuyp4HQL0Ruj2FvYDgISRmOqA0Tww18i5i8uUkwL3DVlRTeTCAGoTmY1XDizGhy9LBHqm+10+/
LZcloRWjFKaPd0LGzg3vXNJ/xkKRljQWeddtRD4Im/tvbMpINDdcSQg2pQJ70SnthSwafM1yl0Bi
bwsgHXe2gczzIyomSf6X+SCC1b2GvpFVhmLS7sn6sFNQP595E+DClb3mEepmrNOXx90qAecqXSW7
iymsSinFwGoCVviRi/nbBE3XeaCtsPrf6hBpck08Ogg0n4OrhSfrw14oJGYkQYAwoG4XOY782OfA
ThVRp7zlSieLF0ccE00eDpzrn1TCtA5Z5FDy/6fprJlEykv6IQrbvEtZUvgeRmTpBVb3KbTnm347
d7+PYzeTL6MPY5lsrnksbL96PlbTQwVShntMSUBUPS/v2m1bgwEzOJIFjiNzv46nM9OcZY0nCf3G
3IXJgSDg8GKIM8BXeqET0kdXsLs8PATsQV8dMZqVjUTnhQtwZXIauvVoGzJ63RbdEirI86CZX6Af
rF0eGmG4FKROnQiE2duOiwIQrikq/w8xZ8qu2ulQ/ZTkL3azDnkuceKeDdAs0D0ZNBQT/wI6aT/H
7s+wCwf198NBklAPzE44kHHSPCrNE8O5MmtY/hEYcov+YvcPB8aTv94Y0vLgfJh4DXw1m6BvxeTy
6sXjEo7XG6LR4Ie+e2i2km0PyusmMjYODb+eHbezFYycU62rOh5nMFz/UYbG2/opkm1paHqVmCBi
3paaReA4jSfzOC+onF14QaHhOEV1heIitdEqJZTyLl2jshmVY6sjjRznWw8GBV6v/d5ymBGQ85kk
vjtAfuH/cRjN1lsjnpQV7M7hxRUeaJICOrSAhzyP9r9A4fdkBGpqrH61VOlHXuhGS5HBL5ummNun
YPoIv0W+Ygmqy54SL00CYIlrABqHX5xkry4XaORG3R3Nw16MbtfBLDCIluHYAvOlY7qoFoA5mluc
3XPETzeDmGf4gSeTKmEK0Pe71OSNRdI/68suIHGa4vmSh7GK86B2ngDuS+6aJERb5Os1G4dUdjrT
JhWrZnEejMeUlm75c5LPLx1ES/5JVps7mkngoU6Ha5BuDuZqqwMsMKBEOavWCHEVXF1RIvq8CjwC
MZMrH/KbxlQuIwirDVlnkK6sZJqTAtwsMR3pzBP+w87KCdRGgqjWemSTOCsrYKM6+PmuabjcqYn4
p/N8XK++CnB4SRc4X7mUiPFQpzE+LC1a9HLVRpDsZoYGnClzEzKbHcQqNwksrHcj1FoanYuE2a+a
eQvf14vtPc4rce7SddbGL3L3N6BNPqzsjv4NFOQP2UK3gVHdYEBkXiUvzokUD6h6XJVyg9IzeAnF
QYb8dPMxJzj1wLz8TEj3yaaZFH91nC5BJbwIX7SAE1z2crBiHdYR9wWEF1R9L5+5/5qmRfVaTJhs
WFbxn5iDKPc+sLbYgGBcnb+6cz16iS/f9aaiwxqyP00X4ilTdCpzfNBhAjpXF3YI4M7K0vTKML3p
mbMg1n89nnUSCa0Ne40sKGDzgG3UrDWMS7U907b5PkHGFpmFg2dOGF4zSt8lTzFG6sD0ZrGL+a1W
rYKqnIMmODWsBn75ELD5GDLc6BOT/BGvDfGEaf4WLIcMbd6EWrGA36b54EDHC167WwnKJLpO+2r8
FowagxlcDecUVXdOOdU/MCZMjzHloy5hB9rcVDvWygGqKfKmtUluas1maIh7Yk5SeP3aMGtP7VEX
Ly3sK0CDUNyZZ2OFeMXoo/pgJZIBxQq0Iz9olZOpX6odDIXaxH4KlBhp6F0S1jNDs+CuLMiMxnxz
tKN+DQIthNwfr9eN5HIbO1xoesYDs3jsYtJ8tds7hGuQnI4CMeqdCfHR5BFA1AqK3ZF3YkIT7itT
nLXmQFKS4mGjujwOUOnZmkcj5lMzbNn1neu6yROK8LPsSlAikCUnc4MYm42KY/d7sdQ65vhOyKZ4
K1xsAtJkYPs8HtLp7a9pdmkHkg7X1+trhq3N7nCyylYAxidWAlg/84HMke2gK0IdhPRSfe+u81/T
oo6HlRucxFMToryotzIdoW1jCKUwAXcCUeT+miTgL8objbIu4A+SMoAKkVxeOU+l+BIhNwqtx0mn
Y2lwkHfg+26xceVw1xS6zktTLPxILaUwOmhb2/Bk7BuugHyygh1TVZZTp+MHBnHB9G4v6LzjqJPw
VNCkOG7I1zjtcsPAP7FZMfZmry90ktgEj1pv2uS/v1K0jQ6DTQOSXS4Rmz6RSwZm9NR06YsiURE1
F6/VA/OYzAPmCO/BpqVd40OfRAoG5vgboWx5mkfLZD/5D/UYUxqWuIkY5lkFW8C4yN1Tt3+NrBEx
WORBEvGfqKYJ55tnj+HApuwi1WuUMgG/XQ3hghrCaORoiPp8oC330upJ0uK44WZEKz43j4KKgkWt
eS4vBi2fhdJ4wf72h1dLGezz+VRivydt3tOw7gJKho+RzuR8inXa7sfXq0MZWA2YB1he3pk3yaB/
f3XFuZvdnnwrhiemxC9aguseMIw/ew+IBAgRq64glR9xi9syFrHzaEcU+eb7Me+J/JAB/IuU7bMH
TxscUcb408yVv00HNSKg3qMxjPZkE8ej5dfIuc9Z9bzuJkVp4NzABmdRID0Yf8FphwLL22per3a5
SdhBLTVQ/Ly3bPaJO5wyX0MeE/rqXeC6WzAwQI18Ig2TDJvKolZ6vrKtFXLRbo1F6A1jwjaxV1Fc
LcN1d5BNnwAWDEnMkMZavEnTSzuOqVjXEuD94EAN45cBZ8nM03WSJVp7PgPWMAMmdh9OgZiQqfIk
pQyKynPjiRmev/+oOUfxYRJr4WYLeKFQaY6m/hNkRzVmjEMDUljgPe6X995imz5YJNtdtdTsdTh6
Z5pxu2Ar3EP1trsLDiMqCpAZY/EVWYafWSrpjMP1dFXk+KDamSsOTNhglSIrkuVf6TPByL7cIKiN
7J4eT/wnNBpTCDZp7Yq2ala7xOu4o6LRTAzN5cekwjmnHEd9bYmuf0YXDM525J9UyrmIp54nKhcR
rZAeZKvWmLCvD70xbRE2R7fUkjKyGoZuRvittTm8iAMlxLq8WdONE6b214thCXVO+++Jh5moOwZF
njMx3KEhHCmwDs7VJt4V7eVa9cz6KeQUTVUhmJZD9LftfwFqXlQEroEndn/uAcMSkmZpU2N9mM1L
DPA2r0Yr/WkxUoSSowXneifvK3Qkoe0FdT+ObqHZcVg181FfRrlDgn3CE0F++n8Px8W+hoNZFu2m
E9iLiJ2i0RCGXOpYCal8mtLq3pdNl9TE+3ZoE/tk7U03VQkDqAo3sqwbyH6FcSQLNHrqKqGIrIjH
0GbTbFKprFiq1KPYSO1hTWLhrAvmEzeH+eLUjY2+F++/3XhwCgQ27kE22d/LYkMuiHPyl6o4aeI0
2zXLT27yfZyh+rn8vr77rtTJl0yKItRZQr+iKV5AjPr7dOE/ZfHL7J5R+ri5S+7IppxgwjZ31QuX
JOTnZemJ+wvVx3ljZHIsEg2C8fqPuXU42cZbwuH6JkqcFvoxb+u01/8M0N7UsvTIBLgVOHo+iIO4
UvIpki5VE8Zw4ipDeaLY6oRutpLZLoH+X5J7MBEW0eYQiIDlrUGKL6Fd1YWjrJb0W3ZYIMSkY3zW
oekBTiGLxB1C19nDztgLcAbmLT15ITTTJx8H0uf3WTnTCPngO0sHGf0YcRm8hpQY/GKPRyeEvbNo
ADaWCXIwXNb1H85k/ICP6KPgGxZs7YzvIxTkmV8JrW1YMzfUPahN/oBIU/rRgsm8ubO0XN4yVWC4
BJ6PCb5+kR3VJDCuhFDmjmhCOUnOTyjwaaivD8iYGhXqu1SEQkDNSFawUNs9RZPAnzWZpr5pJcnU
urZbTmGvqnVFyROdrykROq6qKfYKZ54T4s/RJXAKY/+TOg/YeFfVcv8u+xsK5ihEqo8FsXev89WW
fz70hQa92ujhs0xWSTIT1fP9RM+cUNBzfy5AWSpb2AYa9mwxVruyXLjgA7+E0fDT5wzyCGHDN0aI
8xxc3ZXuoFfsYWUHwPRUV6zpfyJ/hS7SbzkcbCSvMXmd7etqanrIp7VQZoCn8fn+MYshT51w6qZI
Qu7v85PuMCkpS1nLOwJ275KLepwqK+2d10v9bJ9p6+rlwmXo+WnTHMEjYONQI5J52Q6EMQzzgorV
0DeWr26WvF8f5a+8x4r6As9jss9rSiE6wmPsgT3D9w/QoqaiYf7QyxvRF77etT92La1uW8VxqPJR
eneTN9q4aRX8CRNw+ydWdVV6YmcoYHWfjG79T63z3MTsccB/cHA1oZROdDsQ1gxqSTVl/ax5UhVe
ob6WuXJ2GvcJmo7gSvgyys9inee5a5lJUT3VvoRVV8wY7x/8kWuE/mhpW5jtZT6dE9eYFgkTB1bE
27CG4HFWV/8jEMMEz+Xq9PL7HeKV+hrI+0bQAbXXKv9EgZsbO1A+NujD7yVjhXqUTfhXI4djw5xg
I6+QPce6ZPvsy77b6/W0OaHKVdCPejuvS4LjO7DKRlEcnzFctkBV/iLzYohU1/NSlH+38kabgd4p
TSV8dcQnT6xMfmV8qL9ywLuajyGnF1B+JPmQ9B6xnC8WAnDO5BSq9lRgec6bHJwngEV6BDMHGXGs
LgQ06XPCe4e7syZISl1meEnxvuzTWCoFKNqKbDP1NlNp8IYIHiVIfhhmbrmHgRmsuhpFnSHWgrQU
rcq5geMp5KwERPcYrpG1JeE2xZEMtVCMXA7IhIDaUfJ9oHutLMlR5k4XVqigE4RoCrgat5CRuZZG
3dPEbgWPVJ2lTUONvzjdFFNuzbzKduYQDu4SzupPYwA5flHbQyRUX7Ts4QblT1zELKm8SSBXgKkz
xMSYpFsmZOPVLQv+ic8/qE++1WTVVe9Kcpe94zTwe4yheDogD169nY0XfpWJqmQT6ViHN3sIUDm7
vQpUisp8WBxaCvFMbZsDsyBINXW468c9c+vMB2jvBKltS4KMfo8TGsdF+n6LG9GaDn6e792jjzlF
1IvMzs5fcl7MKTVO36RXLd/dUp5EFYjYGq+nEbJg2btE6I74fE8qv6Rz2FTGBwIqKU150eSICzN5
O8MGtWg2j/FvMZ057m3X6P5e8MKXCENWbyPh13QEx4mbueVdDp8s65bCWdhMzj40eYmG7QNaS1BL
BmtaJQWDmyDRRb+DulNW9MZtv4hOMp+wkwKIDO3lFa4pmb2Cwt7X6CNeZRZfx7VACkt7vkp/ooHZ
rY1rW9iAdMkJrmo7hDLjdTwYUqbX0KDy9PnR6y+lQ0UJI7vlDrUsNv5RgQa6oL8Ce/lLc8DB3ccy
e+XxJFP2OkWXbI+qdZYs5AVKOZGOxqPf06edAn+HNacshKcdqdS9Zgq5KB3X7tVqluul0PHMDoil
YgXdO3q6k8OC6ewKuqBwrES4e2qvh8zaDoV6k2win4C+vMfR5qp8rtTwurB+F9cEO76MH+m7hihQ
7gd0sTU261LUjo12slIlEiLr5idB8DBbZQThQf1NVlHr5PoQON2+xRd45N5Vu4XoAeGRP82EFjoB
I1xu0JCh5vByvhySBhFzdD9zXbHm5qCscBg5xG02qKcEfDEwLw+YSfZLYYAOuj7rOikgZTtI+u86
t0ULnsTcj7AZ3Mx87UbVX364bWLSTimIrVmpkUSAR2xT4f7LuBcsF1acxNUxtoB3CyJJMASru3Cl
cT99AxGNi1ReLy8L2KXannEXYBuwVV9saOnHW6aHTQ/ZZX/RazSTVEu/b5fu1Ep3qi5OyQgk7bM6
XfyzlcsErBf5xzW0/B+jMin1y/YEQcKMPSF0Z/oZEs0U0BssNHiRNLE0x9I0wwTW9Um8Ps3QTlz3
K+8J3NwalRletQbSOurOwFiX7y92I0dgKgz3kcqCWXLJTxpg6vlAH4bU58Sxm6H7AXdxMj2fIRew
J8j3lpnckzOIRARWm1gyEDgzXurhm5pB1P3PuVIq8WM7xKyvnURri9O84s/lON5j0pTRrH60cnau
5MvG1R49ZZlV7fLdDslxgysiDfJq9wnFq4h8T/FvpW9ZRcvdm7trYcydXsrq1AJolqPKwOHxnCee
TJwG9DB2RcZJPeQJbqi5l8pIHkZzotfTXthSdQ8XnuVrM7HVe8hnM7yxVNjwCwKgrrWyD036CVDf
pibVs02QR6uF1KQlwChVNjX7d4S9fgdnmZhnBeND4T3/FHP5oApS/3MkXHPrgdVu7I3YhwFjQGEZ
0XnJpG+U+Bu4qeN+sxdhPSkJoTjsQjYmUSjguRVPWFzuf7smD4feB30nGD/OaQi4Q2S14g+y+m/Y
MhnpI1hBVQW6Q4BRlYEhEqMa6Ve8d8xKrtaYELmbGsyfubJAQlUUJN2hiG58tGtewPBbqKdrwVjz
wWYBBHRBbSi8/Suak8QaT2mJ5Sl1eJU59dI0WzJ77BhMvSdC72tQON6CR5ngtHy6k7CqN1v1J4v0
ocLcaSvt+El7OgcwQXOnNud2Av0pk9wICrHzknydAUcP8EIqr46XkMibp1EQL2bg8TLAZvqM+8RZ
rTIBr15QsgHnJS4vwUOfS5OHFj39PwnrlDxmxlOrNXdU+8Ca8MSuEAQAZk6CZXjxKPSQX3jrkb+n
jRQabNECezHodIVkdX1+JbMsw8LcfdSyH4RaNdznTnpBZZuChRn5JrlfUN+V9D7Ir5cPNdPW9Eno
NxiWTALuDtQVnNJPxwixVkvrLEMr3YOX/ZXwZD6cASJrB9qzba3saVngZW4C9s4z1FWn9QaLjcW3
CbajliFxSmvlYvE4nDX42F95TyF6k32oNziJhJzolX+Kr2wT4D65hbqWRIv0ggXvlWDEcDZMj0Jz
8wf3uUFcUHw6tLlwvgmd6JhiBFTi37i1CYyNeNiPfwuTojr/yshOeu87hHajXovcKkRCr3WWn16q
NDWKWIH0BquySkpXS04xbtw9G7p0VyAXvYY/t8YsZZIppXjAIuvcotfTZ8S12DXVOEs8xlhVYoKp
rGZjTT9qR7buRO/QLvu5S8YDXHy3D4PK5Pw8OB8J8JfSIsegaZztrTvtiVXK7aW5tSXdqiH8u03i
85EUJM+Mj/0nOdb+qNVfcROCg6lK06RJGvoxL/udLurleT9jAdBDuwgzJKGLTz+hFsgVZ/ZOKFz7
kHqCH8ZW2ZOHil1MZVnioNRMt+ImkHaquyd7M73KbVWvCw3E9YAXwxr7WUcJ9rfgUZ/tCoznPjzO
QeSfto8wO4MNieS9fjjvKyZFKGVyQqioa5QQQSmhulKTrFaaIYv+3PuGhrJ/PQFdLZmr1MYZ0jyB
c+PONW00nKwbrfuniNUyfXBCvbsvji/exRTRonMi6t1olYuGjZRKjBmAjhs2F/MT92yj9FJmjllI
MsQQx5NkQR3CYfVOAMgFPC0lZ4pCS38KGnLLXWRR5htAWN3vfRBsWpEZydo2BLVlsczqIpzdgM6F
gCroo6+pTh9+BV5XrF5gi5dDWRMxhl+Gdxn/jLOnKH4gVvke1whd14R6hBPui2jVrlBpxnfVXoHi
2fRnh5HznbBjxO+ko5bT6FwbxLqmGbNVmZUzRWijwkxzZZuhNpNy32ujI2xNUGd+2thMIC26BHx0
BaT+aXoufVkJSeXAYOzT7DellBklUvsjyOf1hTZbkJIN97zaG/G5aH3EA2SzxOYGRxQ9Ik8uxo+Q
3dNmFx5V7riHhKWmgkDwtJqAo8Mr1XpkcHvmisQJ8DjSliQGplllbqMKNCOKv14IuHY/b3dP2YWp
uszHkyT/DQloRLWfcPVYGv0Jyht4yNkJyn6t/9EJF+ncAifkR3m2csxU0T3oSBeSHUDnSji8GDjG
555iEKatxgoqtxY9vcKbAs0uo113Iu4axea2XaD+i+EbDrPt5TjXmsAn6CwtGgU4vlh8E56cdU/k
N5AB7CIaDCtORF+qQo6YWErN69g/jyGVaC2pMQjgwfVAb8h62Qq1yvLSZsdtDoWBjnQPNigYcLJR
hvBzf4kfDfyfr3MvkYMKajt/IjzYg49rQM9AoLHPZRJd6YUPdNXV3N1zZEfOLkw5uusOMlBQ1fol
RVJWOHqXyRNESGTFdA2mmYggBqP6fSxgUIk6XQbw6RFd8fd2o4OSow7L/4DHDoak8NhQSikUXWMJ
URMvQYj6Mf+9DkhlvFOwT8WmClhnMwfGULsDjUrB/WMwk4vGE8I0DLadrmpkDN0FncMaEzKfk3gc
bHog7m4xZxjSVCrY33ZI+REkU3ajTxbyd/6gXaecgmSarpgISamlgB5HV63N9yHgnnHeAUBrxYOE
H1+AmBB3IIxxtbQ8wY2qfv3dK0iFzmJYVY5byP5lvY3CHUpyiVssJ4p+j0axjLyNgWjK5K/xbxvV
yL5sx03LKX9cRvjd/Ro3YyRaYJ529Y6a3+zUfzXL+h911BLwhfXsWsS6xJetLrDTpSKoZahEZ5Bh
r9TBzt/EV4TxMjBpj899lGrVd2WNeiTBLlnudOgHKzDQafRFvBY6FR5i67j/e2/j0AZ7FoQpPw3P
FRa+W69qQy8ddZWEJBR0iFkueDUsUQLCsX0H+eMF9Gf7wIMq7y+uPW80Kz1IDW0bUB5L2/dz3WnO
mFDZOLUZlYjIEqgP8qg8RxhMQtM9kVgNbyjx64nnM0d6opt2BHO8mBrP5BX8yCTde2qwm51gvdCf
GIOWB7YdpDGtJGD8RSheWIldyUoELaKsCkYCmQ4COp9dKl/UAnF6mxa0xo0DRz4cH+cOBgIkzntQ
uZYmZalrFiBWyVGAa432MO2cRy37t2b6wMp02fXPpOw+VeRG/5cvWdwH71MyyxW/b3CvyRpPPZwn
eQsZK1Vu7YvAdXQX3GrArkJ7l9EgfZHych5+nVteRmviciwztZmkiQ4ZQuB/HMQeHpMSL/QduN6q
b1ZmUIphSFsN5yL2USooQeMgmL+qACezG0z935MZvIlr+Onyt/IblBALuemVTGENbVMvMhj0xEZx
oJZO+jKz3s1JATySn1+czvudkXO5c5lNMKw0OnApL9K/9j3o1mKFLC89IfK7bNBTho5rZMBqfBsn
xRxGvwJvDnvIW3tpy7ec7nbT6WNRzgxcAStT3dVs/xS+CXBAO982tPmY8vyZ8APNZTaerjVMExfT
2moU8HeM2N5zennlOGyXMW+48A29vWMHkjcCwjij+fcGh78SPKkRKljZBQ3cdUvbj5kS+C5auF/A
5YIeS/uEt6uqMjB3++Xery2fxEIeWqNHEqTCRehmWX89hEQ55NHo3oeOjQB9tDlyHHp7Qn0nadj+
adYwfxQPaKoXPsXRoN+SV42VZKA8+J2oZnAF6fvK1E0OV578+upF90AmuQ9i7nLlUlloKW5CBjuH
fLuWjppmikLjZjKmRl3cTQNfEGH6uS/JCH0a8uzjjJfTrVQfxaT4bv+DMgmgaLBlclQgdZuSDObH
rMy8KLJ7eWl/0mLmuvUdH9x7K0/oH5x/Lbde4HTtEHuMc9DagzWqjrBcEkfRIF8MxpGjJw3B6nOM
9dKFXFFsx2NVBde/eGQy7wOzlsjGMEqhWHVr9d+c05CJYeSFO64Kr9Mq2pNkz1DAOdIL5ubtNy+O
Qacm8uI2IeugagoOCq1QBKYGGEJdmjDTG9IbHl7ini09MNFdZmrdvmkb4erFkxiQ82UaUC4yA7QX
QzSIGUQNkccVQj3cS/HGA3nKFtuoZDO5Cv/2+mHR6tKIc2DkRVUUADm/o0JkLFNGl/gFws2DXcdl
7EHy2w24BYOFtNv13VqnieMBx05LGs56gHAn5Zd0U0sWKuLXAkCR1ENBgo+98hQatg4i4jcXILJ4
ZGA9PvDT7WkWlwGUzI8/yfRxSFtw8ZkJYp76mmBsZy9ZfpVvf1fdobkkEoY+yVOVxIdzsJPB9iAE
R9FyyvOWxf04fPeb5Z6VUQVzEWQwcHFj4xZM/iOPndpssmytUx9LaMsmeFfjiQCswprCDLTaPUkw
VmuMMN343lrPTfheUgU0d8EUpxi7zv6n0Z1KRX1vISEf99tz6Av0mSW/2//TjD5EbjKIUVAmGHIj
s6e4lHbnehynbQozGj/RVPOacvmdJ2J5gPefG6eK/D96i981SI1hPrJcvcmiyvTvQRij4eU4sCxV
if9XOvis5+3mQVSCd+PSgEHP5TaKoRel2KQ6f3jDmi1b48EM9BmtqfLK57unhub9yA5ngMsWssmB
eAL9xvfI0duwwrZiHdHY3c/iaBj2Ii0i8nwf87q8/WBPGWu5llEgFO+OWi/L5EcrG9tx9L4JBM2Q
DsM9f8VSYShmMjBcFq8OOXjsrDK3dq0j1iu/JNOzSXt+d/utJHmmM8HMgrNhHgorKXVsANUfMUzZ
SnTEYRoFiV+lf99xXsR47Xg5AHRdJjKftmCNZsVs4NfXs4YH+fP+JO2KIrc69jnK5K8v82a8KPlO
OfeYtmMcqe0zrWTKbeQ1OXeX7xpEcmEYyB+/djRzoonS9s6+0+uT+J4E3ZT+tiXCkXsGI2gk7WRi
Mcl7oyYt3HPSdM4awfo/7sbhhwi8GUhwKghvcM0SWAv3HQEOB1U9Dn0hne1wazWhm092FOW9UtaU
jYnG3+pQHrkrXUWSfx57G0+5/0jF6eiHgc4fytLR5jP56Hwa45kPonXg5diUn9rcOnz195+9gOgT
+55opDrigW0MQxBdcePp473K3SIg3IFh9j2aatLXjluYuL+m3naqVhD0IqfdVwRv+GOe1oR5Epxz
gZF+gyRqXaojKtCrERaM3e3U7uVyl1LM52U6FIejnnQMyO0S3jTWwN6c+kDRbfciuL+G8ibl2apo
5dD0CbrmgxArrzbDODY/CzKfuX9N1sp5YejAUH8W9+MdYFBkcjoYFIkz/oOnY917sKCXuH+r30ml
Mbc/QRXHhntwslQSi8cquYgoBoiY85QjQ7JK0MLqZl4S04IyBQR0/gL7ztF8N7F2/P6pfyDYsm2I
lzswOeQLUPADhxTtc4D76vTEUCIjqBmohzkJYcE9/I/HqKXiBmNXQaImjvKBmftsq02oYZh9vkZ3
ETkUNgkQzTsTscqgCgL2vP+IsxBprHGGb6plObfpJVS76XSTdoCtFaqBZ0LWCV+ZRfz/qhVhxXyu
8SB0K3u0bJbhhTbU+h35bBnSUr7uPK+yKgrniurtlapifBjqt7craxDvVJPBbny52l6I/QgTHKKx
s8l0228Ndm2upXha1H3S5muo4WxNmU5fjnb2OdDNmk3fJ0Sb6CxWgT218BlQ5trlMPm2gKuTpIKy
MIbouKZLHAhqL6qh3R1kaJ6yWU+1u4jnqgZzGRsjJrwngut4/dEa5A2kFyaswOMmPA9+AfnLXwsc
u9q1Wo3kfi0vtmAO1/LhzM7WbK4XtHxit3r8z4Z43N5UqH0eVaFRpJxSgwSCcIP+KK29KC+xmyak
CaIZ/xKABvDwpTggr5xL43fwwA4emP47+JaC5u9UL5qdoh1oCLM/HGmSIRBNbfD86QPIEh029Nsu
ib3KamBEJHhXqUD/dVDXSidd15hYq6ksZseWHl91AyuJ57np21pGFmiGp+53rF+oMxsDi65Y/TrW
tqeJfDYtC5+RtKwF3yqGx5C7AB/MI7gDy4ZMC7cGhepKpFtQKqYM5Wz7rQUZf7Z1DMN0aU9yzOVm
bpLlz3decuBPC72rksMkwRkJpIeZup5jPlNMu1GDV9/hCn3+7vJRLyjsYfcfpO/67Xcj+fELHSoZ
4B12m6EF6dMSYPAl8GADKHAuKvqNjQ2ghZ8Sn+J9Nzk55I6K+J1VyrG8akJx7kaiEymDJubzV9kK
FSH43PJUaCqUbxjl9ZnqCK1pSAHsH88ZvLdqPdtYUZkd4IRHBl2FbVdiljQGlIzobk32WueZ6p89
8fjytoeBrOuukqoVAhXACYU3jEDmhbEYB3/++epeXjyDG16GRInmICD2Aoz2QwpVoO6eQaMfIJiy
w7sjhuEuwcEXvqcomnEtKbBVFzyW6pmi5UsJYRCKLmrS45KvUI/kotbTt7YgSqv7SVcnexH5Cfut
Xdbg6ZhgNbip4WsGaZmRFCzWEd/+1l0tTjME8jd/e5GI9leMxoj4XENOzQWC4K/7DBSfifcphgGs
1dZPOKzxL8l5UI7GqKgtbYn3JNlrmOX2qlhPhsWl+q6V9XgAmh8wFqGVOQk/A3zrv9zg3Sm+9PIs
rFLFe6c8j7gGeIgOL9nN8IzrrX82ysakdnpzVML2r0kO7ep/oRkUJWBDYmDrY6OS0eJ2JP4xfaVH
3cXXvFtoAtNSpZlY1ZzdsyOVJKrLP4Tr8tLoDyu/fZFKBdQhJgFhEQJcubk/dSb6hatyNyUxNZPD
oyCmTRDub/88e/WF1to5Vs+BvkSuPXYzdQv/zzriT3neTDPb1cKtN/IwxwI5ULDziL5MaFaERo42
LLNyyGo7Hld7UWIDAj/r5jyfMws/Qfo70SiRn3zr7i7pAe2p5o4RiiQ2t3z3CQJOhktT7qIiAewb
s1ngo4qoR9MHVIiBeMZyRlfUuNgyuFD4lj2LUePqvFV6UukaMEXHl94xyV4l1rB2dyHavJ76OON5
3QP/rmMnScPZ2YM/7CeEWZJKEUvHVGK1jKNFMKUmrIcX5w8O5QnPNY8QIRobacD0iA8bgwgXW6Xx
bzPtm3ZwYzaGcPMe9xDmq1plpnhck2DENQhOiw5MpuUGHizlorSamd2+ywZn/P5AHbqQdwbnlmLW
5fFQdqKl/3q+XvE5EYo/oqEGW4ICcLYSZSy6smjmubp5D7AN3ChotNFOSUhht7xk6BcR7PvvJH8J
/BnrBK3S4f6GGbDhku7goToQv0R2kCVXHzVbzrvHbwt+3W39K5ysg22Hel9u+ulJuwAkDzABTGuC
VfBI7DVwb/s3Lfrb5ZHvNwRzYxvIhLmyKbeXvdOJ11nkufIfsH2HIU+qSLNCX/9Tcnb0WIjEfMtx
8jWmaMd9wTwMMRhcnRn1BUigSEzjhPDVqPVMLnqcEhjn95gPi5IoB4McBPvliHBtr+VVgxDbJ2cV
eR9H1GIKkoQyeBaF+2yHjdvLXKVdHnyPjoTzSKn9Tb1GjcpmXBEfnD11f0IhEAE5aKqxtCrCwjCf
9P99wJcSsozrJGBKz8yB+7rCa8s60yKrIKD+2hTlp0RyUWwhkI/qNUJ2fydfVQjR41JxOhYLlg7J
AhHRk9mRaZvJMjPQVJQvgKSZKFiXpW1TuPs6/H2xF5wOf5lM8JUIsDxxXHyNYkb1XKVHgKHb+F01
NKI5J+j+PUxgINUsLf5jBrXeGaFzUOHAavHGiaQ0b6gDDwYkZMMh8TC+rWxcsUVErm/e4kt7HEU8
5NRre9FmNMR53yi3sfIARJbRD97bTCAfFifiv7O6awDuvb7aO/PkkFbXJ5qdu0egoxvxc0goMKty
EOYEQDd9DLYS2OxeDwqx0pCQvwqZ/uRGqyM94ggN91/GkRgDTqgF2PhsnrM/aN1JmY06j3tIMiEr
W/uhNc/brnCHmzaxEfSFKNcqbbkkIXAMWZsP6I9y2s+O/hoxCO7ZImR7pZgq9p+PBAkmDZI41m9T
QxNbXC/Oe82frpDHxdZh8hKmp83uN67XAmNBCRIjinMEHsrQGqdcyAVFP8c/NL8/pMcjmhc3ltpt
fAeGZlI/euGJ/GXM1THXdDdNqZZLcqPjD/21GJQY3IFGFDE5/Cpv55RTNqr2K+y1dvsH5kzVkjgm
ij6w+sqska/ETCsadbNViN3nJPdPxZrNcsnStgvcwtsjBIVVAWws2v7WSaywviLODtWzcG71j2bb
wyq0pcYQeF481eLuH4kNEFBV92IIaThuyYGQgKxwUExZZY1RA7ZckHsIajUI0fr7RPeEVG/rzfxU
9Jq3ZVTyljlFh3YAxGSR8IKU8t0kfHFIFXV3pQ0uBiZvxQe621dLuXbWfTuguAS7NSiUyyD4Hqh3
cb3XSTvZ4t4QkSvj/IysiGFQxvqEkyUl25RTlncP8Zz29qtJmX/etOlqtu5kEtXlioH8hA02kqFS
cFgWJs8U77ERyZfuU2hAJoderYVhHnF821XHnG1960hHIN1tFzp85VkubxaBGhAlZTar/kKRo2RH
x5ufHRG/foTh+efgvccllJI/XrhmPh+Rnc+T4caHy7OhVbVPomrH0gMFrc94q+2Hy0Dl/Cc6fTa+
jJIbjGEtFa8A3udqxm3dJY7iO38ZjjSp0XDHFvuaKwIOcB/BzPFecF9lxo0svI1C6df30h0mkm0a
YtedY93+A8+MADZ7lnNw7z6UUn00Vq2EEA59JGDHEofUAamzqHBVCjieexw2zipA3XTPQrY36Nkk
iTuvRa8gMAUonec8gM/Lcwnyh2/TeKZHUvbkft2mEzMw70rwweYlCb4L6pg+YJJ9RCbRn3YFzAWH
agG5yUdTR4o7Ub7c7G6epkLSJCCqxdLH3XLxy76x0/9VhxjiVDQNeW/qoTc4HqXX/eojDZJwRVJZ
A+sbGpQmVpYkQcsNPEToHrKxSTyMNBqPbfLlY4AfMlmcnmks+BtppwFBx3FLgmwYN3SKY4Qm8cqw
whdBn8NSPrLjAgA1YSnZ+BrYZ6b/QdoxNnySIZVA4xSMx0wDcOozkEZcwUzDgvW/pL27COlmUI1+
/4aCbaSAYBfF4A98v7XGEgq0tKMsa01Ejs6JDtlVAxnEG1XPjuJb+S1C+am/9BIG88U6IMWM02Ys
J6f3vfhlVt4vwydCzVDBgvFS+52q5PZcbw9Mz1ZUhS9e52TG9JNAycFkaSuvfE02ceXRKSw26JB1
Kosuo/ic1zeQ/rN5u2l1iUnPdU7UhCmmq3SJG0MWh+vGKO21Yj3axWaQCrrCFPV7gqcL3HOeIALb
8aX0+kuLukZP8APP219gVC1PVv/zzob4x7mcqK49ChYe41D6QUhelZ4TsF4QBbzMiGNOydfPS0Yr
Ds8hMf6PiAiRETHDHjdcCGPeh0dxhuqLNl01Ejz1byEXUwXEZa/4w1xnU/GdKeADi6EddZX3KCeH
gxBItGv9SGuhsZmtD9thUims07bV2m1Xpd82chZq9wZwMX97msAWD2hZkqbHn3HUGaKP7lMApL3Y
l7Ptlzho/oYpcgHxWr2x1CNTyhVDuLzAyhv2ZgX1Mp0BXgViJtQh0BJjUDpuK9WeN4TJkqkXo/Y0
GlqDUdXcdQ6WYNXkNoVI9PEZKAW/TlJg+oqxzSfF2ynyRwQEXPwT4tzJJxDrgNTZoENKenqi792A
5oUbuspzNBZ+M+Ne24cSQKTWITkWggHG82obYuNFwyXYJ/DIdDMLPoC1mxok9jwFpF1b7R27SbN+
pOorjHFuk3SsjAdWH/yD4SSlJZBHR/I1AYf1075By/DJBGYjyWe4ukFCLCwVXO7+JqIH4NHOSWS1
1pSUSdb91jV3y3kCLZCjgYWvQ7D7BDHo6D/b9tdIu9EJeby+3sKXFc+IlCXt4rh6dSSwhZcWeRuU
T3WYPJJNU/ThG8fjGFhcgW4esMVBMNjf820IgjGjup6ovvdC801zbZYMLJJQRSZNungTeoH/kE1K
5YSCmPw4EMN0bSzzzRVOOiEise09ZYSZM2vFuB/f9s1/I/5TbQeCh/7P8WK3tR8lYGLPoHEJEun7
8RH3Qs2yYnu6Xh1c2B+5ufth9xdW3+vorhNg7ct80HPCUuanjJImYxw/l5W3wDAyx0zyZlse0cI/
hBr9P8uXUudxKg2detkJjyES6ZnwWHfM0wT/BIis88kUvrfctmlUVV5d+RtWIkyOEUshuF7PMt5j
uviVJqsEOZi51PcGEcuQ2ypnfyLnMbYl7QOOEplD4I1AOr9m10nSZgl0cSwjWScRV/7WVAPlcw8z
FOq2+cJncE9OUlkVXSCG3Zz1s+cFAvlv1cQQ7LQJIIAq8FWVPnSkEtILguhgoWV5J1zvD6pRKV1s
g0ZDQZCH4p73CvLZC4QB4qYrebwfPemixXX10Tc/Vo2jAW6GdSpAT6xOXcVWMjVDPxwuuba/JUO1
Sim3g1OioEOqQ2QVy92puEpZu1SdxUO4Lw03gZ2F6R+S6dbgfUIMHos96AyrSzckFPv6Ocg4c117
vJGN80Mm7ML1wTQ7OKDLIuzApR3sMuuMmuOca0noPWy3bgMXRx1lHtD+EmbwA7Zda4qixiuf9OQI
/iNe6ISpegkBRms8Y/jcIgVNCfS66bNihIDCfadEpbuvTTYBClcTHn2uue/z3Z4jl1gzqOG2vIgP
qsujKw04aXmNJauFaX5cxPMos+xO+h7fAeX54L5ZxgH9s1q7UCHKkirx5hiE0AkhZVWrlmp6yD/X
JIVcKXbNuQ7SssWSYJToMSkAtMuanPBLZpv99/324tYhE+zudyA9vy1K7Pnmlf2mcFoYUFPkClVe
Duom04ccpDRWIHqI8W5ol7tJTYtog3KSYs+wd6UoEfM/2S0hk8ckFgPqtF5y6p3jhhaEbM1Z8F0j
CtO/MphL10ccFQHsAnuEBechVdk5Je1hnHjM0CvfNslciR30mkliPzegg2Tu+AO3DU2r/WZC2wNH
e0eWrEElJjx8hZ0k556NGz/431f8xgMUpDArXihJ8GcaLxw4D+t9Kjmp2UPxnjMFPqxABCiP9AdV
lnx/5KGfcjn5bc75OZdZFxQK/ti3m4kdei5D5Jl2e9XfhXMpZ+pa9djypwtXxSiZOCErVkND/ZeQ
M6BKM3LIuondmQlwkOYNQn2ubjB2Eutwa3ec+QCIeNCC9b2euUbvIwqXzQ6fDLPb1/ZaSJQoA6Qg
D3FUEsBRjgMfhjPNZPmrg9jADGnqkbod1y3FqaTgzbICnSjHXV8wiAqHNNrpg/ZhvLA/XarXUwrC
QSdZHQyzn1DI1DGvi114fOYxsYfmgpEh4KtTs7NOhLrmE6xSr0B3DptKeFi+m53iMlXDizSyB1GJ
amk/6Eu0rfKnMBXS03CO+FINQ0My5clQLhw+hcJ6MA3Crgaoy7OYGBYZrprjN8Y7fBztaxuEl05z
G2kmRBWGv+YpgVlrTAat6CCPekWBicLQKH8Mji3qlp+2NogYmZp1ePWQw5DbyCLNy/uRYg2NUk+d
FORT3umQ99Z7fQU+gnEydpvecrlfq60dMAhPeAbEJ7lamujfX18UBXRqCUnHweTvCQjPHcp6Fvmh
wcUlBSXThkYKhiZ1Wl6BiWG39aBL1IPcfbG5d/3dfE16ZgqUiazMJlBSBDLIb157RcWYUUvZN3Nh
suiHvPsxU2OqF3ZJjIW8zy5yIftIWdlJ0ynAgzvPwFb9Kb0TzPONPQGxczPIjvJFT9/Lep0Cr7Rp
8dZ/KmGYO1Yb0mAeWwLt8ddukdWKtdkbViyn4gWMkdybXg2WveiunJHfwfJD8koYApNAsfYU2NB7
6ZxUhW3OXCq6rk9TlW5eEk56vTLSgiSMBkGfdjbMrRwlLioOatQ65dduC45U2aIgLcuTKiJsQpNx
k3AwOz5IRvQADKRTx9RpeANiuG68Go0L3hePVe8cJLAWmOtrFZFUnbIwvJk229R8rjaaN+vbXBx4
9CNsAW1+FYXuftLxBOrEWQpJCyGe3ximPs0NywY2KOL/jMm3QtTlisVn3PACpD1DUJjZ18mkPGuz
AAIuoIWUVAabzGtcHAYs/FaaQu8dPujPOYenrYOPSVoPxzvHotawOR//zqSHGnh7v3ayNqLP+v/x
HAr9piLqKxrHbREZOOaUTc9D6iGdNAqDuvRe+Rr2he++pmYrVlfjog2dvFBTN0iK5fkGuRixlYQZ
JDPFaV/cvQM38h3Eb4X8pXHhh+W55lD8YTUUQvubaPPyya43N6XWJo6sbQK7cRzOm+j0Jkc8cBsm
KDtoYrK8NnFcDNeromY3CShzq6hK/ONlje/sR6fMLtXdgWKy034xan4rz6jeLNlpXz1im8nlKiKm
QYPEGiBmxc1ydmfKt8kq+ESB7tehUc2VGdN6oOFR1bCALxHyX0M58kUw6UjZwhk2EkYXLNurP6vu
uXY43FBZmmisEoU0uGCfQOfjKHKqJHmG5bu69fwZ3DFRJAHJC9z6SWtQ7IqoytMyLde+iRk1tGgk
H4HralLMTC9B6p2xTYE1e8Vt4DG19U66Qj0wmZLhjIDL3uBVp2KE1KJcUQ/b2SK3GXvcUpyZYdN5
2qsHsYnl/mv10t5PcH3hWIuGveHYSZZ6hKAY1n5Vo5721KRK19yZ4wuqAXf03xcA8v9F9st0cTDa
7pFYtbWePTyK8bpyM0wWpmkOlVg7qob/hB69b9xQ4kUQq41QTh9Y2BEaGWyWnPJjNSeBhfEHPuH+
IVp0op0bB+Fa1PjrQFioVmQgCcH09RP10dcY0MfpuqKGvoWAQqFaMS7676QcGz2SksqWNXRdYBVz
GcIKhdsSDXWjs0J3zn0gDmFC5OuI7j83o2Lmssojarx/GWqFG6Eym/WgQ4UTPWEnilhjIi8bd1XO
kc36oisXAQ49SdvHF84P89YZlj6h5Dni5K8h2csK61ma3PuCgU9xZQzsPrsmpya0pr9uCAi4v8PW
Cc5HQCP4pBmaw+TTNfPDhgu4UZ+gGXClU0b7AOIcvrLTSkojY3Swb7T16Xe6kece2qkeIeKO1k9c
KbkVc4d+EfXW6n2RtJSSkHxvFq5yiMKdiAnWAsabfDk/C9OJrEGvGJSCIbAQyFJ6aZmDcx6YJw7I
dlybH6R5PgtyIWMkWKqBsd2FARpcyeuyISrqGzVYPpk67t76g7V+mcM2CIhzNTPm1dr6Oo6puaZ8
3p6tnx3p3s7gEAaDXq+OfYRsj6RzpBT6vsqGhXbHAdiBIDAWOEPcfPJM9OOTcsAhhbneOv/iP50W
LiftscGKZINgr6tStWGlaTg0/LvsgNGswd8dtM0zDqkTwt75VIOMX7b8623CMWzo+CzhR9aM8hrv
BEyU7wz4qL1GAZltOshkEO8piuwdCf2b5xZWS0UXcPrUxHBEFQ33lMidVKP8+/2mCYLVtiuApawV
4bKuQU6r+QRQctqKJakwNkjS5j0yx8mgqm0MGmRn3hsCkjxCIqjVTIisSyCIAHbVTH3BjM+hJGuw
Zh2iJUDPO6PptZfm/eHtTHeZ1tnQv3F+3C9KNtrS35FGWfKZJwHJrHaw8F8GcGA2M+WmUjUWsJcQ
XxhxCdvXQTdKAHOQRD5roLlTaL7y+8fkSlt/lFgloUAtm5JCDfvsZfscD8oR0EPQXPSNu+T7L0d1
ItipK0erpglq2nWu/OHJANSmUqZwbBUjZGS3z8C4pUGrWJjgO0l4OhnleeF7BLCOeMiRBwuOehIX
ZlG8Q2XiJx0MZSCz4jsJCRW7RmnYMVSjKJXfpeNf/5nys3k5cthatKcYSa2BqCehSgW7kPwaRSN/
95Pf2hcPjm32YqpgTSXLGKFOfBkRwC7j/3yWEOBA0JnshWfEhksAjKH3BUiLXnea1ES85ANQtrKe
z8YPXPYdMcSvzU0mVwTmrzpQI5QLDs75Ny5fUYSnHZYICYbP5q+UPVJiXMKdpRF2C86Bqe6KeOWE
YcgrlRNrZ0WFntGyG4vVrD/7/r9M1jke6gSGHhfifWL7gziIcfd+/C0aCbwt6e6qr8LQ1PYel5oW
H1iDV0akAWw807vfjbOnHYTlrBvyUkN3vxQpZwrrW95x4lwwMbN4Avr3sebicTBXuUD3Omk80RIc
fzxfb61fuqMlk1msERM3bnpI1KgdzUsz3c2dHt+cwKkUPqUdEbT+Mgyg6CO7smGHz3CrOTzLcQgu
SRL3PJhFJFBDk2neMnnCQVNBZcNNWFBepk3CeReoruksDK1yHL+29J4eiaEzsemBwU6TbtZlWMUQ
2UEh9pyw/aERH1bgTY/89+RpqeCsl6t6SK2HjAl4d72M0Bu602I9qbBeG+XjDCV9fSwokd2GJqaw
BBLLTh0c1tjQc5IdUuL3KcT8d1zMI2sdKFDqw41kz/oBtBcOj1B4v6a9fPQAtjWH+C+jJyvmbKmt
meMReFmNJkX+BkfoYam0rOaO7qK1a8KiLg5XN5XPVdNM+hneGsc+hWTnhPJdI/0wt0S/2v032BmF
emxUNyNUaEDgWnvBFBoNcQb3GToJvrIFmf1vVp/AGW/SUkVLrIQHZmZiOgvHz/PZ/0gA8vSBSSDl
BTNG+szhyEW+v6jiJHWNYAxsKg/LKXRRueOVpxRrDpiLtJtKvWxS09FHYp4kCqALkXBLRncmHKlV
wo7ekvrdPLgpZqJlBr+Ni7nkmqz2EhCkyR2DDXrlBs6LqpASw6FyQjtdmEfUeZ9w6ITuryYc7vg/
InX6bsMuIXiXI0IaaCRH6KCi/7AiebvIkZqcNoeKEFR8T75CfumTri/GnLAdwjukR2qL7vZLPgI3
eguQgh2YwSEdY2oI+c7PcxYNH31bhOrVr9hy6Og6WZICZrqG0A8ey055djRs6YN2966OevP/tluZ
j2cDBWhexCMlMofQgYVkLX4eH9Y+4QhpR8INIOsfhR4ldHtIGC4g9abwHrnAtCzFPjzmPmmt47Ce
1dBsDwIzDaiGfbUIzrIHG1ZfLg05mWQxd4m9z27sAZep+gj209y3x8cgzDpEsS4y/fVDA7kLRaad
AFxDo1SLHVi+3DnrQkxJkUDobrL5k9+V84EDeMnUFjt7vvuTz+/kiw9fNb7cNYpQgWVL97FXav+B
vKBcBQNGEvKLotyDj5Vc0wETjnB2ejz3Baz2M6nDi8tyVForQnjbWVFGE20P6GRln7P4NGX/GTph
KhyA77f7Jrh3G+Ifek11KkkiArOk5rzUIJfV4QG6em5Cj01TYNQPV/GrQpe/Ve7Y1bCBixpmMaXB
VrWGm6TyseChr8jSrFZyQLVNrNQfKHH07NlMMMrWkwaK4SQnKlgKj7MIWToadsItRlaCl7bDhu6W
AUjJOC6qB2DgK9K5myNu2IourlSp1iPjAwDAqIK/geBfZiZrAP2LZCUjl8aN4Ft8AbDuVnqgNyMk
YMPkd7cRKnxAIQ5I0Ml6sk6HwIC6cKbC0xSkeaOhdLbvdknu8DLcJTX22jDzgIFwSCt9+wXWEZoQ
wxF9lbXDVohjbnQtD/TOie+jFESzqr7SnGoc+F6zVAIvli/wwliovR1VmEHbDhCuPfX7azOindwS
fPBbD7iHM01M+d8Q02bw5JhSUu7D44fZWfb8ouo0PU8WcPHWO8wZpUwWFi85RuhrZEkrI87R15qF
LipocCaiYGJNygYlLqULFv1dgl/iZA1fyGUfBEzjHpSUTPmHh77+p0hShnT4HWEdxrpIclYz0kaJ
PX1Qk5O8eSOhAYuKEeR/mv3y3e5ouikUDTxjrlR/zLGZVYrVchW4INx+O1fCZusrtB+etk7ZvOqq
dl2hD+zUKgSO8AZ10GcACMA21UQpwYEr22J4itkGrM7UARrnJ8kiInI762k4lQEl56HhRWMH+4AW
mhQiPZ29bQpdtUIUxsylU1wQume/O4Hx8q6psWi88STp+vUtycUoDQYJu0LDlkllfIfifhxYARWt
n+nZ4mUDvvTgGzv/uwF9XVpA2zBv21GXqd1wwGE4rBGIYYkEqY6RbBu2akWygs4yN7bTuQhN9st1
/HC9m6+h04fieG4qTDiXePkznjgJ6zRsU1+eLuR2WClJ2TVA43ROL95BSXuoUGqMEMtiN3fujyZ2
huOmmqrpDKitEVG77ufwbb7+oHzTY+ndjMLpNyNg/nu2JEntwoy3xZygHITJhPTmmhIiq3GdBg3x
T86hNxUvVli7TDfVO+ZlECtvUZDRzIiENgkHuiFSJ5NKb+qzSrl2BuqXEVGXIzoQGu7UtbIdZ+eI
/nW+nawlhjEZA673nPDbZMBKJm4Pu5YssI59+Fsz1+ejj++LtFMGnyvO83ZgxsNzogt0SDCCyRxx
Q3Ay2AqgSK3vmWKlqbhpZLjjvOa+qe1UzgLkXHexp75i6FaXQFpoHOn0TFsgqPrIAC49gFpzG9U7
eZW4pXguwwQDgFzlhGlZKUHJ3vXNCEORDFpv67YdcvTp1Fq8rqQcus9vyi87g65H7fyXObI8lpI2
AX5oybDr2ZFVP72SX6uXmqqbWkz9qlnnXCOlndwQ3KcP8vK9fxrF7tPoPCrStU0F6gSA5qErnBYS
26dQbFe99n5pcLrdS2A281/JLdxDXn67TTo/ox6mz9dCGmsKL6pzk9wKagbJwQ5XVz6Z4DlE3XkD
u7LRKzBPyNN072WrZ7pSQXtxHx88KacEM5EjObHMR3zecJt8HGmDlOwGSE9QtIKXzS6D2VEno+y4
kT+ku3jg88rvlOA5UDcIpAVXzlxua5jjPE09nEjhtjq/Cc3AffKsxkzK/T8ubqYn7Sxhn0OTVvX/
R5KynoNNDaXIv7Fi1KHp/k/HNgnFgmm4vHmCQnKTryT+kB6VYkBqEKELXteq5omu0tmxVFHryIm2
ESXicyn8kWiYybAtGOzaaoIPyj6RYjHVoy5dFbU6j1D7/W9tGHFfdR0154NToFmRR2VaWAmQz1hP
69V7OAUcwKbRzXmgYVdIRRWTccH786+STYvR9uHX2jvVQxDvGM9+vWJ9EdKq1/4EtDll0fjitazr
pAytPqRpXgsvxQIsaRJ8Ul9f/aHdJoxe3WhlUXxPS7ks2Ky+zoIwcj713uU95jxEJ3JTpsHgsBX7
wKG/Mu5n5FU3p7v1xJgdFk1WJE+7LdaDWhK9B8oGeoOFddqbpHaOCovkde9rnu7I4c34l+vmJKPg
R9xfBysTbqeXEQMtvzFEMaSU2elgFPdWJhhVQP8vRkYZsxsZcxezrhUAZzvj1cMd8dswQ2cpcOrp
rFGXrkGZn4k52jScQrLZLJe+YrCSmN9j035d2jzoA0zTlMQZmFu12ngwYspwpUmPpXMSl17WvapN
ac3bXF99aUjJ2PDIiyxmraVYBAUFq9/sOUwQWoRRhcw1JkFHOsIGX9q4qncw01pEaPktiSv25IxN
fUqfCV7p4LRHWsKyzim/YMxTDbvYQTJL5fgj5youTVhfTV4bX8DmIca6PVv/DzBoEv5QK81V1iFt
oenJAUfXlCkKVibqzo8WwAuBvcgEQbhRSqglCsd6Hh9amquYPrB0VZjEKxqPXFuT3z0U3Jvw7Xkb
OyodbMhO1cYjbiW5GUQms3ivbckIoGc5CKc5+3CAU4CbiUqynJSek0OMNBXTirF4t4d3e9nS8Ydn
SRtNLWPpK+HbtIsNHwWKtOxRV5Y5yvcVj4fwiEV4/V7kGPkUyMgxsSH2DkwIkitk5Dqk1kkDCvlt
9R7OedDDMZfF2ON8Np7MwBC3b85EARSLZV6PBUMQGhCnovwCjlD50esfzzmKjdoeo0Gz64brnHdO
8JpkdlOVHLfL6julwN/8D6DCFTsGpBslaniLRn7SVg2ILDTMXzHnQV7f2Wh9Q20dsnmJeAlXXOLk
Q19boLlHy4NR7aCQPxq5sri91i7eHWaLcoX36OhvyenzEMOorPPXgQt0Gii1XWttDnDVIRfv12ue
zZ5pU5bx/bLvXFFOp5OnVBh1gpTDaSOYHFpqVHretqxIZ+h2yfDz9WtopOi07DRBEz9yWsZ1bWd1
l2onV2y6kMhfi/6mewzeJi8u3ZLivaRrriEmspG5Z9qcG3vNP1QIMa9H/XAH/ifv9G5YzXbWBpLH
h0zzUc17QpyKltMTcG6/x9HXkHNTCL0wGgJ1u16nyL/vkiTElj7w1zd2ReHaXgBFHo4j5uHEGBJA
0mqe9KWglgvpVf/KIzTvFaKK5Y+1wGWcC+lsOTimiSbTIL48cvrtyTiMme/1LbgUPI3epSHc60rv
of9TLTiM3YkI+m9n0+pz5twxr6lTDdopjf7THeRE0UOGUfs8B4IhLk1jc9EQRnRg3QAWGCZ7nMhh
olUf/Kimyss4VokxtF4f3I+fUIRoiV2ea8BeLJeutrrVfBhf6LpBSzmAXBBGrjbNY6AD30B2C7lV
nfBYyU2FBdQekZK9NHUSw50kQUenyUp8SJfS8txBpZ8853pn4T09DvTNPsWFjQEbTn3LWy2DrYGE
i90aCO8C/QBwhH7mhpXGck24b4uOmRKF9kvfz1FoG3LPeEkZHy0OuGe+y2RW1C1xtjjl/sibzduP
Dq7JDkIJ9ExfQD0gTKRYbZSaVi9YHFKw9H3k/UBIwHEYwwlS3cw2wY/KmyqgEFPi/MGXj3BUduq7
FWjf3WpbXbldkwULwxNg2K2h6EIIhV9tUJGZWTTHRY+cYwlDK+PPFPdrrJkV5NC9SKkgHYss7W+a
MI32fl6/5/EvERc6ckKloNOLlInJ9VcCEkcjkiOrSKKzLCT8ezo0NRTp20gPLuB2rr7z3eh0EMJI
1WvZ5ikV1BaS5OBMzrP9FeIlvPXc/iVuYOafeYxf4ysrR6j4d6MWpWCf0DX938JOWzqtjfERJdoR
5Gu2HrMO6Dr89M1z6SvKSiDekqBL3sKs6fdFEGWmouVc3B2kutM0k7wwbFTpn5m1L/fwyYXPJmmj
O4gbDilmq5ZyOo7kQ+B6W37TCE5xUoRZnG43a9ZWzuuyHcpyekKF6Z3VFVS+ipHn7wxxIS5bRxwu
Uycj4Sanf40DipWQbW7CFqZhG946bTTfkw7IrLGPdRLl9Xe0aUIhqNEAK0/e/9cur42LgXkNHyUv
bHQbgEfC8X4Eo9NZixqfL9i1kiZ8Jv7NT/nRbanhJQH2FxFpNd2aP3GqMmWqPvV/XyH1NfdJ0X84
Ye5GAkp2ka4NSzniZDDZD13+p2lffXfOKhwp1zH79eg8+c/rY1L7o7u+xBHhHGV3MS/N0sSTnwLx
klcMqiC+l0dvGbCVFncjavUPLCodHMn0Np6aiHu9SNjXJY2ZZl3kjivE3s10U0F0OvyMUsFu4+F7
MJ7xhejDnDHu1vGTSoq+DWECoxr9OsUJXMgYIyZjo9yIftPCgtzmW7IOCJeTsHO9lahJdeIFQk38
tDcwOSaqt7/92osiXHS8scCzyzHdgYlg36N8MVZ6mOxTi+f3kGYzWvG8njTX5W627WC/Sd8rgnoU
9N+f7WcrtxkKh0H1ijJUMDGGmM31EbaHmsyP0L8DeYuVC55WbgU7BRPV2omUDI3jUMvrftK/PBqY
ZCRs8xSm0VxSmRj+NqG60EJgpwuVb2CK7uLSQY0mEJWULFQuvOlHLYrRWbfnpqVAD1juVVp3p6tQ
0tBxzWZB7Qi2wwtsdedLBADEcATr0uXGYb5X9aVHE2463/X7TRCzpifkerAmucNLbvgFgPmoh+rG
xx/Vv5lbRN96hBPgbVfBc0Sc6v8FkKROyxpqrq7VAzXx8OFnMwheEjUNGmNrx42PLwXywqU3Bx4t
ms7VC81LeO7CYe79ZPlk5GGZiocp78GrItCGz2uGazroPStWap+kgCaoTFyytPTicI96CVe+NlvB
0BrIfXGMbx9/64BN7JlpOgrKLjvvQyFxHwHVXgqTbagZu3QztX6hvOZxLJ++P9myeZ/sYDRu1+2L
0ISShalEYlplLKzmpnAFljWE2n0qbInI1OkzWgIf2nHVJAwK1sYx1ybojADQ423Gc4FYAq2npaIP
5aiWQGbgAiyB5yDSQPuRmojL3j5D7kVGY2+i+3rh7v3kzpXKxqCuQbcZtsgpfOjyxOFqvLLJAtA5
ZzpjzKqi3NUbKscdfYlYCWkRCgw1mr4bcSFaQBYLRubNobB28JSuhwKusJur7Fd+7tEerTv/xooU
znEV3H9mopP9IhyhPxiFrvHUBRS/t7Z9S1ViMYYMQ/HatyPL0We3X1RANUf2F9jk6XpOBU6DPyCI
XnqhE1/Nik6FpFXc5LGDF8d8iShgb+DJ7cv2xRkCBGuR+WKQDpq2YXgx18z5IKkd71YZR0yn8EVD
sdlJyAxZeDCOz7fjgtOYVrgppbf6rZHlV/78737LudUOLvjYPbpr4GYWgDl45eO65y7s0App5MPF
rO87+cxYpVe1FwAzJ/aYV899MVdMTI1yWAdQO5AggxMpaZXghbZYQqnu32HLMA3gnXR48EurPhkt
5JqlhHr6CKNj3hs4+9kHPjuk/9HdD/09rzzJBVHOhjwrt265c/JyjTkas4KXi6XlNx/4VuhOYMWK
YtAL3p3GvdoaAp7oGG9sH9xJ0VYac4IK7Rk4uK+jm2ngSfTVc715J4l6koD0FW2dpHPcCgEDeHWe
IR5BPCeR+jyMDeYb8pYi9LN4hAMRAjGNyGElqdaVEDerI75/IllE9/7goj4pA7TnqDZlgDFlnCpH
Qk+j0yXxtas3aN3gQHuFj4M/Xq6BmbS6E+vpvI0DNg7PFZvEYrE8NhYzpM4NHHjqifjxBKNkTXga
fIK7j3howhFWURU54zw1AJ0NZjGMIqXZIC+pkY/VAfnnTmh9ngl/zRWIrhRXMeXEwxlaiJxlg84j
E9jNNXBXMVtvWkdj3iNvAmBh9lZFZfZbt4akOKaYLTBi6iDgcD1YtSFmWGomfBg8s8YR4SA/A3og
litrqeGYcPv6qbNvGk3bhpPFijXm8YR0hbrGtdc/5YkB3waZHIqwpUbgLTztybwu3g2zMhl2rtF5
nLKV+Pro8G5O8eLy0ZNN+v8Ub54PObLhwzs6DWvuTGop7rGkvc+KNufc7L+awseqwQlRiBs4o1qs
gXs+M7V0nIR6riTULNtN+sCem7P+b6rzlei4oj0uofh8kN42nyezYmF3p2gUnNMYdJ4+bgmWotAO
/fIyOYTN9y33W/R5rqLeCZeqKPACo16EuIBzdWHMkXG+M0lX1FpyIguwNY5sf4RA2QnQYwiF3MzL
zFpEKCLRMyRNfAYapL3lfbCMeuNJ0iuOdtaVVTFC/dfKiMLUZIdCI1bsVN6bkfsg8CxKUf7yeFuF
xcTc8UUced3K6vIaaETqGkPqDLEz7qf/uPU09hTtklqwPh2eZ5TGq+tTq2DupImkEIgQafbcQSZ+
R3P0/D+pIGMAqekNfiTz98aXmzYUSHd3ZtUeWkQ8DQO20wBFfXSGy5aBPYs2UaKIKzudZ13CZt2U
xzL8f+/cBQCVhqgP6XI16A4s3ONdyFfFHgIXQqLiFBzyaBXCHwWqs5rj7jabzN4sVloeyBegTwdv
KtIeU9Tkz8F93GWMJWeN0dZk9bbWG2UZKpn2mfGRJ+kSrluPMCCSsIv1XScxBMaeA2kh56fyuYQe
lxJoHtTgtxvxJxpxh6bjYP8+TXngSgCu5v7wkuJo0ktsWn/BTywDjpOrOhkabg96fV7MhDyvyOD0
o3ouUTi72u9cZNj2ahG45Mrht9zygSLCZk7MoehVr0Hn22rb7gA3abXumf/M8JCAbfsYZbTlTKn0
VdNhaqC1j9N1GK+n41OkWBp+l/T/47blCgDfImJNyemAWweJYv9t17ip4WJ+5wf/Mz/wibga/5ZR
OtAbHDs19oyrDbTzQ8zx82aL0XtjdldBoWmWIveuL5etDZ4OPV0Kd/vl7LjwVl27bf0pkS6YLHq7
89cQIZA6U78IiSVOJ/vzvVDpqExWitrev3rmO8rjBq+Eva9OuzWE9P1agMCMiY3yLSdTwRLLPiC/
T6lQfylcGqIo5vsnHxsqxpDBDJZmNFXpHvf+1H4dnRfHEthsqR3xyLDbon6WvkbbCQOAG/OSJod8
v/wxR30crLDyia+yduHmYAEcUya5xIBgxWfthb7rEywejA7Cen8+6b1AjAvD2xk3jcbPLc8eGLIs
N6GI98IE8KT7CNndxoNTLqX6wzrntNPGqK8m3GsvlqAyI+qwR4/04uHt342lJXvPi37/ztUMq1nO
InF+SLF8KcOArdVpSNNJSWoEyaxKgl/o8I5JVAN/TkNsRouIODd9vhp3byWwe424tEYJCpfX3y6V
VQW4O3fbB3CJd5PWdebZgDUQ5TEsm7YgSlqGqTotXbHSvwXC7ZHj4wbQG+cUv4DsALlOIYkpF+BI
JAybxE4QLs/GugvfAe/UqqVst4AM2V33xXw8yVCng0aKeluc3jTKGmMYEcMfjJCkogfj2U1j6zbY
+Pt+PWTTfNbRchxPdDqdnRvkwKB9sSErvBdqvqHY3lG2qi1I4A+e7VX7Byj0+KTuifB9n+cMVWSR
Ct6H+sQIaoiI/Gu3/rkfkDa3Dm9rrKYcsian/z4bDqTxiY5if7SoH/lInNezMWnqaHYPweLU2s6b
9VKzl3aXz/X5aUODqbpXJN4nK5/CLUmpcBvPS17mx86yne/24nChKduJULR5Rw6RrD6sr4q4ZYXx
dk1FVje7ZrzBqGgphx+NUpWGdu1CTcgKDr4uvtGb4oXaFjjtxIOYUMUsIa3TAtJGUgafF2f0ZHpN
VD6zq4OBs5ZGVmMBVk8wVlUEZN6CokFWu11S/5XUekYBIEtbrAORC6vRG2s8WBG79nis1NMpCHE1
0gPKiL32//KxMPPkkDFPgbtEEX3JX8JBwc1OzWn6G+1rw3PX3/Zs9zxZIXY1+pl8CP2Tgn2dxt4+
X7W4tvudTq0sAf9tDWPmazFObrFVB4YfGB5OtU1ekBXy+PNW1Cg7GhATzCTtJin7Eav8p2Yd0X6T
pJCuB1PlZokRzapxLgFnlLjdyF0uXOEI85L9J6fvc3EflDtGFROvKH/vHWw3zUeZJmGb2aG5C9+L
42NA1KNKBrP5Fwo+knoqoo0TxPpZekHQxEf6y7mAFV/N+YDloEEOeMGglklKrBjB/FB0mRXYrSxw
YLEW2mR3stu9HK7qKChpy++tiYXm8vxDdckC4OWO7/zhUPGGrean/C0xVAbdh4hGaFmpxM7zqvf0
HuLrQHEuH3+m4+hGFnfXXchZUcXf8khGo+yNrXQFZ59MWEE3s6AZsS7d977vwasUXLhR0uNqOAe6
VyMWIwhRUDR6DXMWVAYCUarPNNWIE4bL+HkddkQu0KobFhZPry1aTZq5Xg7zvUBzU28sXf4MHs1i
TUG1ywziISGNGwHw+zNPKuIFpD7z1m3L4+ymgb4GVyS96N+zoeB+pjEJrNVdpXLv1r8spM73Dfdn
NE98fDVcEyDCqA2fmuU9/4hzB/aTd3KeMRWXpiAK1kzqjaJ5pyRHtjZJitEIfAEcfsK+ZOp+cfAs
icIAfsbUEH2RRM6SO9Oo6pg8ZUA8KydOC5q78mBSwQ7heUjM1p2VeQoTMaQCaFfYEGIkuX3qtNmR
+EOgOjjLzZWG2grPQLXIoSeKLcmUtyXbOBGqXd47qHr1XBwhY49FRrfPQXwJ4ciULAdIMEvqUmoI
iSC+x5h57bK/3oKevS8amviGVEic0VWLkFQwR7EPOmm7v34WAJjdtXWrWHYJOiPsfwzTKgOhNxcE
X59qnt98lP02r2IznTow6MkxGyhkCJbuBSHijsuREzV/CkcTVWFZnshhyNcNhHMUwrMvjQfyhEva
0VhjhL58D6wJYerjfOcJVUzKrF++/h+pEijm7/SMNGFLfPPbkxWqaNiJLAjc0q2ML2tGs4iiRSqK
39ovP6WtZX10JWY/N6VZgHkNLtk413vQ2Kog+hIvFGpgQugZ7JSLXE8JOpQq2X0FuXuJOTxsC64p
7fExEzPijU9sy63I4lbSYGlw5YsO2TjXotWpyRHDptx75ynr2Km2W+LOUv56aMhVZYh2oEBb1b/2
yxUKkfPBacWLa5Odd5JoIhg6A3Wi4Ezc7yZvZg07YGsTTq/cfaTgVc9qcAMop57og6OYXMp29hkF
YyH/d2QR8gW1blB18YLJfDfSWw4v8oT2/y+HcEF9xCXo9SwhRt28cYRsj3z+53+hy5ACx2DgJyI7
RkTWapfexSCuFqMxaD1Ducs+7CQcraHDDrO8pYKoJIcXb1BhHMcRQtAMihwoz7CcI2Rl+tjsUa1Q
5TrBaIkmpMw9e0D5nHdBjeTFbuVXEn5XdhDCr/v8KFiVHH5ue6R0o+HnrSatcIFi/SMEHm/hz+TS
snpRnLjfPr1Ijc7VnKa6/C8MZMpKNd/fiu5cCl/xl7QsOiQpeUoWr3Z2zJMVOqzRwoRQXixHT/te
zzsPSugzy7D1Gv5M8S4GAg9dZA3lr1EDL3XfwDE4ETH1Q/9hPtMe+UJ5RaBaSXgfd615y2eStn7m
XWUXo2hFA95YbQapNa50BIaX1QqV8GJKO40uaFUJmIB3i5dwX64CETjAuM5j/fQNeQAGSzwk+6Iz
qFsklUIBMG2txMW7ecQi5BZ9SnPIYnVkf9gdCSbgjePtz6AwSA4vDPIysVKD716/c/OwhfHaFxBi
PhBHhp1hXY6N0ALztnty/QjngBU0Uq/QWf+tGJwGSFiW9Acv/ZqZwnDHXmN8iDKJzgMroM6yhJ+1
S7WLhSjUEAYavVpS8aorXwELAjLSQGub7XW72QzN+a14GIF3DjmjOHXeJULlYITp6dlxLVgEI8+V
t8ho9qqVq1mDxo5q70V3bjK7o8npCeQTKUGTDbPdlNE8eY+Z1tit2zHKTyoomy1muNM3iE2xEt2G
oqt0mBOwpDcSykFhC6WTlitJ3VDigiNT8xPsAmpIlufAXt+1Glw1TuWxp3EUTLRMO3ftidPph/a8
uyB7YAMuyd14WO/uyqsoOkmZ6ti2m3dnrETpkNpU14GT7w3e3Q2h2tk9847MupCflmuVyrlHIfeA
PsabLeD2GjvvjJz6n17+YkoCw4xIB6QHs3RMEwn21UoH7ZkJZ5xqDz8T8V4Doa1HYMvVJOUBSAUy
YG+dUkkdwhKSZnnzs5kp83Z0F1At6pa3afTe/KUICtC7dN/hEi4rqfFeU39RN5ZXmME2fA1j/sik
iSg51hu6dO4IwU+iDdpY/Qqaoc1X+jJETXXqDs7lyBBhClvKQMlgUR5D20E+GYn6zmAPVTcji9XS
jv/Yyh+8wfRTe/9Tl8Wh7FutKGYktvXtZQzUnlLq27K8HHgB4PM8p6NfPEyHJikKDUD3WcSpQ59J
+sEvIyP8Rytjo+TK8R6PfgftJ4YnUzVk9orfD3KtAbRtoVSh/NASbFFK/TARiOjp9W4i6QMenli5
AyTrwoJpOuDeu34cVKxAYp6437A7lwlytJq0/O37pBrfxKdhqkli1FPRtWgLVPcQVIYjImw7x0mc
rfVVrW4ubDOGERlKzK5ABLgVJzPoTob/YThHvcC2efii2NqqaY9E1Zcn5+Sh+plKhwjRL29eYEfG
CGFIx8AqIUI+IAdiY40bE4RNH3J0VV87H3nsaVL4XmKGQ5vCgudDWlJVCMJLjgdlSj7HqKN2d7Zc
WJkJztMHnyG+RTNG5yUW//izJFIp1uqKBotgD48BVwr14oZJhiDnrO/kI/hfOxsmeQWu3vIiIGg1
PQIcfHtn7mcZmxZwpYZwDH5NSmqgR7ulf+jxyGbSrOiJteKQcE3sEhWKsGdrrD2S0x88ly0VGwsj
vYqOX0IuOmfOc5lTdQWgMrlDiNfzGQw3y3Qnt9Zfk5bW1cd/HjQg3BsD1g2QXAsZhYTPPIjqfAGv
uqthw9nNcZiM+J96k3D0Zbzv/zhRLBeomEhUVQGNwqfonb8OOmnDeA7ebo9mJJJvwGte4GE0/Z8J
fDYUuECfeDkOMgJp+zSvwWPbYWUBmcPR40eSYjKskFqcUgmeG24LhPVhwcYySskBQv94iP1NlapS
FiPUtlkajQDtkbYGdLpZGa7CesHtx13K38iEV2ANoNiFrlTH8sIksNXWJsCoxFJZnwxrsgMSSovF
igNGGXPYk75h7ZC7vLwjHlfuvjwG6/vOBPwspopEyVN2U4gs/fRBVplKy7vd9SgQlV9sLdr3cfRn
zWfwmNCoO3DQmNDIkPeKqYHYmbVEjczReJDpVafLrkaR0uN3Ycvt4b6lmnLR0x4l2fqt2wdbctaJ
Giwgh9KWtxblJyzB2ZZZNKt9F+Bqr81UN/5Te0A/GXUgHcxkHhvYmQcVNltpDfrXcpDIXUIfVJkp
QAeS1/A/gzGidu9ooA+nY0VV62X53pW4GTNv4m9tXCBJRAAG6as59UvW0QNhDqqdyhuZ+xySLioD
+NaQI9BaVc9GBb+GnFkCAX74+Tn/yf+1fWmjlWz+qEqSPvivAKv53TywklQuVJdSdDOH6Jj3vF9b
O8rn4FRfeBjYFEI9+0Wwqe91FQJsOuL654B+g/wEl7/ahd8OGv62dHS5hnfA5xUEMfRT1cs8PFOh
dsTAfuHXq/ZxeduqstnVl8sDSy3thf1E6eqdsAUMLYYUFdyxZGK00+2np9NbiXitrnVzw4uSxsp4
OIO+r+oxPm7rMh3e7h2cZUUPcxNHgfcj0kk25qPR8h36Jy37C3S5wDp8NBZuDxPoEXaO3nam7uBn
Skc0GgQT3V8ovgeNlqud7uaGrV6U8UfbKuhCOrqVmrzVPYtolvnGitlPOmjznFwOWAIN3Hh25Q/0
KkKzw/p9OSYZMBPAGJ+ULYTtUJkl7EJPN8SpERU/8dmOVcKaqIfzu0Vq+xzJKXRQGxg+s8W53h7+
E8K52tBFd43RlzNKNEPzpJf6ic0R3yzCaP1GFP2/wXuEN5cYX+mWy6v1WWJYbxZF6LFoNBI0mgKl
QrMvasJ7aneDbsgIBqAG4j6Q1SCEWuz7AXYOqna35vP91hTwTQR1dSubJi1w6tugtBDr7OWxV3ya
h/ClHWtcUeYZdM1LtyUQc87UMQLgj30l8SgGWFIg+PqG4YZuNXTNK+tAsWaTnNp2Z6yTUEOla78U
DkMWgcWrGqk/LLbv7z2k61OZgqB3TDgqXJvm3HwhHoGG0duUKaan1v2C1dLFsWpAR18gj5j+27go
+4qyN72+QG0mgC/wAk6JouPlKZAr3k4lyEnd6bq+yqSmVaITxcGMZeULghgMiWCgP0od7u+8anzh
WTVVoT8VC15llFkauL3i7mV/wd7L3yO/HeW0LvB8abDL4Fcqo0TitR6DdAC30iMVD9S3tQ9wgG3j
oVxSOPhwnm6YlP2S/VenLyyXuwwpjyATSfIqiija/8gs3SPjPv9qMplt6buIRIrUBnUxeZMvtoha
nRGa+fNQrnRahj56jQaujZD4OWC1XaL5ZGdtfjF0EcSpE3y5409/7Vhf2x/FHq5QIVOWiM6trAPh
ppGFqx3Kn1u3tSeBC4pwQL+dpsFrhBc/i6te9jkG9cv7Dx7KWy4nCijrAShuc2qr7VBVChlOn/Gi
t66VUZg2Z7ZsHAYT9vWb7uz94pUj5C0I/TR7R+yE2tuUgsAwkNfu8efzzq5gCtgdB6JruqIn4+gY
asv7SMCiUiNBkQ32e1NIyNf9dz/OHcqnwaQqz62ZM7H1GSR7ttnJ5ptRvrPzbxhRyrDEkEY5tfoZ
SUSoz7wPcd6HgicLeJvLiW/0Tn80kjCg4dphbmDF6iwHdP/H1uCXBA4zV3qEM4yu5d0i4PsRXEOz
afvNLfg/pU2VYN/4s5WSn++uX4jjeJ1DCxLShXXK+JawWoBSBhnvgaRz6OnfNsCe4B1aAn2S2jvl
zCyo2qLopGMngPJOweT3t6z7Hize7PuQlC75LptzRSD0o7OxLKeekyQZyIJ/iFStooEwmxq5NnRZ
SAOiJJky3xWimTIjnEn9+SRYGx9sy0fABux+Ocg1MAM5XHJEJDVC41ndlvAg1zgeiAe2IgCPkIjz
WF7b+OwEqp06c/I8WfP9Hz8cJAhiqqFMibhG/9ihuNBY8LLxFPJj+Av8HjARldDyLgHmMnRv0Zjg
V8jJNH0jQQmByPY5pQhpvrgHCCDauZo6mVa5aAihieyPM1hB18CqNzeg2pcsCT9iktt+ycq2cNfq
ne0/c3VaK3vQD9znBQ+M0nVUlMBjGzO4rWC2ZOSrydz515rid0d8r7o5wlVOBe22a+ESeZado40i
dDHmOS54hGBcYFDUBJ0UtOq4hiPAMKjghdAXz7PvAMryzVigOy1o0ZERPBiLuSTDpHdsp2cZvdIJ
uU+hT1FyeTXj8JfZ9CfHyF+T4LeaSKsEaOvtqoLdgrR0c6kHyxvMX3NlRTzLSi4HeeNI9vERMFT9
GgUKa4OSeNBKw4i15nOONFYkMkY3GSCfsP8CHg4HKTMMeHoabxyP9EWJQEw7VCcr3+Z+klSLw1r/
dgTJZBSAXRiCcMGuEdLpTSytG7dTffikwn7N+5up0bOVx0dJKK/9e3PumuSPFtZT/ajX81WPRxlu
KNkpbpRYn58+pEMtqSDmV8i10g6JFvFsczXwfbALkcg/6UnGh2X4MtIKbEKYiKXov/N79WGMEtPK
Y2suTdsKzsg7HEkZr7SI1Dtjvv4gwP9SELIkHOvlMjO/j92Enuy0jxyWOSCyv1UZ1iAtdI5FjYuA
/0ENmJ563bbntc07oS1/RuLF/eqc3/griq3zKnBEov0VrXYkeOt/OVOjtkLUSNYM8X8mm+etr90X
PGCxlyxUW8KYtxfk0ZjKi/jYXoxNASRXYqq5ySYCl0j4zCNqLiGc2SuxFkq1OJXqNiXtGUGkvxBM
K9S0YQkBg3KcfP6wp0I3DHNH5/U8YxlmIjJ7hPk4bno2ItPbe9KWOrldJF3cj5XmlPp/+yHfVcSo
QL6jR2awiMpHpZH5EfeEdf3aoR6OTjV2QZF4LMaNclQTS+tl+VFC4yd2DInkpAz902WclCBO0W1w
S3XIJVIMRjeUbmreHPlSluUei2as9CJQDzTppTbU0ZSYINw7OSwDF5fAw8d308U4wHco0UuoHcju
3Lekiu8S8uimEkFBDwkftqGjLdg8DPViRK3z8VoWEt5vUA2Vo30NhyT4mIZjSJX0cbqBqwajBQ6m
I251tSvR2NLIl+lCUbT+6nTwhPgI/vmgPQgXjFx9gsnne7lPGo2AH2GqBUa+gxV0JN3lVxyVdaLy
qL00u5X4K7/sZE++hJ5auZfDJsvq887bTSAzeVc97vAEdXEcLbvL0lRCEwt6DRi6negKiYcgl9xY
VOwL7iKHAjSNSttOnVe/8hLHP2Qy0taMragd/0wNMPempJ2njPKspDkak8aKcDm2pYR/6vQJDVTa
2p61NVuhlWJJzfHQs9k9Moolo2I4C95HiiLsj/fnfRC9byCVYzZi+CGr9Y/GQF0zEedjwOdNe3Q3
Cr5SBNleLonunVp6PP4t28IYlNFBgfxUApbApTaVVnP5lmo5GGqFsRlsicJ7CVLFWhDJfTLQNEbL
oze2xJvj0UbFKYEHWQFOxkYTSqe/8s/y2a5EtyQuCCkOMAS4cS+ox+wizmApNkffMh4iZFvwd8gs
8FzhY/uaTmHXcg0gAUviWn9sx5CW1MFUgzbPfqtaYa22i/pNYpCmeCdixUEf2VpWXu1rZqhwrKL0
k5jxoej/LWS1B/NKYEIqSkgs9lMYoIIGBeenKrmKUsjRUbghqLemlwYLRBlPbkE0xOrlvUNx2FCT
HtqpiOOwCHuW+1XKw9Qs28OMA8Nkc2LyhoLkMhzQq2/gN8+sDy7Mx0FSnR1gATQ6CYR4IfKk1JUe
rqkQfRWOKSh9qr/5VyrAo9tDPrqlqoZ3EmTxtbFq80G6cIHSIphBYdGvRhamKdE+M8NWBTGU2Q6R
Z/1V+cQ2Y1qe/fC9Y5h5VGryBvK0Iz+rif+74AK6EkJsgaS3guFYYAdaNKug5BOEY3h5Ky25uYg9
/5OEG5QmgURgTEK7k098rsRz115er0qtTJeMyOzzYf8le/H/LQm4+6VLK1srX3rE7DyPEnwWmlwl
86bGjMsvHfjj9bHHyLKR6OQmDvqHYxgl2Xpp8CZGMvTfMVv5YLNthJuWn8AcKOGwqxfUNZwwvj25
7jnGhB56LekYKR+xHyiA1ghR2HDfr3nJghaq5LIoWwYmgIzVgvdetNN7/R1/T61hOIQYP9z6/ND3
sJ43OAz41+sSeQiNMdm8I+Vjs79vwvbojb7OBRn/fVcAAuLnn6XlBkkKJ0onZ+VTDfNxLeENLnHS
02M45cZcsln6hH0VTxdvJW5Z1joh/Ny/PWnLPgzVcbn1HthB3FIc4UioAPOOu9hYPiHUtIzGuMXe
rwUt1nxnwS6XHVEIii2NGlLnV+8NHKvfeZcQMuCNJeiZkmxZXmgcrWCpr3kG/crEJGmL7DLsEWu0
Ph0QCvQkzOPUd7c1We2HxzGT9ZIiXjrrf7V9WuovsiLudbAi8Aq5u9CEEk42U/JekMe3HlvLfHZX
rEKwxlb7gumHyloY7774JeKfMWAxydKlhlY92AAqd+Nvo5DCVBB/qO4BoRZtIjX6sRH6rjdo4cRt
lnuz571V5a40Ssan5gbMuzHKq8rIXft+xG+3Djem7s847kRyebpKq/Q27FpkkHxtjf91y0xtDhrD
641VrB5rr8Ol5eNHBXtpdAphaDmUkVJwlam31xbaXZ25pj0GgWzoERW8thcoNXFVq2ogNq0Ft2SB
afY+AHdNcIHrWXops4/tGaXgPW9PRUl+USATkPaZyYx5G4EuSeerMXO2Ioc5wkMR9KpG8w4QmbLc
RIa4NRlj/N4NF20pujB1T8twMzbuz1QireWySEzsBtvxGVomFEQdmXsCE1fp24V5YAEKbi/vBnUZ
tPfxge9wP7DP0xqDsuZ6PiV/dXYV1fjBA+1d5yfnVp+dLyVWTMtrtQnrVwUG1NfoP5hfkIaUlg8J
nF1M5cbn2tlukwpffsgq4LWpqycQwEQ9hXKZB7NGXZyDsC0iPsqqw09yjeNDeIHtnV0BOJQP/l4F
CLHBP4rOtliqJe2kOw76CxC2mLNVPdaROSW0Y6gfx56DDek4P4Hh5fMYieBdC6pcOAq8FfZFC/F2
m07pjejSbsIPlS8dR88B2DPPKdTQm0aGK4neD/8jZGSdVAVX2WCOeLOwCLDyJSh7NErOCocO65k2
HjOIxkfga8FK3Dy9D54VYC63HsP4g4euMW5QS1OC5UdMJcB+Glr/OkigGz2ODXjkU7F9N5wgyBAY
S5rUcVaBsX5OejqgqTdZS8k9QR1KF/rlbYAIxMk6bOPuhrUSWUZPFqf9LoB5Mbg+/JJwAJRmplv0
bC819Sp9MwcKr237rnRJv0nwTrkw6bdTvtiIBmoo3DcUXU6bH1JQgm2slkDbin33zT/DnzvOK600
hT2sgmSSdIymP1LrfB9NNCofe1hJIeGoFjEuD9615QZRvffzZoXkSbuyDmYS6i0JTl4xZ+q7/cVD
6CACagiFh0Tawtzmwl56L3gi8BLKJA+soIMkjXc+adn1kkTS+UKHNBBDxCzUGI4/gs5H4Ru56vdx
mqgr58NAlQOgKMzUHojkFaHBDTc9OaCcTaFVxFUvGISzWiQQc2K/GwZHoHPfGNXk56A5cNeesJJl
vjtaZBf7F6i15FLs15l2OIOj6iRyC7eMN78E0IxRoVeQ5SQh6cVa3/Z5MxxA/bwd4GmQV3Lwu3bO
I0TQtbbdfvO2LQRJYI2XK+A5xHBxMWGDqBfcVLfIQLfCXzyT26FeOxALXueW4IMJ8oEFWnhZZnEK
RJ8DvODDymJOCaAl0t0pDAakWyljNqOBKX2MabGsjLoN8sawAneUNwy1Qm/btICtbOykhSFeTnze
8fSHObygoS2kWBr8I3Om2miAdMH27TpvrI36FZniPmcGBskw3RQi7EGdpq8OG0V+qySaER63pL6J
BcU3cf/U9bJpHYkvS9WiaoGqVrnSnCKZCofd+Axv9J+OtvF0Szim3d7idfH4HGuv/BFnPr/RH8cE
OI9Yyw6bMd5xT5Uk90qCnZTG6pn4cuV+ZX+b3aNks310tJL6S2ixhPcIv+N1pY6aoP6vTnrjqIMx
symTAI6CyKTv9YXEUx7Fw8yAbFJuOHbvH+BkeVtfacQW/JGgB0xCkwkLhfoGRO0WB/0Q+SSQYfr/
vVojD8t+TFigZSJI4PvPPJ0Qwx297FdVxzyBYrx9xu1lZFoup0U3GEX17g1CfDD+Yj6aWwRv3MeE
IvKNNUh1jybsBuymirX7JMx9TDe8dLcC1occhuw9A3IEgZSumf9VZcQ4NaoPdgL7CR0aoDV6ayRa
1ixhGncaRGqEZp0uFxWzbLVqZj+GkKReZFY1IQeyNhp0R7+/maLLioPm8YYwShe7/dpyfMLNndLq
BHRUlw0qP/fBTD56K5DBXoYBEy+RLar4O69tlTsc4tQ0eDUHVQzebPYN3utjra75JhHCyBJwr/Pz
L3GpgcHhzUyvEAnaZocyw8m5AdhVF2WNIP0HhCHsPHsa4Na/gvPhXQSD+Us/op6ZH7GwY1UpkBc8
dmjwL1dzyxMWxOEwfheVqMUtxT36P8RYxTH8mRsqxAcfCFensA4Qi1kyGeMtiCu26jXTZ8Kpa2xs
/JRfYGscEKZ+cdZfaIWWEms1e1zFuMBYCxMUPv/wyudipwsPyr/UVKLjIESjdYgLfL6oUtnNMRaP
AipMUrnf9vnyhEwj1Xyfc8Kug3LBXJ7Gw/iGEFJOeZXgUT+lSVc06rd2k/1Y5dpc8CSoZTpZVLMU
LJtJZi78ANydKOM78edAA6zUmMHRQYa6GVUDe7GORHOr+qzHQnm+LqA7O5B0nc6bU8wOZBH1pru/
4quZZKsZwzu+CBF1FSsLz1q0FpUEpL1+zrGrFNr64UPyXRcezOKOa5GqsyNdIeVJ+zzY6LzLqV/f
2wiM6TYxNGOG4O0XvJlSCVU+imDlVlHO64lZzTuMEbYnCwz8pGUVFmuP58UE2Lr+9EaivNLib6JH
BFCXIlZ/3NuBGZWvRY8D8YuQbgXfUX8nOygYYIDfdgjCQp1WLAQfrrecj39T+z4RrQG1c1MUa1lm
JAQmBkrOcl2GJQOZ3T4lTDxmAPyP6SdDBTwndJKveqxVB+kj2UGjPxOji7/BPaVP7KN6reBz0CTU
Z1l4vU/YB2Y05YR8UuNzh1QK3YVKy2GYNpiUtry8euSoz7oYlMhBPlQ0o9RT+s1m6BNLL80gjVrY
A5HFQ8g+LqIbp01SjXX0acm3haGKOR5i8vbAJYKDs+UTDRF44bVMYYp5IQ3RFUuRgumxEU9vykkd
10OdApol56O88RI5ad1Nj0RcMZy/f/efqoVfU1GI3AGlnSc7X8Fq43qvzvcxeeImEcKEmbDVsqjz
OUDvRz1fkyUtlTUyaC/mbn5JAUnCqUg+WvH/TvDGnB+EN/AolcAcT+Q2siBoGmLiM7I98E8iVwpu
QVv7ITzZAqmnECN/8sYw7By+OcuZTC7zC//KVbodZgIZURSyTny20gIH+pKWDScPdsab4ttjZUeU
/YwsrwA4Li8/S5y91m/AGqh6DMPfTSuNS3H0DdPK4pcvwA2cWmplSoXnqeAPxqvTqZ9QUd6n/xuN
lIgbE0IxVP/nBjVmbOpq9v0oRW4mcVLj/iZR4ctOp+4pwR+AQKNqLOdvsh22GeH/TWJoxYeZJzjF
1y76UOgpoOXGJFfyamHqmtACl5bmqYznrzfOPcW/H1TpbEDuOZLsgHk+B+UO8zijLI+7iE9ykIth
/laWBd36ePi6nQQCU+bYiDJAZ+XR9IVRd5ziSfRwSGzqWGKHL8wa+x17EFOT+R21jUTtVkCWnt1K
gA4YvyAClDmqNFtYIw3Q7k/acDfat+QkmCiQo2pB/B0EjQXlmR/n7wm989EZGltGcQZ1/otpGCNW
tB3FYEiZMyPdZuHTDqPNQpD3pGbTbCQYvEr8mk9Y7qVPpVjFUuGXKwYnH9+ZqBsQgoS0Gb7JlMxl
jzDEnWEvoanI5vxft/Ic6F2gG12vMMSMfipxhD42n+F3KgX//CmjWxbXqzumHMP74oufvIwCkJy7
NkcIdcQI5pnvPmuXsjQfqL5gH/l2Q3bQr1AWoi0Mynj7cRruXwCsyE0PeID6Fdj1YRAbk4mkew+8
cZ+oQOQm/nR76gWYjCxy7d/tLWxsbvAiaiwohPkiA3yfzGkFVcg97si+mBm5C3dl+yZydatm3ixe
/qFc8EhB2yMjYsT/hJ0OfaK7xFLzVHTeqb7sHGFfYuYJJbYCcXEYrH5jicdpsf/dnOWa0VA/zFIU
p9pHCd376YaCCmelIHZtDGp5U3G2v6cFRRCSQmrGK0s2cQo0fpnFI+ZP9hTggqCtS+e1JJaWxf38
q0A3CVfdhJ/R41oDwth3bPrhQ8vCP+okW1xTmXAm0t8TA2/lsEHPx0DJ8bsovkesAdAbmp+Y8s10
pcZ8nPlSikMftLNd0H4+fRQpH10wKasXRYvBIOioHyRQO7NINZKJyuxVPHyfSrJLXj+pWqSp7Ldz
8Fs7qJgPKP0KfGDEy0cnCiQdObQakQ23K79dl0DM5LUohSsbGMUE19SnDHFJJ0fqSE80jkiSx+Au
1j/RxNXa+dGPcjNXTQvAVxwozeXSTSU6GG2oBqf+urwD8anYRrwR0nyb0tdaXPQ06RQUmcl+fn9w
Cz65/n+he3qzpqLNC5PfczynQJupPMA4minrorl54DUooVjyTZeWcfc2fGTW4awo/atj+3pLvML7
TNrevhRc1K01/b367vSWGrqooP84cBYzdvlKTymiIgAxWFfV4vHWyYccj4ouw6bJ58+oIjn3iNK6
hEIdCyWYSw880DyW3f3fDTe9Fzy4koRIPYier9nWzZ7QT0N/EZ1Lm+PzJP1RFHraNuxiRxkBYXRm
gQiTkwNWhxVPCUfcVxShKxNEApcVT00ROPyfLHMdNfJasdQcqYifldtFGGTkLPajfd9DXsQZNnJW
7w1cnN5zy9s4AOs0HzTOpzKn/ZeU0Yjrc+NV6hX/tvpPR/+70SeHpkEF0K5bOl0QcGrU6NALHpgv
9LnXyjqM+46yhvYfa9Kqrz4R68cqHADZD2fLI42za4FaMRqdgF+2gx0OUkX6NiEOUYLkA1i1WuKE
n/wwlpk1b2cRatWIcrd9tDNLFP4Nk+bN6oh3TACP0NpOm7mgi4HeHo7pt6FnRZfQZwjJMkz4kbTX
KaxQOq/OwW7Qb7yyCyIU+rt/XoPppTg/BuMnGHUz+nNCMi+dBvgfPD2kzbuiVwfFf92c0qDabOJu
7NhSHlUg76jgN4m9XeYL9mlIDD6V1m5asDc0xCq61r2a5CmkaauuGnWpDe6cTutNOlzTWA6jvROV
9Si/wAvLtodXa95vkA7a9NRs12XPLz1mJDPjKq+G6plCXjcdVKHDkjt4CY5SP8vsBnMm/xndCeKt
UvKQjPYFDFyLTN3mKI3won1Bp43CEypyyJHduOQcCMliAF6D0wD4EiOuHgHK4tgQYLV11GsQotLq
KypRC/pzCJrAYmo5nymMmiJO0i7SphSKeNZkl2yt1fwAQkeiOCQY2+7sqvUE7m057djGS+9NGw6j
DyWhR+ovavg8nmGf3pYO0oop0R7b5wFZwwFU34Z+TCy3ECR++W+bdp+4QEQKXvD1VXu2PT6Nt3Fw
yCCBthOWd7OmPnOMW+2EJFqLrIYPrdJqIMlV6NdbohEBFEUi7o3pyAS7QrKTXl6XnSWJOoB/PaZG
SAFJP9jFH2UyibqiMIS0ru2bK4dHPiOg/tOT7d9Pxj8yEcm3M758Xg1RC0CCUo0ITy/sbk0TK4MF
bciN1gSZ4Wz/Dq0Mowqiei8VftWjLqRpqJMwPectL2gA6Knuy2yZWZ1rsJfZNHDM+MEHfDbQt7OE
Kvy61UrCNaoWcyEH3gSnafzpQsv/JM7vmHOJTsR0WNqoe0uChaKYkufKt+nbqsF+9S3u69ZmSjHN
cujYQG0wZtGiUAxILDN1CvANz6QhdwYge9s5hz78HMsbDHL5dL7Q4u3/oi+7a6CeAIdl+Y/DRi9p
t7X7hFHSPpsp1PR2AyBJYAcH9vb25gBQBDUAgVUYz37TGZ23fI0UAsOXMieq4xZSKylTjCme+QWQ
bk/4bXRgqVmTvwnzULmWiWbW3sNmiFd9dVc63qW3NVnxLEXkccZ8Mfh4z1r0VkU3ezv8WBRek1o9
1j89ak9CbUU6Fu+TRgGVNawTiYx178ymuPU4quRHUginECUF8Vi1Umb4WDn3l5dQvHp4VuFrrNfS
5frAvdbf3FHBeVKUSG0EB3A1e+SzXZby3/413GlowiDolaR1dTlP9ozD/cR5IDaonxurkCwhltJ+
SQYgf8ouvtEmgkVVh6QHC9jUy/JfXYdzisv0UBDPhD6teBS70JAWQL3ZlWP7cLxa0Bv5OEofZBxs
poutslZ+I2INUGt3OVFlXSMyZyWaE/qKhchn4QswUR+j646SQ8rR1MCd2w5HJUSu74dMjougFZky
xrauLSJHOTUavxpDtOv/W7i6AdczK/DnmBMcAZZS0gFTfktXrTphX2ejJMVfqNome4RfAAGUUswl
pTJbz613ird4anBFzAzBNtrCtUtC9K1pZIzTTMlo7IwoO+nIuXZhCEqKXxvH5iuFww6cS/qCcyuh
wydHEk0aweH3OYoUTz/efjQKsGHZ1yEYdJ19RQ4at0e9JtEuStYToUdeQlFIg3+183C41HN/97Cw
OV2GiwjLyEFQ69KMjmU9C0J5qsSHoUS8BBFIfQF3/xO/5myimPa/ETkyafKpqhazuvelnoq0mCzX
I3zefT9eHbP7837Rqg1PtoS2Wzp7uVClta+lhfgrlKGVSaL4VIy9/WJgmFLm+GQixo1q9LWZooa3
rdIcV0rmVjge4/7+H/h+WW1HADFU5lkreYTeJxAjhVGHPqUuoBldCtZ5AKtVB6+G4XwcWrxA0zn1
xxZyxWk+y35IqMU4P6yshpKdgOCq2xLLEvNO2YPL88HRiHORMI0DlmTfYIVUo05kMXb5Moxi9GXs
eFGSWZp61bACV6fgvkQ5wUjF8Mk/OaWWIkIK9zLp/5+vh3mBAfuBed5QQFkXfYsB8NlCJxRpbcRo
G+qK+UWsXNx1vEG3BpBmEvaF22gQxHwkbTUXI2iddTAbUt8+8cylYKc5tOIfTY+zumHCzw95XbGr
2yenLzB7kIkuFPofAoFkOVHXKvpODe/8TxxorHIytZDrSiyLBuic1otZ7NjNECuHeSnFR9S9U9Gh
o1DatXwoOm/POemcaJ3CGSsm4dLKjhzF2JjgrcVWVsF8yxSnourY/vMcP7hvEnLCx89qb/bOl+KB
DTtEGUHHMOch6qejsVn2aUnnFNAWuZhXwMa9TXU2Puh3jBYFVTsVwT/Jsjjx9S94SGniDeNIwDOr
nzPd0Z5z7K5fr0UYZHckbQX0rO04ezu2NHDt+DDKcGrCtQL/J9P2pHBJFDGNrRm0riW9GDWKOjd7
N8d4a4nX5LlWQqYOnvuoih55Ud5niDj4hJKBSD+6DJMs4NQLMNEUUeA+oZbFUxEhB9hJi4ToEurq
29513fTxGMw8rcd9Is1OLwiTl/UaACbvLDqVB2LjE5YNgaD2GindnlKXI8UJqNTK8YYx40GElrZC
d7rdypVnCyC8RfHBxXtOI06AJOkAY/HYZvwukeUE+YdqMYATUsutsvu4J+qvwNNve4h4JxFAJ+ta
tYAqwmg2xLXzzek3xGwFr7dvQcUiuOR/Dkh0U5WJiwwRnCao4LXNBEgy/KCGzSD05tIXd0Zo3OVG
ixMReFrWQfciu7ZGeplzrh7qQ0sPOsdNDJjIu2EFq54/9c62Y4rtJNCcrQM8aVDEsI81YYCFQ0Md
UbCrqjc0YYZ6/+9Lm/nBrWlc+34q+XyNaz4gXEHXyd2bGBTV7OVRofFIYSpmWNsaRd8Lh5Py3YZG
u7KPhXx6F3HPYXGMSCoKod4leVTqtoIZQFZ+EgkxvMwJgIrra40CY9Rjx6B51h/2qu7ADoc26EV5
v5uAXHsSfyGoShDxEZKdF7GVL9ViTb1O3SF55zu5i4G4USTXX7ea8N1uC7kBu3W3lHtk+xMOzT+U
asfqpQkByK2dcUqvsz0Xri8NhjB2r97s651fGehTvcOHsASIXzkB6umE8NA2Fwh1RKvPM6U3wX9t
v05ZtZEhQuh4E0v+4nJp9kr7CsGK5vlFjmBQ/GSFjwF44Fznp+4Vyas9U4gGZNfCcCRzaKOY+zb8
z5A7Gl9lodVxNGZJr0onRgwa+YF67G35QSFS4+BOAMyOvfHgXmeXq0ZggciOAJjSbRMcmQUNKDkX
CikQv2OBXAW+H/Mkn03pGr3zQCAhPz6x7CbVIZqeMD/dWO6YR+sYD/Wqk/2xxi9E0wVtZ83gwmys
7ux3LG2o30Cu7/tXbAirICpwdnK49UF9YWfRiGS/5RtdWx1bKO7661GjI3U7WejVjG0qdEQCyecY
r/DcYpQxwSUPXW/EqvQCOxxXAdRpCe8gMQ3LRiRCkeVjfjNmdc7uRXs8YMKHB9rjmd1dXDpGa4Ep
IdXLMzRAXTksc7F00T5/PYKGSkF+8mCv88Td5qV9Cfi+Y1BrH/U6qgXgbFwt7L1nVQOXBXLYUS2G
bc3DlRc/tMbI+TRnrrVWKoFXLctSwO2z4lcRhDaJalofuI3l/UwO3YhNvJAFoo1amUUD+IDZwDLI
BUPdSrtAvgYDv2yYksqobnSgtCx0OW8tQrE3CL3T9yNO+ADsiI4A9cizojSssMV3XdBpgT/Se0/U
PPA2QnSr+H+A8ngRQdlsG+mHeswKU4ovk4bY/BDyXyktSPx52fOOZTQ/Qj6PwYYwDuNTRibi9NSU
k/D3i0jaumjHdvtSVSKghdVJGgnp/j2QOQKtFso6y1laqZ4fjOHJpken2QJ3QJLJ6dHXfxkOUYE+
h0PZ/nq+UufpLXuey3I422z2pp9Pk57H8KC5r1M17PHjqeP1P3+HSWzRudrl28ZQ4+SiGhtbWd5J
mR1q1mJyDU7zWCbKEdl8NxGiF3frSXr5qUn1hzQKXIjsQv+dYqeI98hkpL70syKNI4/shZtuFWks
gk4t9XG5HdmQuIV7Au0oWzrJbNgU+c1A6EcSCNgCUQOvWExdn8QcKutGIJWRN0CRkwf4tzWWxqCd
To+k1ZdTXaYWYkYdJ0naIE+eIpaMhsQBmsEQryfsCAqSF8AHAFcBekG2WXpfSU7/vJpOqIAEJAxw
wWdE3u1TeNvAh2cFkX/recltwuLA4Ms1OSkeQ9iaMbAasOHxKZtSKDxq1fTSb6OGIfyEfVUXR84b
SESz9en2Sn2AvPczqVgTo/q+YjFGiKRh+9Ep37P1nBcF0m2Zu7iagewlj4ez+o0QhqlcKVz4EeNl
fnX0Cp9Gan4KWJaullQQbC2xBq9wyqZqBFGE5AO/rjCNR0y1/jvabAtyTECWps3xKwQKp3qOUPxG
/9Arm2gZcyk27ZIos/qI6NiLOmHjAYTeFdbwFvNJhNLy93UwovXUDbyX125J3pMy3eOrewFOLTH6
x7zpDndLxbFTSaHrAJAOClEe6VrYswrQAGA/EgpoxYYcdM9LykovhqCXWaZdB3Qr7MLxtjn6gbNY
j/rBCDcTm4PTvfefVAn6YrAh+dfqc6L0L9gzEveTJzW4mBSuhvIy4eGUZqWdXJ9FrzYfOZkDAzcR
NIYo479OQhFX9HDXZHrkzwq9V0egjRzHIasoCBv0KTJPg3rYMfGbWMFp+2JYKkjDNHqO1qzItWzc
TpyfLXXq7+pIYri6h4/cRkEk1H+mJHz/gXwCpTnrdrlmqeJuxik/ONMvhoG9l31AtWNuPU4CDUOD
qR4wdJ391k9TLRXyEzkIk8mH2yGQp+bu9mqFwSsHn7Dp55Q2zpT6v5QDDlnXvJdkIBbZqSNmwfyb
ZAHjzV+pekhnoonabKzR/FvUrZrSnUCdXioaddfyp5+lF480aJYI4OexAjhV5cQdw4jlE2Ermghx
86WAJ+fJYV4ndKK2QTHL9mZuDvf4lnCl4kKXMLQHjKsjXx0h1aP3uhkLNUTTI7ADwFEyhAhqbEmr
WQu/fCF6wTggXa9TiJ0oacQKYhLQ1piSUT8hfirxAuyQyG1r6Is0qqQH6CcLmy0kCB1kDUD+43PV
Dg4XC/V5wONqZ27uwQt9tA8LzG4bjou8KCaCasapPtf/jKriXgUtC3ZqAJ4P7Wl/GX3hLjYhI1PQ
QNn6awI0dpG72jmMRn+LI63/+KA6Firl7rVldrJo9Rz2lyXT93r7s4cvXYLzU0J0hfAO+Or9MpH4
ONelg0mUm5ZKESWzvBscfUIDtcK6bI1WKq88za+zWlQLozpv8Es2irO71B3pQq8UA8HhT2xGqNpe
8SxQBdSKgbc2IrPmuzBixnLtfk1EuR90Z2cLVmrl20Embvflgegwexc8zAwz1R40h7tuZ06cNf1a
tUvbqk5j8qot/3lHogIxTZ28vab3K1kpv9kn/XIwLZpL53COnI6Yf7KfpEHdWBlD7TF5U/lkvpwl
rB9hRWmMP7KFNyfGwBZQhOQ7ohV6S0Z47mG4yFQncuCnILd3v9pALzZFOprQ/Kp+oQ8H4B0blLqI
4OBX6r2O7Dfgj3Eo+BMFCF1CamdyO4y4hzuPZxfDoVDFU5pdogzPUenmajLcghSYO5Te5b+uDXEt
tHFW1IHzsAcYqTBnvA9mvSrfMSG8Ov/MHftWJC9HubPLOpwE2Yy+vc1M+8MFTOEzMJz1YaMcFiWY
aT4OrlEyeTF+AQZ1rfrj5uSGxwZ+sJchg2zJcC4BA+s/VQY+ov7sj8OMJvtDNfUhMGH04XSde6mM
j/KPIecYXR5b3ZMMniApxRcyX91Vw6hbKI6LuwUoIb81gez3/goI8agmq9W7tiFOohBIOXZ3P7N2
1kDm2WpDUaYeic3JGpfA8fXtMsGjBtuk+36+RMm3aCOAyHvcGGGHiTCvs/xKxkLR4srgjOOdQM5x
WQx4u0YI1EKSWU2etYnVqfgfyazwSa2QfG0kff+efFKib/jp9t4YdtnbXdIhLRYyPorl/hhQllQe
eRxnk1W1HDHbxEE1LLadUNnldn7J58tP8FhyJ8OGxc9X+BywpTgNT5enJXRRuMfLREyBiXB2jYjx
lGdMuAfbyPlJzYsPLBSUMoyI8PikArYe6En3ewFgic8bnY1hDOmym6MfKMhBrrUhJ6h+w+ElwBHp
x7oVw7degL3GVUmZTgklf/TDZvzbyuDkAYzZBxdBGq+V+YgdVTk3aZIWcO85MSgH8RNjlGaUJKzS
TEplwan/ovDyekUoFjrMlbP562ckQkI4ORbl4T3HTBuhIaWp62BXBtNWfrD/yICT/5Rh7n6yrMYz
wFjbEH9RZE12yywbog4NNyoQKDm89OT2UGi69QA2OhxWby46UV/mKMUraQhEQTuevw7CK9ZOR/n6
VFF3WfTfuNUprB8jvHhl3bY4rYGpA3YEmYiHxp5LGTaBCQBWEsLq4VbYTVihg3bAq/79r63AZ1Mb
aI8nB/6zEe1ikbarVKcHBZIp+auP0NyHtcUcsdi1tTVMRfbyzhzbyhtAJL2Y9x8qH+JGiQuQXTaO
dvvJygcL/ad/gXmlptAdT/25c+A9Gl8QlCAq9z9/hHFyZB2Y0Q/SsPGbQcWFTRGydULvl6ZocdBw
QNU9GWe0c01e6Z2Ou5UQgZ5nTxilKToD7XQJMXBkJ8U8tqPTBXEzTiQEXAUnzAKrTcLrWg/t74N5
1/dEZKyMnW2i35VqDIr68ORe9ANae+k8QhyLbZn/Ft9cwoQvOXuaR8mNwwYR9h3FtozjU5bKqh+Q
1TBsq1yogtJ/kf8nt9bFSFbFBcdScNpbTQY9PgoRv5iC/QOS4n55BvWhYegm2GR0bjaOtS6vMozq
aV8b7ruu944fDNt/8wL3oHFJs26ApwhRi/DXGQd4aEJ8HGGvYblnxDAasWrlYA+0f4yVghJ+jxOx
XB1QuTsEbl177cfXQsD6cyjddh9+Nqy0wOEIRox+USSbgiWcN7odSWfWesO6c5seRY8DFdJTMovP
2lvJVBUfQLNR+X19a1eDwLMVNyCU186GMsuyoRuAUlKG+voEYkVw0887Z2K+UccKaG8zJEPL7F8M
XNkKq+eke5oiphDMXeLEKCFU3IREPtG6NYMmGW9TyAk90aDFFWGGCEJHBHSzz1lawxPEbO2TZYVx
59Gas+Qc+tgHxX90AWqExjhxiZPmtgjlUiY7N62pZCpHVGhfR/BP41hElVoHDTdt4Ejr5xxtApZV
F1igoGrUyADMs0d1LxL96M0kZS5nF9vbjRxPXSAP8r2zr6zqlviLDxeLNL9baASxXAffAOBmlblZ
FnFuDDHKlacViO/ICYf8b3WVOcjVO+Oh5bOc6KeD4jMrfN15D7U0Te32HmpEjUw/j492inZvyNiC
vkEdXvU8aVbax6/vOaPZEtmX81iF288Hy2LFoC8IE5fb4KvqvKjndOGOAUKbv+zseN1BXXG8uDzm
h7PY/kZWJ7wOiedoG/PWdY/7Tmyi6+jezZpiEcLegd6MUPVyuh5kYD/EK0/WZpOMjTy5YCTryf+B
KsV90cgyhhuG1eefHDTfDhUGLYkrsOv/Sbtf1Umjl4mkaotyzf/BPp6lnJZTcVrllUcSJPeclgOy
0BmLGuCVm2UM91o4Y8SstN7QrugCC8l2jfzuYcmiLWGEzz2908/gmffF0Ej4LinCqdLOhw6zxxC3
eHbPAZOLhO4wsH/KCpsZaPZEaakejiPyvi6+W2gXtBm4p/uF1pVkmuX1t/gmMmn5R3oCH2z7far7
0ixDksmAAPVeNHJd3rDYIjmwNJSOxpDYK5uyMkyNo80F8u6twJ7cXkNOPZymNYJeQTBYwk0rk6lV
6BVohxfqD9+6S/+uiwL0WIVXpl5wFcFZHAUxlOW3gYPXn5JMhOP+xVDmVSVlktSc8t9qXSUnIHVW
2JVW9eRMazBgFJ7Cs6DKC4hghDfFDG4AgJDzyIjgdOHnFPqKAI5lMBa34w4nRhFw5drmJfBBAW9E
5xUiKOtSUigI8OuBJejNecC/SS7RUKWLCePOj1OSfqrTqHFHqxDURukWrWoZ4kq+SzLAY0Sp+oO+
RH2kqkJ9k8+dbl4xAcZrJq/PpVPyD7fL/HCtkZYwfuLmqjpulNYXrEHl1zO7tPhO2YJgBL+U7j/v
PKj7FnVfE8zrHDgZLJporkE/syrMxW5X7Qc6A04EL1TLCi20j+wQrkV0Lso1qQAJskrisPrJ43+q
uJhEztGtYD/G3Nj2D1flJ5Yp65TiOzorphT3qK0OrA/0s9MBSpRpcywTPcsimnMI8jxkovZXVsLe
cw3qzJlnj+mXpWhpG9VA+MAoMLBGy0qgoVDuWRVoXo35SQaeNe2n05lF1A+drtkSxfnTLuLWsK55
yzBCZZJwNC2LBl4fyU4waYDhEmZos6LEEhFkWmq44JRCJfOvEc1NFe5+qPTZ+LuoZqCFHRcVlbNT
bpjrRGndShUOk9gbNL2C8B6V1Z2R4NbVb18sAGRwV2OdLJjOdUbA2WitkqK9AJR5KSX3AZyworEA
54C+8YpOlmdaqTS1zITYxS8YJsiUzUKyWeeQmT27wmRhSws1wU9ffgaKW953OGT9Tl0Hoa/S8uyQ
yRPRFTYWyZDHg8ZdgTp6/mkGGPKTchHU+TulSQ5VfSylTLBlUISs1I+gBUXLoEYZxZsHWlLG3oK2
SgxRqbHSCww4ATQsOs2u61XyEoO9hTpKhW2QuaPQFv4ffWeHvrtdmrVU+PQZ/b7o1g82CMB6Jy6G
gnRYfFDq9PE6SQ4+KnK5UD6KXW3FAt8Le8fvoLby2bIYfp7OtyOJoRypA20Jx/NM2GAB9WLSHjrl
y/KkOFc7ngZ89JzTiuhLNSOwsLRO1AgGQ0IVZrprPLxAbMovArn4LsPQ1hqkC5fGAZMq9dV9XqEl
QbHynjI5OCFnFAy6UzSOM7j6dLAPKHIHX9XjHuDNsvt/uAv4YtO76l88ru5vAJI2mfCyi3WtcZsE
Ma9KqhicZZefaN/Bm0m06i/3DQj7DQBqxFQv/MIRCoTWNGp8a82vBk4debXkwBf9/bW/X8Tr0e2/
+luRp6R4CoKswpYB0MBAB5LZAqEIHRr8kTwkAVpDyFL0JayfQBYhGA+w+0wFk0P4QCO8rYD5BP59
I02gR3A0oC9mbwTHYi6XvmHsYVPOrMouKDQAl+eSSHvvMulqCxP/AS64unfIObCgZpHsFbTF/jRA
SgdROgIGpjS26/iJi2oX7VQ661G8/9teq5mVohzA5eYAL/GrD2rW6Iw6yS7msHHmAkdgUan0l7oT
oKsgbB66sYjZRwWlbvcfrcU7RJY2GsTfKcBf8Siq/TAN/DpQtArhlUBDOtNDSGvWvTX0TPJVEOGR
QMbnMFFB3qSwbuUmQ01VhfiQX+iNzrVENgguiuihHPMA357GYsxqLpJDyOKf1FcHcPgVlcBXYJIY
mcxL8ESZTq09Zr7IKBfB/yEdBA/Es2PUAnVRikHzEsPjKbOtJChcSb8pQOd7QBf0NMAY9hbRGECR
C0sogEW0D3E/g4ORPkzCMDxLb0er5PkzV17G1ItGbm+xJfnL9EUaNGEahDhSVwJLRiohsbs/PjxF
AsRXCgFQ8nc33Nxnrb27ROVDL7bZxs61I4V+QsCxATqOtrffBICw/B7V+N3sqB9su47fEJKifpp9
d4eLxoLNYSDJpI5U2mMr7lH7sAh8ZLoSXG0G1V1XfrkjDQzHj0mMY+YL11MFnbjYiBM4hXxiNrF3
MJJxlCQU3BzCnTD2Y/7LE0L7nY2TZVGgKruPYR5S9vDtMr69vUU5swpDJ5UcbrZwySkVBWpak0xl
T1TA9N4JXkPArOsPna3D/YwtKmdX9SIdx8bWm5I+pzinXi1ixtejGLtlzqPJrNifzhM7Z0ekriNy
6OC1tuOYDItGbi3nslwjCjE6o8yyieJI3iBkK1reQg80piYbla4bhKjem32z4I/ONb3o/jo+cMum
xK7zBuC0BGB/K6zqfNG8N0cUjuZW+W5awTxsDHdmqhiNScWGcZmsmy//0nrNm6ITqLTjMs9n98Pq
yxhA8xo/xoaWvCZSEVd8Vjh4S3kyF21jOJccr/CO6lC0srPIGCiwLrPF7z5mKLwdgMCI/64oRkXO
OCRu/e6ZWPaJpGMZwkrSvXW3Wf5y5wEMgA7A0vC9pVBS2wxXmyrxf23oq89h05AxP9Y2LCgAXFsa
K70F9e1inBT0HUZbLjaIif+glLhm2Ji+2yZJeu8gCifMs4KcC1UZQhfZlud9vp1iVmQxGxqXMU+q
XAx73QoPOHGem4gcJ0xnFD9CgFx2OzDEvcIdw4J9vdTLjja8ix3pUeOSrKisEpHSHCb2bvz8gcGx
c/RrMm6WeAZyBDxRNFFImKbFI5xTqA0r9D6hn6LjJ3fgZ+IFGqBa38xim/kjFF/b2wpU++OF9aK9
EWikBYrEh1ICANErrHYTGL8X2whwa355LzJQqykqOFz3/ChdNMNBQvom39ENsM9RowgdgsPEQ5MW
N0cKuO9/ZDvmTkqVcX/N5m853ImQiWxydsZ6rO0lts07Tg52u47TitWXYah6wiLMYLOOVlD/Th3u
q3GRHR1U52WmqKcpRZYFsBBL3DYT/vl+PkrxXJqqw2fAYOsHcXIfewbnHER7dS+P0i2hHF2Wg9e1
uprJ+gFbMebhIQQVEM2tZaoaMVdFaak/XuF+MJzGadE5HkSJJsowK8vrVu9iIQoHOyv0MntVsc4V
hIZuVwAo3LpY0q1JZu/e6SOeCgJQd4Z63hK8qB0VHgjwgYLKdwGJKQuv83RWMo4iO6NHqNoBcDrM
mjfwnm7dL9mmrellCAwG76Jh18MnhpVE9ERYnbTdZL23cjexc/BvJwI8txCntY6oZkwf07HZmtp5
px1LEv1ibBx1LFxDYdcpkUY77KLrmd+e+V6lKfXIACdRjm/7THMC3vVNG72rgQ8VEMagLo+ABDJe
ZrWomi2rHVRH8P5kCcwc4IulV+E9LSihB9UVKdxg3l/pV8mZPh/IcDNb0J+njcl6jEpY9HRnV91q
GBZl87n+f0sdKGYmOUTa05y6QOFo0sT8nfpV7fP5HDVri0E33sMx4t6VhGJ5QyLxhB2IkImyOlcI
3fs0Ak8niH+0UPMNc9caTVrSEcpTWgPgNoo/lFnXcMJuzLxeD7bVj+NxGhfbswBKOnhF84ba3yvS
oK86g4mQPaAeZVxGJ4jG7wkShycYGC+3smOX+hbFM6Td7n3riMMbFtTYceBOYQEnxecyvE4QZDwH
E44g8u8JEJdHetkSFLgmqVWYE4SkS64UZLWRX7Pnn7G0u34ATTeWJbFZvWvmlcndEYEgLT58BFG3
ELrgm3nslBKTIYmkvLRPfx3BuByFRAwD6JCm6clvHLEetDm5NwYvrl08BANgn03cfK8RQVeGwhGt
rN5i/ss+f0ht0h45zd61a8C323BCrDzdRzS3M/G04VSRJmm+zIPkwCnZxKHlc/SdAm+aVRsYHP/P
8i5ELs93ZgjEPAJABjifjuDQ1HZnpVka9mdpDeF+QMiFqbY9g5lcf8cIZpRRNGEzABG0dVCtOvCy
5vusHKv0/pKNYxoeMovK/3zgsmTm7zdOcZP8qnu06eKjBTLqkNiSz/61lvUTLTa/rP+Y0jVKeDEF
fQCpXV5ZZ0iI3zYFJj5lzR9JUIeZn7SzIMa+G3NL5U1X6I/UUWMc4tsrKawYmdjI5vGQpFS4zf6B
eUDJfKga55jEYs5nxTEvx7sjepWb0B3DhAtYcR1Ahl4lW9n6i59XWwPZkQt+enAi2tJh1k2WewGV
JqfZdMSGvDpcMImN1bfpmYMcgUb7IIOLgkZiRRjPGW95EL0ENDUxJGEwmryf6Zo3n0KsZkZJV0sA
pw3gQ8+yMFneqZbHsZOXDwRfexY5nuvD+pOWJX35KRRttU9i/qQtzVPYPp27wS6Fwi3QoZEBdEH7
9BMeiJbLZ2SgMfJqJ4qXRFD65KVN7kvtd7F34BZuOnfTEPBSqIiwut9eOZIczaF9vTJ71lC+eFKO
kqoS11O8tHHJKp4v65L14rsGMzWRcreT262I5MaMPfTLWw/PQidRveBCsP5q+WR2mXZp7pY4VosP
XKU+JthK/TOFyjQIpPAl1Y0yA+jjq+xU6togOjjk7MG3RVugcvI+qRuJH5QiskLWGE4nu1CpmYTg
OXMnV33OfBotxYAk3Ou1ZQmEO7I39L+55+o+iEdMUYjADKtf66Z3ZRcvJztd64oytJEFctVO9D8n
Rzprx/DhyO4o8xlFqSrCuS1CCvkzezp790xZn+s8V6dhTC2Oys6VqKh/A2vMHJ9cnDUuqow9PruO
BTEs1WANQOXqjkuH9L3DUc2cZYCqQZExc9BWjqAflqokHDe2jnaT2Ww/tzJbCoT9RdJb51lTpXHK
+OZPuPbcq6YArbRpOBgwTxLm5IDY5cEC5tG9aF0JtFX7Wh+BzF//0KIRAcUNBXlCT39vkdhI8P5e
KSse9BwN+LOdlOEpEQjsmvPb9G8ZVaHeFNSyCneQvY12GMSlaJJTJscE6+dy6DIpRUEmbXsq1m8P
tEJw7O/4ydiXo3EGRqHRkymRj1SwKnsedzdHvg4aA+1EyCGzQs/4OAqItAhZx3H9Yr4s6GqhX0kd
jIrlvqw+wMgkrT/B6zveg7cKqosV01okHMOIdx6Xo2lGhKcZdMD2nKWQh6h04nGHAdeCK0RO0NPC
DeqhfRvxaIzLtCeznmkx8AUynO84kpvnba9/yjGoOapI/n6xQV7Ri/6hgKojnojToT/kzMl1HRZp
ghq+5S6i4sWO2yYSuofoHw9nAOViCDf83HxC+Of/2XwcxOAp19jiFxuJV39pJUkAj8e06OV/ouNm
afxBCXOAbhEdWuz/E0Q0gzc2JEmeYq7ujGzw4A8+Yw7enEEcWCSliYy3EnpKZ3mRTjKDkYsBgDRb
otw46vqhOxLqq5apbewP2QQfOoTCfCVtBX7eVRPmZS85/DiuJu+GR+FqL/RlW5ijtORGXkISZQ/T
fdNfIZ1fbvfQqfFjvCQriW5sZlD4paVNUg4if3/H05qJ06Wf0J6nyqZOVP5b9qqY0figivyJKTNg
gkZ6RLRxuraU1ftGnV4wsVkYRkwfzZ84K0WjVzqWpU6Wd0WF0NWc3XV4OSGWNqlYBcAE5xWOJAYr
2nI+rAV5cUnnsXbhlaFkNAlThK081b7s+TS+Fu1h3f7au8YeiXMQNOWUfxDnm8cHjbhGhOCvuJC+
xxmPzUhO29wzTj5sSvDSj/CFDOl51/NTnorE++OOvBvsNBBpdG7oaPbI56uqvCuL91Z+rdyF0bWi
2iwMf4dO7cu26aWSPwoLOPuh8cIOR8iSeBxNx7OQv8L++owMCXaU2vIwvz30S4UC51QBtVNObimg
4+QzjIbvjitBdSzd3vNR9C+yd6th48nNBT48fBEgg352Qzr7DHGD3ss4iFfwyKPgn3ftvcVJzx+m
OhiPJW/LjOvSbNlT6tS/gPGwsuYy/9fmEgD4L8hFPkX8eYPzsgV69/UYfwV2fL2TNymM0JHnSdbS
D74ivZTWA1yGUSENJ5Qn7FuxZ/k7L22VcVrOCJVOEIa1UaSM558ejoRvDKfBmDgrWD0cMxBpF8aq
6QLKk73GLZMzn3CTJDN/bQ31BVlywXmySSHNC+BBbk/qjtoYaGEgcwbYoCKMYtKKdcH6CDT5/K9l
eQuY9JZ+IonhgSMlGfg6VvO4gezWGS5M1JmsGRKSQeMhddBhkAW73P+oFR7M5dKlPHeTLDpT+qHW
D+7lWi+omraguffOCw/cAKsfL4boKj4J8f2MRSXJ3CNsLUUaXMIvkVSDgB9qn29OkHXTR5rxVDVK
PmeGQ2hZyTjlH3ym7Qpkc6fZwmhHpvnIm1qhmGXJKda8W+JZfOiWRcfjuBbrnqZjLMnv3fYvi6jZ
1EB/Dz2ybNmX2kRRchRamUe7JNrYGy5AsFNiGWdmzlEJb0CJcl0Bn0fmzyX5omgkFIpxBHtkebVb
oTMBppFwnw8A0QE3yxJtFJ10xLnLMMt+EvN2ZbfNM1j13MKR/RYiTO08aJXBabn1MKVLJweJFy5Y
4vUTiHYRUNXnWXruvx25fh4ZJww/KWleYOyMHh8RNLNE/38dop/nCq+MIp6htZZgi5cJCPl/LffO
s9perOalIbdMsBzmMaPmIZe2fRwFwailEBppPWQsi7cALbSHozBNo0U8yIWQrhoQa/n1IO+yjaFu
rkgMwfQQcUU0a5fWCO8eNICQzq/M0ctr7j2M909qQWhjHx1V8XW3JJ3HhiW9gZFTT512HeGOdmjh
0CfdNTMxkMnO/nmydnyW94YMxwhX2hEGfr5YdgmHQC8wVxYqkGy9TtHO0BOA217JI+QxBue0UcKI
NvN7THwklkppUZqXOa88h8BsTIt4lUTfoT4XXnCpULw2m/VYdGj7izgmlvOurg8Lj/uKJUU51PUA
XhC7wNU5blu5YUrBWCCWf9kv33WUEJny1/CNniEXKMwjLcrL0v9rCnNEVR6tr3AckqGhLMxwqLXo
+vsUr/YoawrmrojoxfeL5D187h0sFtRaOwl8hIUcgebcEsAMeWwOR62lvG/iDZADV3MVDtBfEvQ9
gyzK/RQzcL1OmnmxnY0hUB8YlvbwdXJdr7Z01cPAZ3lhUY69CDjf+LIb+wKpe6ip8wDqC/pk86Rz
3MZ/P0nEI0Gx/pZaLaNDF/IEse4epVS3llaY+D4RICAFQWG/gKr41WHtMgQiPyflck1G9OHiQYrQ
9aR/ctVRKHx3s4q6ZsicjUMBCuwBdr+kGYM1w2TpzPD86Uojw17kWqawVHUhPqUkCC964mR/hsOT
ep9IbDVjoY3p2v3r+9iaYOqZ39k/XIKbc6YZhATQW60oLNGFkSH3//X+hfFRAibmVSbp/gxaGUa+
JkrfPuAm+nEPMSIVsWL6WuUzUfwNs44ek1HNucq/cucS7bg3G5q2yn3eNzqthgVjZXCQHNm7SXb8
LwLeUfSega4cBCdpA1NPrvwN7Q632AdQn1EJdeLnx3lHkjQe7p+iZ1xBH16fOiKbysBSM+y3steg
ZXh8y8QLc/GXw3tE3AnGatEGr4kYWdM5sE12GIYbOcf+VJJbBlfqCwyz2Dms6QhEIp8OpevtKujj
S3jrO01ZzyBRIjjSHG4iG1o8l/gDn9MTOUIG4hGTBOegB7tp2STcoJBWX/htBV45UwB7zJM2fABI
npDKr5/NCr26pLTU9vK9ZaC6rSVKt4nrClj0HgIq9CCLAuHrDp6Mj8ZrQ4y+hMxhW8oy/EFkSJJe
NhvkZzF2jp7OqWbKmqOc+7B/S3v7icAgPR/p/xCyz7yR1RqFBiuhKybLU5jxNRBVwD1Stn60Zn6v
0BG4dJFS9Ebsloq6TiBrwfYldL65AF/4R/aIT1zkkqVkn2nZ16+VXo2xgB1Ze687R6aRBFJ7k6Fe
K8yc9xT07U8SpeOXdHEgHYvOdHpxolzm+GWZac1my95r4mG7CYNMg7dKIFakiGIhyNbBNRvs7jEK
sQWzXbNXSQPW4nJagqEh/yMcIkkn+jJYz5qemG9y0nHU5E1L8UcAxqzcdasbOFdx5vGGmkf2rJb8
s06vY+Alzul8Jx7+CnslkHj+AP0/iYCQpX+hESo0mRTMUU7d4v7fGo1wT2sg9trrC7AsCueT/GUz
6prFmpWub42iNZdmDPUSuDF4HwhTQZ0z8/Jzzocg2KwaL49keOT9vs5C6g+QbgBSpgqviHw1O3St
ITIwYoA8ZbiCIXUsjiGi0z3JwAYqvTF7rm2gVbKIZ3GFQ4XTfGhIDhyzE3FKraIXnMNQIGS1/v7C
HikKV0xUlWEtdNRPHttEPxZ+BrxAhL0lHmjzqHSu/Yf/YtTwspsWbtT7GuPQLQ6TooEuo9ccFYU5
JIQ10ZfoUKubjcQIYW1/gv3+s43oTAtoYrcUa3cg/LgtY/6EiKfTGI7W2EaV5YIns3d3CKzueXve
1FdZN+bt5OADbkPiGecEaeYwbDvzN/vN3VzeD4GzkrDwSP2kmGtj7qN04NpLXvYQge6J8vbXEplx
U6d8kwb7140BZuP48NwWDEVxExGxH+aURBYdfSJ41Emu+Ek9xrwe6khomOZmVrPJJ1Lo84hllIlW
MgYDReQTLVbqOOgDm6Q9elI+sf5/AJXoes/mCjdVc80d+22ggUlF01Qd+1TLyyM4zszYHjHshU31
rpZ5D3Iaj5lYU3nphQUnPgUvOfoYQthH9My6GtBNrdj+KsFKKIMDAJfXtsAulUAO53YqoclXJftu
QhjFbZ63hotzw8MDOAEyiYdr1hw7n4edDR/N8HfkS150x1E4tgJnrElfmQ8P5C/KHI3IJGkjmXtU
f1nWxFtUkH3esbsHVrCnqJ8DoyjRiciOrVh3KIrwEy+E5d+X0vmTvvybCGIMfV6Gx5uZyhOYklbI
gDK8jP30ImLNY70aiEddk6P/ObshX5Abmf1j4KuA0MpNF3yjG8BpMp06TRdhUl0efHBhr3/i6sdv
aMGdRJMqLzrQ93bC58hgQidtuBS9+Ro70VAl1/C0CVM6C1/n/jOIn7Elcb1CJQv6OgjhxmOBLYJR
wKowzhNm/8VnnYpAeBva/xT1gAxYj+zTerxAOx3Vxa7p50OcYAEmp1RL/zsE300kro6/8SQ2QpUi
qe3cMGo377hxJIVLvifl/hOHwFY/Rt2Y89jCEAFTAqlO/MKJVZltDA7JjI0jZsPlV+6PDZkK/q+F
i4+L/4Azr4eMUN9kAZjApILOjmD1ReRkrgUQocSeqvYVMKCM5Uz2aldJOKqBxgl0BzYkfyZP4vz2
DAnxO/Phs2afqWneSe/OScanx0sYp8FL0QR73nBj69FfZrTv9JGHQ+0dOES3rhmY5N8HCtOU7Y7O
rZl9ukdJBr7mg2PMDAeWAoog9Bxr7LMkVgg1QKQsywsYXnBlLopGcCrKev+Uoxu4fIfvsbhwqrnw
+UVrmFfjD9oymE6duhURZD9uqkrEM9UQSQCFbO5+z44N4iKgGphrxW3nAw0ADoZAM5HKWbFpX79B
d62AWlMRxFYu0UetLW4S359WIIazezrQEfkIQQ49yYRHsBgKPsHVJqY/w+guSPLW2EPEFy42jCsG
O6jm0SToD/95bRXkWuWsKmRzHqYjfUyh8RKi2VO3ApRDUcCWKodXr1Uous7fmIIFzvZBwTxpT4Rc
3jBKyDCszupUSu0dTMEXFX+ep9fBW+U+gOPahUHBBugIRckK4CtGFGageN2u/cmLAlFR6IyxPP4+
1OXcRZapdjDRGcksfCOjJl9HByQZ3ezOeB4mlGR5p9jNaINRyka//QpNFyawEZDagg2RlE5bdJfw
USCZ4KitbV2fCcgAMHkhM79BIjmktk7nbBdz2M0GMX1QZqMtsZQNRJ27qWU7TiMPTbQUE68rgq9r
2gQTZ2ZBQWFDj7BEuralxUEg77NLCsSQX8R64my6Pe/dSpanakZGcH2Nf2DDuzUxEATbYn/SvYiP
KP/D9iQ5fjaUEMGJ93xLMWq/1q1LfmMLNJMru9hdpXGlpUy36mU5tJUlChfp1lTYLlAB16Tf07LD
Ny/Z56Nfw9i3K3/iSmJj+1DAGojzykzI9AnYsoDr2HmLV4nKwPLNkiflSm7xrMLIAsVSb5mCIsdv
L3wFdBozfWWjGEuG90sysH5k+ZD8rFHyO7xC7mTHLm1a/8p9xUzL34OZDzINGa9KY0pr99RJgXoL
p/n4onPYQSxkQIaT44Dml9ijXSRSDyZJOy6PdA1vlH3unHyy3POScn6g6/Sq3MpFpiOgGR4LW+iF
bCKUbbAb7r0XYhvGxkVRc+i6KQTAxVIwmuJTi+I0Ui7frallh91F66kAcvtXQmP9vEXe+NfhhYi6
vG1JOCqYIOnNCECiFLcBeIHUmq+KPwTGbEONJQGaT3AbnM/4h/ln0iDaQeGIQpSDsa6yqtNfKjhb
kHzcQi5wh8Q0q7IJKjT2ZktzkqUodUINpOstui6lto2G/fVvI0YhntEt/FlG36e61hgB4FRfMJg7
WPXf6fmdDSPT8zVXIzZj8OYxR+njPtKRiTLzFMFhQYLan7HkjPNaXwvtUqAfkcfiiN8ZWxv6uy+u
5IKBVlR22Q5OHVgb6wPs6MI3Jk/C5tZ5qHhoGLGLTQh66L6Rim8hBXsSxP89USFuUmV2DN+fN28K
k0w33osU9BhFNNDfpaTl91L37jXIZf7SN6NmEPbTTWAX7r7kTpGvHj5nMmtVG89036X+Yfw2ufvv
kyxFmh3rYL0KSXm1bG6bYJ0jIJBcZmQzPjZQsA3awalXE4dyXXFZdQksiErog+9cp5f6YJ/Hm+wt
lq3VwCbrbK1WE9LPM124YHcJ6Z3Tv1T27/vM43r7fS/NrgBTySWRivc7xmWRxHGDnlshM4Siu9g4
w6P8DGmJcA5FPRBVbSbojag6ruTEub0gM3THC2dIFTxUH2Fi/LPS0G79f2IIe4tYTWlWJYLmwuRK
O5ZobuszxFwrxuqUrFE+IHqYuAsIeS1eoDqAFmuvoxSQ7TYP6/vGfTeS8zn2R/EHu0eg+C8gLs4P
Iw14rsQxqjAVRsLSqkMcKy4lSLY+7Laxkvk6QZtzWgi/kbRT9YsZcQPOThTq55FgwTUh7j6gFfc4
ePfczWy1CH/feYjL3/lfWEY8UdGsr0/yydFKwmZR+1aF0xjC+yqgJ+EH5ab5Tumw6lOGCz5seKb8
3Ug0Jphj1xNbGbrgkm+Ejo1ndCp6pZKv/IyyFIOZ1cN/XFdhu83NL74+QXzxaHJovTdaKe2hWFYe
IGDKN02xBzFv8jVYrykzrddrzMmO5q0MO8WIranWWzVTAH+/az9cBz16rhv+kGr1ISGilwZGk+H0
wrkebD3NAtwbhtyszJSQ0F7TBS6auVSD02HvvPHwfVrWRLXo1l6/29bj0O1BW4XimA21q7SUa8Rt
R4m71gwd5/umyKd8Ags7v/A9B199w5oiSEH56ZOTmUSpgIe8OaPPZnyFWbxmDwmD5+Cz4kpcgPKh
QQW7kWscKqxywVN4J4qu7NJNLPNhbNOtSKXs2ML0QXbHaGQXOPkEBQnk233s2L2bbAtan6nT8eZ4
ml1AFUgZHRdmJnnu17WcV0kuGM3lZnKQ2t/TvHIX4tozghRC/uRJb1OWrmbxKFLL5cQ7Jb+8IGjD
Unwd3TmrFGc2cqtG8hmyo3ypxtZ4IXwXQkX2vOu5jL4C9I6T6tjJ7eNv9Ab7PsfSwDIO3qTYuRv/
UDKbgkc9VUpyQaDrAqGy3twasSJRRrroP3rdKPf0wfE6074GCvUNR5ExhsjHofzREHBGWVfWZWbc
5tNC/ElkXawmGGqivz/l4jug5VGdv+d6KWa+WxZeJ4QwEcuUPr9gSy6X+0ELy61+XUgKHcDAGD3R
iPzUeZn8EpECvRacZhCeeDKKMW7kA8t8u+DlwuzB0GnrIjI6UZkL+WCwOEDMySPr4MgHrI7k3NZk
AMSx/ZoQwntOu65AppwigoGYZzJMJmTnT9h7PShFhV6zCNVLa84P/SJmk3Ya2frMjJkU5SFtf69o
hV+moHnbbr6efGW2cea+pdJ+W/i/J+iwsHfs7lBUr32ufIBgJIxETx9KdImHg0brksXs8Qu/hqV0
jfWRg1+qOFumLNuMlkurflwHyx5ImtMwN36Gl8YtNqnnsjZpwdaY1H57QaqoBPyAna5mLbsOLX22
JnI8DfWHuNKojc5p+V60pCgetw61TCdOFl6OQR33IyJUIB9YFFRTGqUBA9zNmFQt6u54ZdG7Ee+L
Cpc+OZRl4Dya8F8S9U+nYVpaT+5iFGEjTYW/AZSs2kCxgCH/WYYzm0BtZ/RE2bp2xTjGFLAd6itu
65wc3wfeRxODQfPK+NY7PNTd391K957n1tD8A893fyqqxqC+PERdXRdjIOnEgy1EUEp26uJghwyl
qh9y5yfHd+DvDUtdG3QGRs9dOidwowX42hMCDRAQIR0Vzgmw8nzJmmfCD07KVaVvab4b7sjsH8+j
jVjWGAo34nBK9ZvBNFdvSeN3cAqIFAiLdtDdNrD/aX9cg20PPCpLdZrzGthX1HbK2BhgnQebRE4t
uIavCJrjywrvXWruCnVlqPhnsrvWjyf9pO1irF8WejR86eUbRrj/yDBSV7o0Sixhcm6t2kQoBKMn
tXEyTDVlDO9pz1u/efL8Fbme63yQaF73FLc2/gxDy8nKmaJpNB54HlIoyN2ItFahp+AwoLV6qzGj
3SbxmYd7GGThKqsDnn0gF/qn2cUYebiNS2vESwAb11MHKQUz+VuGj9Z+6tBqmvjen0ArzxSzmN3t
HauSTDT5CKDxsclx0O0/+CcZfRGFUOZWNJ0zfoVX/0WHgrecjgqMkFKesrZt4yfDP8O05cJkjO/7
sQr84Patiqc5dewFlVl/RTMmays9GeNNDxbTVdZ+Zj6kSiTQCcS5XNmJQQrPwTU7ObDwiP8CCCZB
DnwAe3V5OQQkBHFQvikLa/oEWNAZxbAOFgPCWqlsU5v+hfZtBdQonin69Z7tChVW49JSgBEb5VEC
EPoV497gJ1JalXHcGvQ+gDbTfGPDuetXn9R9PN36t+qJmLl6whHd9TymmSptn8+DrCqdAPoh58vN
+UZr/sSJBv2qcbjPrNFevTmWknowkZGOaaSkEKTqEqHtwjQToqqH7m0ma3/DLr4bmJ8iB/GE4GdB
O6RHbhL4j6chLpkKzQILHjBJVqUDkROWAXwdVCe97WMa4DR+vs1T4T6QaNujjMf4aRdHlXiYSc7C
SyeTk1dRs4gbNJ57d3W1BH1QYns+6BrZDA6hfmYwiV1uXPDnz+HGAoU+XrDU4j2LyGnHcAdC93la
9hGNP9RqUo5Sl2AHGC89kaWv2wApPAr9XuR9vpq7z+P3r0KToe04NE9A04zU27A559UA4UFGzcQk
9RT70mg/NQKFC2engkHZWFC+L9bF7geeg6vVFHRvKgPGFuwwBVV44wcjq0mFO37/UwznEpwsIY8I
g4Rv/AwO4woDpUpm2PxVuX02A3Fk95XtM/2jRIDzKgbqPR+cDALA656kDEpY8gswTpMc0TdvA4xe
LMXXWX+FihTcy9wgZjyX0kWrnIeqXT8pu2jNXp4OLeZKIhuJ4UBf/5l32t7DSz4mE2147w1AWy2L
LK9t7nQtyQ8BNyY3pMIOEJYguxMMILLJL3lz7VzaBIruhhDWz+KLb0N/8o3onDo3amiCPROr6d+v
+Ruphh4udqgKOz/ULG3a9iJ5xZYdT5n04LWmYaNRYt1RVW3IhI5sPDLxqrMQMLXIKIh4lsvRA12r
w1l9MAmyt3sFkkxGzujGV+Y7cq/fyjI3NIkinB233CZVAugJxhnN8YrjfLjQmPIwKbg5Y4wcyVV2
IirRV4lOix63VlJiW1pogMAWxdA5nYI5VkvvRuqtGRqodfH7yBvxsK7XKKneDJ2UlqZ+vXVTCuNv
yCnTn5Vfh9P4C9sl53g42XhI4w3S+uvphNbXDGHo3NYDciZXEicY3kMRYz3n46bI/6B53v2IdyqG
3xNjohU8vG0ehBmjZI9eJW8berLyuv9e5J+1nGd7ydMBW5YleadGeL21KJ+MqFTT/yq5ygHrTLb3
Iv2wM0AaTrLby531jx7RDiag2puC9fV/ImQ3e6yKoGwOye24c1sM4zy43DEDKX1TbL9GgYGqPTrD
2h1/jTCjxA6rKw6OUoRzv4RZmJfwNUCCDj1+yCBl0PjsSrWBDamXjJNpE5ZhAZGK/9EnaZfQH4gL
dmi6hptPonQzHHV7pJPOJbMYvLrssL64AYSPODkKjiBR9gfgVA64EzLxRnNqiNT1cH2GKQ6FLL2f
n5/kDkMaGfVvQ6kinNx3e6ypduor1hh6jlaDPtp/Y57x6uJ0HxxOZIJs+iQIjGQ8NE7GTfEYjWG5
O4n9p48tKsKyRXV4ZpNbeS/2CBK4s6XaN4EahaHvkoW4qmJ1V1It9RDFeQWTEFTmsNflMRgV43wT
sbfBt2fOTs+/7eIjnmD9o0GrkGBDPWb5+yItCXk1tpBFT8ozTolEJEVo0r8eGNYQJGzgw0wF62qp
Yt7spOS497mjdcma+8wqOjQec4RiuvBYr+QOX9oulQ14WY9b49XC4vCmnGOMyexBBpSXxN5dafcw
l3q64/veC2c4JOwZz9/SpR2Y5PyCLb7iENvp5W9/vtyUuR3Ug73/h3pHbYvsO7tkxdVN0olEcOsX
4hKisqLj9oGeznrnvYIjw6nAY6wJV+tmpPX7yl5aQ44EArlte0xKynfkv5eZ4L0yi+u1eO17jQ3j
iAql+Ou41cnMAVki06EMrNhJK9UeLXLOfOcyLa3BjvjlvGZHxEoHLkAVmCl+c76xME0u5+KoU6oQ
Op/mIdGhFwefp4XBto23reb1RG/zzIU0btlkXa7yBJ4FoNg1O00SSAsU8WtfsorSR/cj3petTwf4
7GT7lb+PCjFFhFvTJoICD35EW/+AXyuoFeb8xwjMdLRLRwmL8eUmn5SCzmM4MsSiA5L6UVekRnPV
4ckDehkrGckk2TfX74Kkv3XCwbq3H5SjR7cSSIeOTFQ/hJcxiCIgtn35WLubuwvUntjgOmko0NPF
xIiw3FJV0ueZfHAPjE5XG6JzJK7Vx+FQhw4gaGyGWZamrfRNMUUM0gFWUpn320R42XRf7CC9t3Zm
BBMoSccxz7sWKl+LeYVe/q2W8fr3PMA/JWLkEy4qcwPnghpdw3VTttXV/kC1PHMb5lW0p8ET82bh
Iu+HvMMjqvt47B04nh/fQvmEVMqKChC4aSmU4lDLrEEjXCTkWXxM4UmGI3+YkZ0O/RweCljR9Ucn
R43uFwLQRN8HgdHVvQuTKtHv2WXg59dwWvRmKQkak6cFFRc0ZQbK9BvLDoBdRIjx12k/e7d6SveW
ljk538QC8qTj5rLx0Hz41pe60DIckoGAqhnONA6CPejjLa3JFmdfIk73d6DQGgx6GoFcug5ILma3
tdG76P2j9PpeL1QYNZIbMAc0ZB8ocD+gFprSrcD9dWDzls3lrc4k3qThCbanMyFy0lDeG7jABKZz
84nLhXnR1RSv3zBws36qcbaI2oDHzevBbjx6ocOTcoHVIk8+O0n41FT1dq917NbouSnsiu1yxGYJ
qnAbsthLTiVHhyblFDrS34E5++NYxoE3we3VEynGfbQcvhDpVMguQ5fWKfuvuwj1qXpH8q05EXTr
Zdw71/dE4DKoTHH8TsaD7CmAiqpLfKeaHHwZInXWHMWSDOt85yePeHIyV1IvtSifLdQzgJpUDI8S
qtMbYYyn3zkEynw45bn+tXQU5IM/vjtrbeo51uFJV3TbfekJ5s9Vzu+cHB/SyJqbH6juH14KDz4n
dVemGop0q9bVEAUaFi7FHHeOxxegDVwKkAWA2SfqtwKatJvbQOBXwwA/MMB9gkI5qnx9tQEGmLTO
7EO/qibI2B9hlKKCWxQ6JNvi+AYVzoLXyYv7NcSFbTJmaQBHcDnq/9udd2x+wypOwGBx5aroCEkQ
9rKhW4TsUqZciV8DcqM87SWz2cCAu+NspZTUTEFv0WrBrlugFq2QtxgPrm5dFmZMA32yllZRNQz8
ccCxEcKPpfTdXXBUdAF1nS0NTes5ZDmSImwMSJ5BgLUxlFuAUYXQ9vo+1TB+BHnRYh8ZPqY2iOnm
13JV2VbWkFyF/Q5AwqHdlJ+swfgUEHZJnpOt+WMjaMlAy34jbL1Q3C5sduR8eJhGCw9fS5N/yAm0
DpL70JI1Y1YB2lft3F1XCpRMK5apQajCCWdI2jUcXBfsa2pbEr0b0xXm/Z1Ltl7GTB+Ld/G5DPz9
29KjT+PgWh4bdClMKavMlbim5n13TYFSgaqbNkF9+9Pi87BuyrmJWXVCW1TLBSV4jY7nn3HN97T8
PTq7rya0ucK2QQieM0UkUAPM4WESCqt3hewFugMRJJiZkk3c8ayt/hBSpqaOUx7diN/GcV2Sdpcj
DxBlQ29oEVLhUXR9hHR8RkC0KWuMy7Y7dYZAd4aC7H46T5RVCpKE0sXtlRPf0Ztx0IRADFcgaP3O
vtesm5LY50f4DruF9Z/1F7BgBlP83yfquuTxyq/6V2dBKWevyvgCWhhPgEySKptLK+Tb+frIrwlu
kZAGMO4G8EmXC3vzGhVybw2BXDO4ty/3/rWtmYI9W+DuD89U6iGAeyiV5dZh5A1aIK6YrKY+UnEl
wl+anWQvT/J7Rd6IurphHdqJHbXdelkCdA4cn1+1gBv1tGTdo0S57p7PpAKTUMYgc+dMcyFYriAn
nrO6qAv/GJS/FRreRA4jl738oZ9rQ8vHWPyMmgFmb5qeYkB3N4nbesLKe1H1oc7h2KWuKOPUhZs8
TMWm404T4fghHO3BvBrjftk4uTOh+DZz8aqBmbQkt10khqRTFJV1g7wbSVz1HiPAYKqgt1dJyzqc
p7ESiZuAZa2j9Ut4FbE7lSmvCAwx9RQkweuDBqgCCtLUS+QMIa402kVTA7jYmgbVNiZoqksJxzbN
XYz/Bz6oh6ilM9qviOgQIhrBLQUxgGudnql0CGYv4NH8Z/JfKQzDPg/eJDwzBYb6mQBM1JbSxPJ0
i6MTpnrSEp5l7MlyZcKdb5/1D1+HjN2DeNNddvf7MHM/48wIY7Ipia9Zu54tqFF5ySa7hPgX86hq
hZ4ecqh2QNUmbIp3Wus8wIs0N6zBy84OWe3rfpagF1iXLX/GxazHDBB7COlNmbeGZJI6+py+1i5M
xF8KM0nnhGwOGdB52C+NFPVwmfQ1ghQ/dbRJhxMLvnZ/l2pgSDLyLgIfjx9LpbPUcZnj+E/7aeW0
A6nHQjPex1CE4nW4e+nTkvttYYYDwBk0Wia9d7gPb4MhWGIscnbkUfcIl+hw+BOZF9k/Ohe2rI2u
EL25bsYvVSzmOFxrviO/fVCRtVtN59dNwytZwt1tm4RLsro72mwZMWlXdB2sD/4kZwQlTvkLCgls
bF7EkWpqdlEFdX/ZU74TpCmP6HgTClYpqjz4M3jfMaDmx+bJxRoDg4hOj6XEYzEwnp4keesb4Rl6
X0ouJn4zWjcsL7xs8sH6NJEs4JolDPZpGVIitL99aqVg2zE/jGQFti2ZTCf1hMzrHeDSFZYm019I
5y4X/5D4ApPfA1lY9ewGffrRSa05d9gkWfDB8oqNIXsl57jpzcNpYvJzVVBJKKxps0t14cKIGVHU
c7S1gEJfx0mAh1A4FXfP5x+377wl7XwlRdXzd16t7ykAMZjxCdF/lAdAf9IPcnd5Sm3xPlhY9TMH
zjxfFCxC6HOtJY58oCvj3Hz/CYwTXNVo7qN0b2EtHdUlc66nzuKgZXAPGhHMQT0HU87ipbBCKOBx
swA7+qhAYEZ1g3OBNRj0CMGQ8deg+vO3+YF2n5W18hJXPXwNFCCHafzfpeoKHyuCM+l7USaKLI/k
FxRVdZDS79VMvj1mqkojfPyjKc99riWWf/C43avvyVP+fPKB/C6kGcVLc05z7yk6/wpl5QslnPDA
gqIk584SoHkxRWPheS49Mrc4QSMWj8jOoElLecPfxCZUpgWd6Bg4ToXpIwsyu1wWZTHOb/eHFfsn
zMXyDvQK8lGUYm4wb4121l4tBayPE1AEv0if74wmUs3JUpA3kXuAqS0o4UsztzjtZfTAKPXhxnf1
c4PCm7Lcf6PI5shCQHmmGdOaruXFPr7II9fUj4NL/ApWOTVl9wtmwAvQqU4wfp0FkVUuKt5gtoMH
phS3i1zC0N7kD8oZTzsqdTE9EWv+JUwKBjM84FqXPK+L+PEWuhlZQGqMScgUNltQXPnKqljxVgTY
NbD0L5nsDcgHMfe+83PnO8YTJgYPtea3CrF5yG1WzSKw3mP09sM3kL5xy9V/bQEcbZgnoh4JoR5w
P8Z04cVN5lZxGctnVjr466iCCw5bz4gXsn4+GpZErh4gOEkJ74BanVEB1oX9+jWi0QLYSaY51Mjk
MxVuWcjA+jRyK4RYg/KI+kAWVom+hR2T1/16SeGEwb/klG4guP3XiLGCOE/W+xDqeZBb8v5oWgYy
mDV2Wwgzo76rG/4qOJYxbtkcCJ8qjQ8KJxvINuNx5MI7a1imdSAbWQOib+3XMVEGQm5JeK8osPQO
cxTCik9+BH0j1C1as6nlyFtUY5De9AFzogZjVzYuzyASjrTHAhuhDJKmnzD90HSXU/4UjfKbjqXE
nwuCUvs3OUaegnkdmo5nc2Kb531kbUqxUF/TQ2vIfikTmSVLV3f3d0x0l7Cu75jhAn2EYLZ0VnWm
DeapidIyVjVKD0ixlus7MQyGw+cPGhTuD5r40uTkx4Lw3gbWeBFiKPwdmql/lIxb49h8z1fQUsKl
BkLZQlQrH3i7oDi//fCoxwLO9uvskPEvYd3KWhgr/O3iAB8erbPdEg4l42kd7ubqYKlBmBN+4AwX
q8zcbNUwO/dQsnQRf03ZeIBqERNKQMYWjJcxU0laeyLYgYB/hTZ5EbX8117DOFdg79JG0gB2ldSB
5zdQsftyhNTlqJn4REz9jvRL7H03q+leSGJAqrFB6RCxDCEiS5LalgdSca5FCevGReZbFqnWIEDd
cYmYxL4rhpIgLaaNH4GQ9+mwL0uV6dPZkHE5ZY4kjv4N+CejoBEm2rplv383j2l9H/isKS+Y8aAT
s4ZLMTJbBj5BFyr/hFg3QSYNl7oMmi2E6Bb3e+zOZStzOdYaDgBgE+k9IoKlRSEe23uVck/GsNxA
+493vs6lQPqGFb0QIC0PCBBvDfYccOgEpSuXHTn9378HGHiO9o+xD7Wkt0IQcgP+GBbtYXXcu+4m
S2mKzECxRy+Zc0U7f1CiOHH78wBh55GWNBXnqT10Z2RBWXLz7jmwGD3tIfT6e6mqIoBqdChDOpiw
u0wH3/Aj0LGR162pXJxBykIhX7BI3LUdtfn8colOcysM8PHhkTU7tEAFF7BKDpXWQhyvQ4KwgQMo
8Rtt0Q72ETB++YbzI+9CMgO/GRYuXNMK2mL8G0GqPZA9CXV+vJiigdgE/mrgH15gA2gZ7kcAJ2a7
icL+4zKx4i6r2EN/F6opo44cwQ9XwePEcrgAHSYAUCq05p2GC+EIaGdUm4BBFWWLPrdZQ8J7dpDO
shgo48vwNuJR8d01s6+aDJ8JOnTRHHFNHA84DY2gHQbX033xOrafqRijNGPz4Jp9FnQWsG9yAE6z
8JL2I3rI32Ul2jyNBetG6akdnsb5wjn8rUTglyZ77Lb1g5FsQKXby1TJxGRPc2E2KRFziwoMt6Xx
BPqkLsvPeHTMvgk2kMb/nTBrd1Ipmst8e4xXjNsjEWe9R53vmIuIXPVTAxsfT0S5II2lsOv2BSjm
wiqsyqBa8WYGkIBBeDyQu1JNykX6+Dj9QkvXVNvXHBNPiMtcWku9TzpLqmv+pvtPK5icD5ZrbpmH
9zGh5lnc2TEr5Dvc04V6o5lHUxvfPXCm8tg9/uvgmN4V6H2BJ/h8ozS3pgMHOL8IB+J5rtyCOLYp
UnIjObi8hhLJ68CacuPk65U2lvir8q3eYVBd95Ok9Lu8C4kgWsfjQuMU3gjyOOGUQM82UQ4tbp62
tgqNoJF6dZHEcaaNYECDtWERhCjZu/KL5A17dLD6FxTpgpSooaNJn94gKfoigovxiVbSH0YokjgK
x+dH32OuZYJ5IIIxwxr0D95EEJF8RYd2Oxwp9eK9kkFX7fy8Yaz9U9D6pDoEQl7xPSRNboY6zSY4
enDV3VprERfR648pez/36ELSVLXETUbIJmIW+SuK10v8YLErJXAAAa0iNIC7nDpobj+Agzz4+Ez1
l+9c8vwZogsZaWXCAt10aFx6DQoDV/6mOryEoFdE0gpTMs50n1gkuuHBlnvAjN3oVU1N4squuf9w
TmLO5ZOddHQzktLXDwVzOrLmfP8dtTEgjID3t96ty2F71JFjth4KURqNDlfkRMPLu0Ve5xzYvpDw
gUGpQQcNVrTzKcAPnTyzRHVdOs9Cy9AqvQFVvTUZL5NxZSCco9DpseiwXsqalXWen+vpLgGbD/QD
eBclevCyZMmbbpGNGGRYSGawiDGiRGD4+eqvut0tLh4YMg0wFm9pWRPAlhY5aTd7wZ1XHZyt2MTd
liaS7bnDFLaxcD0c0qHvMNcSVLpMzVC8DuDLi80IthuMPr+CU8QONZMSgVLuLb9bhcxm5h9LpaNr
k+qizx47QxbZmX55qBQLvUCDiUWB+PvhOeV96avGTsHuwXPXJHvwTA9ruiZ8I0s1B8nRHkz1pZvF
NgldANh8uVn34gMV6vka3Jvm5YOXjNap7MlOgMB0BccKcMnxjgwkXEaB4uX0SLgOe5axWgwi2DGJ
fCZu4RLTqDNfkONw58+KRjzPZATho4Y1wFz8g9jkEbzsFSElJFKSjZEWN88ZnRk+x80ECoZrhpU8
AGMh2v29L8rGWqenmNL7JRL9Cvzvb+YX+HxTreGTf2AmzspDE5UXDEaLZRI9Zkh3vrd5Zu99Mews
POAxIDQh6y/8yTJWFos31hPYO9oOs6TsEhd8oV/EkaEZxJGBaseL27OOxFLPE7RUGgsVrxdwbZ/J
gPCIbdqmbFjpc3j+n6s7zPuOUnf9PYO30d41CFFYrHan+SEcNEsoN81raGGSIGpHJ7tM1i445ij8
mK6IhpRq7QCCOsQ2U+JUldIjvATBJAL+QxTn38+uQjbf+NwFBkB/8fD30GoIiiIgBZyn4HzMT7NH
mU7eHR10J8xO5cWm/HtFG1+zGWMFvDJg25AzkPHZTIhP9risvA5raVrIuVEbbhgu7GW2ddPi5sx+
zjR5N0PlBV4wfTx8WR2hwVvJW9Sfv201AE5boUwIoxcS6YdidI+R00wfQcsdsMhp6lUqdUMYqVHc
1PeHeQ+4SasHC0uHJ+bY3dRqYya6uKqUW6R7Pk+I36zDXBzsyNMRJ1BOaT7deuQmxY9qswqQeaft
jQtVUbY9xCiB1U1+7SkfjuTgto1AGFCCVlRBkrMePstk7UH6OvoS5KHJY92MxjXs1wi02TGTWGG3
Gickblh8qzBIyheXWpCOrQhvvwj+RvuO3zA8OEC4T8FFLU24p+FvxmsCVgTzzYFUVjr/s7BVEUr8
ah0IOxAe+RWFlrF6JEPEz4DR/lSbuFohoR8ArjNkkDOrJ1lwKzZOMwU1F4kOjcdBK3pYR4T341gE
BYSR+L9bTW4/AcFmHSxJyUBnjMdMSduL0xhiaBbG1ha9jrSFNaNyq3FATgrXGIFYrGF/hGJF2rwy
k5XbN3PNpOhgXqGatvOlFQJzsh0YvEfwnnQNSLUidrpxZhaTS2XU3BO/WVoKaENNgvY/shNiC84A
uV6B9eDqeNzVfHui68E/QhjzBEpY2xOa6Ha0fo1v4rh6v6WYWisxFwgGyuS8WjYhySnZi48vOU3i
vKBblXb1OL9e8Ed/X1jSAgt/9Aru8mKskZ5PFRz4lIz7WOtlxJM05NiEhJR+WSm7qF7l/0H4UlCx
2f/bhj5XBAQGnAbngeoVZxsvt5JAv5uGaBE/jcJ9ze+j/s9gfVSGeG3EVDvuqdgcJbn3qmg8wCoi
mBXTfwtEHJP/ShY7lQVWyXKlnly+gpbWY/nTZ4TvNqspLAEYWmleZ+j+kbqrh6T0VS9LP7YH0jwt
ShFO50t6QefuCuiP2DPu0rv4ordlkNkna/SOHVjCoOCBVuOwFNdSxiJdLsoYppeX7tfxLEqyPIji
xlZLH9coeRdHJATi137QV++nxxfWWHeLn4H8vg8sFYN3hb/3RKmziRhM460trfqgv4QC7qO2rCt8
4TlQ47kp7HnXctnfiLdtNbrK3G6DeAbFdUzuZHjnhPbvPOsAgQiwGQyH4EhO+WL1PfzUBaXBh7bX
eUp6qmr/tartjDAiKfV7y6T5UK40FiNZdqQ5SeaO3lFZHx60KU2fzv2XqSIG9Pq4fKxvUs4Sn6SQ
6ioG764i9yldj7hmHh3TEmA9zSAcvW/EyR7IAeT/DdCJkxfgETzNOusXnJJTbvaqAigbEbtV4nOu
bTnjagxImukm1f+oN7oCcmk1/cHZmzGyKD9oDzUFd6E0LijYJYYLm+LHZEQGdKoJdfXaaDKTjca4
VHkE4AsSBacKwzy0ePEroMYgE9WuXKiO/P2aDeaDVoRD7E5Y+rC11mN/wm6I4yn/9WO8vDXydYR0
TommrM1XylYZYUBWdrRYW+M1xkZ8DMaDM+HoD0D99sdRNjw9VjRR6miZHSXLeMUd6UNwxV6Plhi9
YPdt8M7NyxS9ih7gDdAtbJj8qBB6hN+pFLWolQTNQjlEKWecAlGRCS/z/6e1o6McXlsbcYBbxLl1
RH5OGmrspqDkxtA8RImUU+G3RDRMpazwXQPI9Anfy1FjnDCvKxPyLgUMF1qez7qso+xeLgfa4b3p
MjYmWHFlUzD1xtIgnY+6ee+3K6y/Wq34scDb0ix21tVd9IggSYxh4r6CYNd67x8XyAHlR8rX4cGS
S0vGiwyx1CmYAD292EWDL9ISklPCLNWwh7AwQ4lW0R/Lca9rTwOKo4ay7C61du6NTgOSvFtKfpTH
FSVpSJVHrVscA8o0AnVIX10j5ZoK2Xj8rw4d1FNUZEUApr4ctFS3g3hA1CNfb8CvaksHcnUfnY/1
ce99HeJ+yCOATyTzTQU+B8IPrUMoxLoilJkLUKu/+To5o5ww74dWpNBHk6w4Z/CtFGGziRfrXQHj
Q66eeSjfA8WIXmPXECrWocSpRcP2LtmKx8uyqGU1dOXMbpHSr36tQN2ribQVTcGeCRbtICJdEaOc
JvSpDTvIDtYPm2m3UqvETpeZ4RRb3QiXa0fumtSAHuUAuQNbJUkEwZDyDM69FwswBuM41s+M4J/j
8JGhaUyC9R5+Cr9ZCAjqzI+9/3YOjNhKklcASvKcBFC8iYTbW7RL6S/hRYVbFoAGcQyUNDlfomtm
w3IBbWiu0cqdRf0nu+NZcVbz5XuRydiwunhAyYKl0rAXjuRVIPnr1DJ3yGj/1XVBPVZnPhHUHwWH
oWJfP/qZioB98V8WSGfMyGtOzIoh6mliFhg8p/FrqALXtfuMTrV6FOy+q0KZ1Eokjij3aUKrIuEp
BLKHdnaI4r2GNaXwAy5aJH1NApwIvEGeBEqvZb5XmWXLP53JcGLWe/cgThUr+sIe+gYitdUM99/r
WqCLhEubV4H62ITL8nD3KFpxF9lDrrP0xV6+kt89FdaH/iqK7iq+V7qCWi8C1+ChYkDbdxyKRDHb
nXo+qMGu50QuRyteSQK481aMayb+9O5wMs8bX8FVJJzwCmKx6Wnrk6NYVdkFq2On4JBMoWpSz4XG
Cua363O69hUF5JnCuJ4Qpc7kwFJwQb5YI0k5GX7VMAvpPNXJU3f25dKdCsfT4b4eUraRRPodrTHK
NDlPOkBXQBk7KZqVZcEil9auxOKZXG2lq7z9IRHujLELxzFRVmAXEz7IMwl7Vv7NQVIJWLIr/41c
5WXUNhXR9skkads8Zc/mGz6Ww9ifU7qSklptewLmIjhD9nBMGXij/NDrk9KuR0Zua95qTtDTFLrw
ZaxduuAE8u7LNJdtTiNjLNxkUSujNh/GSIv3a0MSR9SQ2PiuVoc9U7nz4q+/agINJSd3KEtZBkN4
xu3EYCNuP+d+uAj+4qsRk1h4uyj824mPhDs+zoG2Dl0ren16NbsQdlD5Wip84+Q5bj0N5hoc1u6G
u2N0Qv25QcQd/EBL6IjZCPD5slNV+hfmIX8V8mrt1kxYYStk8QPfOqFNcD87uCnGe0GWwUQ0ali4
lKQzUIi+FFjrTl86F49vZQJiG4CBST/id+xPMAndu5wgdlXrbT4YA4oQf+VZhCjqssXnnnR0OqjL
zN9+6/u1NW66y4ZYvPl8LJutHwBdnfx7ycrOx6Gk/yXDimMmCnmT0RvL+VZQj+l5vjxMWbJYA9Tf
kUS9kVxlLUBznAbbRYKjoyFoK2L06Jg0tlLJpHfJLtZu95qR62sAvjIFtHuerdi5S1iTaqhl5jMo
s2JTYvCDHg68ZNO7+8PK2sPSYXwqsof7JSPYVOy8ssvMdAbPW/rb1XJpuJCIkYf34hE1Q1XXwRnn
05qn4wkrs2QUz4BFpEEeSC+dsw+v8S+blAZNm4ZoXqq2XU9vwnC9RRnh+QaVgVKtpJYO7SvE8hMp
W0g6Zx1KUohHY2kR2IH2+384+YdLtnXfJX7rYsL5ktXIPO01vdPn6fIpgxvGMMn2wkhFWdy815WV
QrP6qqsdMnToVSEYlxRM6h+rKmc51e8skYIIwKjpGSV+dIVlosy1biTGqR1m1Q9Fd+hK+ZrKCyrw
LPwYi9lVrrUKJohACSG+O0JU2pqw0WVXuIUAU9DfxaOOrgIAH6qBTGNoM1VK2vKSUUalokp9u/eo
n9O8JDP3LnUApfNGNce8NuSk5Q+DrwD1NU6Zrs/vORQbcnmtzSsZ9Pj9tGRGSwwI68dZdpz1E/A+
xlyQhCzUbSuAHl/BurTvLDGpHbL9+t0m70zULRiAdPaitmkCLu9ACwoNP+WdSz6IaIC3CSb1TyPM
2J/Oz9VsBXMWJ/8fCeiPDtUc86xhSV1JWL+z5SG3Lej1kdPGL6O7fGYm7DJaOWq4BkCy8LKtVdYq
vuV3pOg6427a0/1DR9MHhURWfnpnFXMU6XgvHxdJrwnurBdle+hBxlwFnSizD5paqzahLOixW4tR
aGYnOPsVMDr5MQ9eQRzazmHtMaC/wtSXmRXWhIagVcczE//0kQUs/JN7w+P1wfco4Of8D6DYfcja
yv8W7tI8UO7Vkvs6a8PK7lhT3csBezAjsWdSApRDh+gX/bagwPUeww8JTRtHZUL/fCgnsfXC2GLG
f2KoeYI95HqTYQcqIVrwk96h2HQmJKpQTD4CmuIJMJuwX8/tWz9gOIBvdy3V6XsLO0SYFpWTWEl2
t5Z+94fB+HCpWN8ubDHU6GRo/DvojpoyFPQngLc9wDRuHHMUB0u879uSHPqxSO9oopu1hsFuHyyo
vHlVbhs9M2z1jfM4qXyiPR1PWOlwOnqiMb4ElL88q4xLyf5+Q60kFvV9lt1smruv1uLh6WKuR+hT
fWoUDMIo36++6UJOB2pa7HvFPKeFEttJ/GpiAGtkjlFzqsYk0H3rqgx0+h5T/hFJHeKzD5era5FL
ncVURuhju9k1mZoz3xyAhBi2hXbgG4rsOLL/Ga3P8Qur57rysa3EjmCHP3GR5g2MZohev+CPQ0pO
xWSXw/LibkZbj7lUDk9hvyDQ1LEvs2SyQ9g9acyLm2cWwcCLj3UMTupw1/hQaJTEV563QvDcQlEI
IOzjt09E5TuLsqUmc4WpTWuOmnJ6Oiv04+cWCDdIU4i5Ugp5S9aA7GWXgi2YRPrm+C5KTEhXbXSQ
SW7uExUpBACN9Y+tLLnn2fJRr3vXAZBeM8Eda2kIgn/ge+Tw+dQVF9jt+zva4H7Qj89MFDm9qgz8
Oy1+ayJ3h2Q1naiH+P32hNlcS6tjek98jXfxrodd7RF1nN+ScG7koePLiVUAQWPRFdEyLDzzkIrg
tWK+SXACRd1TWSeHEA0vSDUspAA6xtbrM0BacJJ07cjxdvDb+n+PiIe65D7sD0ju1cTT4hhJLjmX
C7KZQ/kLh1ROG93j0MHkByzC6LK68xYQ5SqN7OkUm23RWU381cLGGX4qnKI22hYyAg1XZ0fOwUJl
HftNPaYI6isj0lpcE4EFEFJrMcXYzHZ4/z6ASnH6zZunUdSSlsQuPdHd7pKWMCwDGbQeS1r3NLFX
6AJjfMtrSIjw33lQB3nXAdngnLbBXcUaQknNQbOsQkkqoH8QXegyPJ8yoEQHOxONwQ8QY+4dOELx
AHvR3tdVOu0V8LnuAyGWS16HrIxyAebEHVUkMjZ+6B6axAWv+86C9ekGBeWikfYLRhYQoYpl9CjW
e1WJ52bkHrk+BgsR3tYHG74ko07jWpFBnZNHC5sMVNFd7QX2QuZnLVdDtOgPb338Rktkxiauact7
kcCVIl0n2IySw0fI+nXm4diWn1r5Rj+AQAypgPJ10to7sAUAO8cEugEft7k0ORz4AC2V2/3ObEfB
pVol2S+NsnY3I/DJEO9BpC89Vmf46o4L1Gin3HC636gxIR/wJg93jBqiKRVmek56xu2P1zy5qs0G
PiFCnKT/FRRLMH5rTsFeZPzoYswKgCgb8I5y53tmwFnDkEXtl8zQF7WiExTRVrRjrHwAPovLjl8b
LonQB+zxfiOchQVakCcwVJLSTq9TwAoWSbYIu/CFE45iFAdZHbBADdzQi0th8ejfXQSTPDTUcg0B
w34OZDKoJhT2pVf7x80LlUfH7qTWIPQ9amqw9g04Rm/2gsuaKoz5xoewlBLUFfnUueR1ghn+8WUK
SrKWDCUyMTmER1zsf0cjdCJjGFEK287sR1gb2JJNp3wORor955oBu4YNaEYTwGqhozDPszOumujo
1LRtFCKoTnfmkqsfbplcXmBid0Sf3xKD+6YQynhLa9yaCu3Rlymj/B2ZZeb5VYi2nGr03eECT+c/
lxdncHlHG8yAAtc7hhBoEGHz9YHoHTjsupo2c2KjOP3AgyH3haqCb80nOr+pOQUB7rFTI1yMH1/k
p/jjn46yVXM0TRoDVeqhYj4CiUzVEfKKl9mpopF2ixt9MgOUM+ZmWDgo2p5xQZVQVRtB3szHsh0K
yfxjX5wgjAuwzpaoyJjsMMcW96zZuW73M2qFQxOORtTbhVHBDPfhk0oVLT+LhJTbJhhUN/jo9X0v
2TQaT1pPbku/nj/zDCB9V8eJiPXvHBvosGQXL7QT9YJb9DlwuIZZA1pzPp5wyfJQKBOW6uvxnUa8
PEeVttgp8shxj1HvMiD/5Z8fosk/w//Mpu6HcjGK6bs/Kr7h4dKoLLoQuXAkCUFx6sbY66cfDxbq
L3LeGPyKvwiokdE0U06M5OasDJd5yxTmS0y6YbxunPSmE16gtgbNVQ/l4hNPzR+KJ+rfFuryL+MU
VH8MUF/Y3vpz9dBQTzfS5NCvvdV9lUoppXwMKIUM0S2hdvB4tPUeJB/HlDU3oqG/Jz/otw2rUi03
6UuxmEH+/s/yd3EOliNsGfLpkZD9KsZxLpPE28JbrKRvU0fJSDu9SYMpkdXlnfr5opKQ2xCRhv/g
89NOzFSCD02U6VR1A/lsgSdSdpGuAev/JlyX5wyUYlrbr/AblfU7adOLNqU2fXcgET+e3Lypxec9
Cp6yh11XDARXPxWYBu5ZIZQ/zlRIuSqct1QjPcg8fEzWBs4Uf5LTlX01fKtGjnB4CDUSYGRZfaKE
uon8xatUNejT3PBc2wNkO02CMYWQWs8yH+kD08z6EK7wiDmiQau9E/kSuaiPLxtjAJ7TIb+jdYPh
1IQ+Fyp+L0Dj4trF6l6anh9m1hTHvxpMoCuaE4/0FPGVcSO8dsCmjW69FyZ6vHTX0fXCB/lvDLLc
igxDTEGx9lp9wsHritdoPUtUvtloaYaZLI3LepOzzNZ5hP/0ysxIdvX0egUOFwmnEec2gXHbJn3l
P31tZe8h62HuYt1h5cuykigLyu3OdSog86IXekQ8SMxR9v6QgYZThGX0dCtB3gASMDsFO/XGvQez
UOmvnAi6CwNzx1/utAcAT6acd0XsBZY0ov0Ph3NCbnas6T3Jixp06oheBTFDdMPsMPNsKqV0jO4x
iYFc8ZEFUJeHGWydUb2EaVvYlJifCdDc7CyCFjMBE3qzoQeV/KGOrjBKwhFeQaj4VEOjGZHd4FXi
jSYx7bHqLWTxNq5V7EyJZNOc1WngCcQaoK1ni9w8smUpRk1Mzxj4ylTgm4xc9ps/apG1BaxkbKbs
8TzO5RhDwnIwdb/i4lgbuJAOwbxkz/RKzgAPMuK16TFwzEk+sXZxRKYID68TtZDrZoUVIvhms6Wu
KB81QBOBWSoMpKKYKXgMIroUvTHb7iSbD1MB+USkw7m0nj+Zo4WYp7p9cLgeKpYw89x43ob6bGWZ
vwCMl7uDBIAFMBuDMtTNMO1FYtHzLOS8ZLM6atf1Bo3p35/PQN6eWKgjVvlRTL2W741Dy36Dy/wX
X00rBB3/R/lJKpZt2MC845ShdFSfnY4/MVasQPmwp+CpPs9ZD0ydPfJLGNvVE1Yr+qQdh0h10KJV
d6epMO48WcSLlBqDMc8FqkFLhFI/NwiBRkTfDnzj7tJyjDuiFg3ekA4yS4ksbS5KUeQ13YMUR6Xz
9ZAgVC9J9zWp0f8Ycuva62KFeOYpyY3RbbouDVlsAWxzqJx1JPg1lURrkxYYdMfPvI+enET1vr+7
GQVYobbVKAkWBIyuMYJ2YiSFgznh7YYn2ZkpdjNC9WnMq8LvOu4W4FXa+xFSFFHOPErMouGvQi4l
5qvOqqCSadEmzNiuvyo1abjmEm8LrQNqqdT3HeEJSmXnha5dxxwkXP0vO9LekB3i3noRno88Sxrf
zk71ijCM0wAaQDNRXB8/p1vD9xsMzWjhNVEzq4ylXVr33gaBv1gOCJarHmdfFfR5QWkDZ7gh5VtP
b/DUwUV9K8t8DRnaKfawy+oecLFVIOAI/osTUQY3YkvnDXMMcnyPbNXXEvXjPghDmnAjXYApiuex
AGfJBXzeS/oJcsyuJq8VsNCnzT98JcDLBn06EgZPyN9vg0JHV+vFFPf0ozDnwUZdkBAiYpNUeXEl
hbiU5ftHbdn9ihYYfhrTBnfz79zYY8v07MXl2S+ndBJgbEESk+cWbdNj90DErQ9CrUTGpazHHzgk
82IOvjYKKBoGHLvCboMxLJgnqjWZCWf3wBy43Ax0p22zYKPjfhtowPnCHAfWotivGaPjkF37Tf7A
NpVRczEzm+GrfC1Zm3mDuBS78VSl2EeNNa85sfCPcFDPPE9677uJtvrnsuX4K/J03iIiMD3ADec2
IxGgAVDhtECud1ihAbB+R9tYzZxseEnOh/XYzU0UK8PpFXVy1KAUiC/dKCkqm1TgO5L1lxl53hgF
PqdAR2xFWfRfS2Gyw7Ug0w3Sl4RVKMkD49GWj3m5ggHPa15WaS7QbNt790j6VCAcgDRUkEBWotkd
xc+qYBNbM7BXRLws5jVth8IAqp6NKuYLjedzNIqmM9PtDZ5z+V492HOl9US38JFxusQjb7fXcyU8
S721KD92dYt4XKCxcg/3699XEoc1kX+pl7z0e66a5wG1UT00b6Bf/XFkFDxSQ+KAU1MDVzcc3BPw
hYhtTgpcxBKEPgzNUgLjYNTfzfklfp03o1wOqAiNMu9Q/OhhRkYQxoaiQOxYKNUxF6iOtv6m64Rz
sGVnViJMbUtoW2LthgT8TBkGRulhGxbEllYDfCzJgXLzEQarvRQcTsgk0DkInMvPL9zwYd/CWqze
ngyimqenEVqx8EkO/3TdJSSeps52yKtS7VtRxtpVPEZIiWmyT8URYj02eQfwlF14OGC7iyA14CuQ
iepaZ6F4usvrlCEem4q08aZ0yPoHMranOIPmcknQ0QxkEIg6WJptwCJ3bQZNMBykdQPZ1qzHSVW+
kO1haM6JNF8CT2EpPmfY8dD26R/a4rSX7SULfP4ZirmyAN+eaoU6gLXVlwAbe5LKh/yUUG6ZfhX+
ei7oalx6i/IJXdoD5+iHJRy6lOUtwjKqTu+IZdNySHvjuDlknEUAemxlVH6YN14uieRYcxtezsRS
s1T98YmIWrc4ceCX8fOOYPsh6mw/LhAHfsCMEUqrIRA+rNeSq/rVKYsDUziMXVFeZ1UfpVs4q13N
lA9FUlDJjldZFCm6luTg0LLo4zbCUql7TIE1sBq3AMfycgh4qACEg6+G47Ceifq2Su5S3uQP/5AF
bGrsfKxHdydVohsYO4VmS4+U1t/ePdGvPsVTfHRtH5wJ9e6ivP3uFmcGXDc0feW/XAQaD3/ev5QZ
2GxZkL3Yxek45v4kz/3fF9JivYEcRwtQyDtJrBs7NSCLCdUiE3qZ9xI7NZ/G2kuWMsQFkLZJLAq1
8qIsEQXC8xiojTZAWU5xDXXYrjubPCo0f35xYOpGtRT/wszCUdD69Iflhess5UKeqkxZlitjW6PR
b/wCCLrbRryi4zp60vqAIANOIIJIuZj1luigMF07xNAqcm5y9VTM3CUgeE8uJ8MhvscL0VyY7PDT
Gs33ENQwjgVHwIAt1vAWc9DKxcj6a0nCos7ol9ZeFHVrX5uWCQwks5UJRBrt7dSyZ9mFoH4kY3Qo
bYDfP+qNwkXmfCgAOOv8yEe1yTTL1M9nzmc1YRVLkKQAhLbpPajEMMQ3J9m7usTj0W6ayWE5usdL
pSHr643D8SOvJzZysk6wooIyARa6ysC2uMC98/UX3YfTnLG747+Xz7Lv+EwvIoNbYp4UEN7WXTcX
SQrt6GN49sxeTGO7KBPXdHwT/SKHLMfBTmpAxpgd05/b7xPr3gjxtPjtRMCJIp3+qvPsrA0UO46G
zJ6Y2nkFqh9QAfUfQwqtPMx7MuzaJpOgtPB2FUM7mhosvhBuuPtd4U9K4U/aYZf0VxtmHyzi2PtI
WlFCy0kqzhq7hbKVwcQ0IYwBiWTXKcptZyb/Z3pAXmKlNhvSLzOwVarXU3mMkqwoYebklyMfu4Ct
Op7n7hfaiplfZj9aBDj+ex5G0/B1Sfzmh275I6v0MXvAWyJtGKFdqY9q3J5HN0EW4S8XcmzwTrAJ
Kj0bIUyqUI2B2lygTw4O7JZysFFvEP9HEP4svB7iuewkFAQtih/YmGyyekVpeTZSCeT6xGTnNJDA
apFNrlYthYcdNzIWL9L0pVYg5OUmOfwWCo1MjBmyiZIECQvMOLCbC2Gt8ZOfRabmIQzPbPo9oeWe
lAWINDLYox2SdzuGtr5G8Eacnar5RNiEJVh9D9fkb2G6OCj1YUh8ly9TzNBNlL4d5Z4tBjins1dd
6urVLpXCxX2rY/5FPHIbkrJHvvgwRhPxc7U1/CyrXbtNiXgGpL/Wzmwx/AEDGLMQty1qd/Yd/3KN
yHzSW0q493g++hQOFLsP7nAaXctklhwkv8tv9K9A2e0546xT8+xOacounxCLPYyqNiO/HoOd+wBu
l6DcrTywmIrlfvJMLd10+jIHRnADyoi6ZImiMOZt6Sueh7l+XQK6G2lo0hWVBpW0JdU7VO84oBGh
K7f6IZFC7mNLOVmctTKoa/wZmpWBuExppk9yyD9IywQRPVI1deQ3P+CvO8xDO2hzAPKP0DbQ9eH8
MWbS2vaMLLKNaEK14mziLSBuzOCYzZTwyBXOfhqm+zqva506IFQD6Fs/o0eCq3x+sp+pXdpKY9ro
nwLDfaoaSQc3RazUBxPxhwfXVWwglvI0WfywPd1zgNFHwQwpGSurQk5WYThOHFSHAZvZTyv/NyGT
54uOKhKd33sY4Ym0WHL3mKjXFR0TU2Cd8qBLftKpUpx7RgMUNwg16WdjSRc5vgQzvgXXfC7Mty9N
zZA25dN8+mb+rMhbk/sbPMhorsTOg+p0fLjEdxq358HIYAdmayhRAJk/o4vdkoo06U53kSoq8Ctq
pbrxpeX0AE+DrI1/478sUqtXADFtsIZeK7TDn0wCpsG3K5RkmnqUySxUteBu4R011mWQf9YVLdcM
FoTwJUGi4ojIe7r24ujuj0kJSoR6u3NB59nKUMXG8K+veNoEsexaUobWE1AMdcb7KJjlv7MnGlGn
NbZdX5bsWM1KnyS5pCMReNNQ1s2aYxup6P3RxcUcw/+09b9FC0oqmNzgoGr9hKlYX26wX0vEbkAs
HhXDZD3aMql8klaMRge4vel9G1HEnzS+bZx9gkXwq72X2+MGQT0f+gP7+C3ZoUZuuMDqi0NUqGHw
hEjt4ZYPc9D3r3OZjpQ9801fFzOk1wPn5I8y2fxM/Yvwi+eFPTR19WzRJVOyoRPue6xoGsW7x6wI
a3sa41crtqqBf6oIaZFDjY3a2wkrNKPoh9MAl7dpvwIyZ687lZ2pnYvVZxiF8Lyh43wH5NDrnYPc
0DbFwA63ro1zcBpAh3p237Oi/Xzy+3BgsxZfgRSSZVFMIOira4JyQ7FQGFJ8XiYVCngTu9nutCdC
itKBu2/Y7srHrDRC1Q2T17fOogwuHMNAs6kj7/L91Pq1gQO9e2vQNA16tIYsmDhTVZH+lIMEKgdH
gdk/p9Vnauqwc63Gnqaz+6UPMcqzlSf5v9sMq3FESpT76Sh1RIVsPhaQJx38rEMVZD+3R/Tcl64/
b31RXc06QheeYg7pW+pNrU3KBHIXqW2ukWLFDqwst1/SdzfEeUL4kBN6x+ZpftxC1+lfhE2APU79
fCi4qoHXVjpiwLQ85Hjg3wVumL/78pWrE/iO0RzXvahBfJdq2sXfg8Eyryjo9LRwRV37MvgNtp1U
wp/UIYZ7tVo12lnRz9aOkiOJ0sc5jkO4EbjTJS5jiYNhDyuGNVeGve3CoYH7rj+EdNch+MQb0PPl
tcf0OWaI7L0ccFGyeOA6xJysPpcBeDVdJK50OMrki2Iec8NJ5GJyTo7civMStj20+3DvBy+toDbq
FPFVV+OIZh3e4pSpt6H3IyGYUmMosqUfzid+TlkLF324LKTa8XCxghjNgHlTIe5NWNRFmdx4+ms+
mGZ9K0bvxduB8PUef27POw+T0gn6Ey/Qv/mXdgrLlwEjjV3bmSkM25sbqkk6KzUBNXcU7L/Mobep
a0F54tig2znLPvxi+Z/25mLrVWXquT5HPCCKjpdoOi4xjU2gShmtb7QARYDyYix5Bst1tQI5gWng
8UBiQJpZqTbLsfPpz9MdfgFFy/K8vQjDmJWSc2XPFAsMSASaNNP0ineo03ePq+tDkj1sZzU4XrLk
kGRFfRRiXwYckcJAJd9wSylg6DRcB8l8M828MRhMHoi1Ahpc/m07hLcAWwDDM+/kiVEWZa3Sz5aW
if7dJpLR+fMsDTQcUdd/TS/VrB+n8tRfEZc+oR81TjpdE4vGVTggh/Zvr5YTbjwt1ARglxMN1A78
qnrwQdJCGhBcTeOOPMsgmmwbdcLNqr5FhNPWn3dsSOnui94wHnat3Wzqc4iQPt4QOj2GWKeEpt0q
xslDGhfNSwdiNGHQCUtEI4JHlq956i5aEN1r25c0yNzbOb/DiROaqxYyLZA+Ch1Wwaf38xj7GsTH
ZgDBAkmNQaiVl2Mm14VlhlPjeSz4n4yKqVSG2/lA9tIxB9uIqlo7PnSdOTMwiD8JkJQ6uVaAjUO1
0FT00iFXxHnoaaIO57FgXDKBb+q+Z8lK/d3pMYK6OlL1als4u7tfCvoz8eljQvraGY+eySTYvwux
W3fpsFykiEx23wFyV8gz/STwcG9OJzlHmBZgLVf1TOvLuNNM5feCM2qCz0Yr8jH+XDYaw1M7qbsn
IAEIJaYgupE5P9Z5t7d0FYlEwuDYh0GJvy/AaA9GjQTqQjZPA2MKttdexELdXkii233FKhmkHnZS
znRCt5YyEnDul3bw6Qxm9B57y9HWgMUukM8zWQkFELJeZ5D9NeHRojyFOjtz8Nw26t1w7gr1Yh7C
xw0YmVmKJrHiG14ha2K0eQYDgprc4qNEoiX4AW0omdP/L8RMwCOKS1VfzLb8qkrieMmw14l3FVCo
Bq7pAc2PF6dO+ZFsOXTz289MUbzLKFP8YwQbpU9wAb9iTti3cZ49it0Fpj0fb4AemsK8B5g1g/LI
WWXCPwIiaru/Up3u4FhxmBCTfojbZy15eAFsgupZeKXea2rW+WCm5m9s6gO42dmKQ226vxT8Un+o
jBgGhU0T7mDQ/1wUgtNHvCYcb9ecw61aqcK+MClAsA8B64ovfT3YMG5yBOSHzrv8h0uJEPxxV41M
03ba/TDk3i59LmAe3g73mBaxXWO4h6Ey0mKi5KD5ohWbh9CGTo08iEnSf6N/vGEQUaImqTBuW3K0
oiSU4KNw1fhBCVRcAS1Wj+4CeNWpT6uHqJjbWFEBUFDE+GRY1MJmNjKFc3CrNVjjwmcVpAZWS4RC
mEHN7ydGxy9jGcyaEjbyLRNTti6YPaBXX/Bi0rsHg7X+JEFJRjY8pLUBdILrG5MzezFgYED5GK/v
ilNOH+mXHBCF1umN+/RreBjItrhPq1iwvJ30K9L2E28RXCsCmDOzukK22rVxhaeEI0kSmVOU56BE
PPhOKD97xPgkMI0FS7TuVe5RRg8bp9maTg2pXPcTR886RzfoTwM7WmCTs9tex5YKP3qymVr7wWcC
0MmOQy5f2Ac5vqXlHCWxb4KEBQwQlYn1e4LrwVcflq84POG3ZkKDzvHwc9sm9dkJbi2o4XpD76FN
MLyfaJWzXA/KSFJKiavmrtTc6PfKeiXRgNoxZoEsuuEhZqSL8g+FNDjRCQe8O7gq2IyUS88p8zYf
wqHzLUZ3PD9BuFT/YcB/1Zxz3KVxCp00wIEAkpxz+iVwd3KG1n5puQLRa32rviIbdmBWI00Umz14
lyMwvN4EW3u34tx2KWiBcFAQAjYs0z1pKgQBfVhOv5hLn2daQYM54/cB1XQAZNyLLBBV4vYDIC6+
t6OwJNr/o8rS5ZaiRlsRXF7p78XwvGbVNdlZFCwNBj9TLkIXhn8wbvaeqd3cZQFOGpbX+3T81zfm
pSMrGf4twXJzVObj+pYGQbHGNsM6FdKu9P5+Lan5VkEFfWX4ct2v0krWHCnVsGnDg8Kh8iByQhrc
wpk/cyZJnzEHw/nSJB2OuCUnGfzNieEESnmrmmo52LzwYfC9V97U0kSBaYRWvXSkKZ2x/Bokfqf9
5iAQ5faJxfRTpeu7ZOSJD7NZvdfc4y2yzkckH9LPK6pybIobOjf/oXh3PGB6vz2pUb0a1h4CvDYj
XLofffoUWDHf7y1EeK6/8DGBNP7PJh6hbli5e6G+ie563FI19MOsvabbMANoCYRBGhC2puoDcLEp
B38Ic2jETc5jKidY+9qg35UmrrkMQJMHC9OMvyFibJ0zunOwInOg82xUnGcMZqg43wOLZXoeFuBc
cxgmB4T2nzfCgTvPmleLDhBjtEn3qbApurmUywax8rG92jbKPhgfXT9zAqGraihzGfG//FJQFmZW
pL4NO7Ovp8eF6gPC2HRWKRvvD72iuMx/J1SZlDEI0P6cyIDbwcsjredFCuzGAgguXqBGpqOa6vW2
bM9A10iJfHhfpLg6EED5oB0/fSsbT2nKYVBfQOOyZ4DPYZ1NnXMoPc9jPMTcOKKEpbtw08JuODX9
ADi7wLnkYsqmr5rO2NrtwgKG8rWwVJ5tGq6X3mHkhQqd5ebqa3HTMw2xsye9OeTMSIGn3fsVHcnK
F8m3XPwahjum4JNrI+kv8R/m115hMhJPYecA3VJWjVBcGJweDdy8khZSYbcwjU4JoWPQSISB41TL
9Hs5T6NETOyzbRHN48WuzzXDXtW/3kZ0aZfCVFoYuM5H39RIcZMCarWFAcb12DcQVL6LASag+8YM
/WCUkRJrx9T7rZNRDv0r0Pl+/JIFuzWZXDzJsVizXD8S7DtTGj0nIwv6VCG0fFXKrWOuONdG1Hfe
gElWlQ7uaQKQ+eyGGDpGUBFqb/tM7Txw1bCo7Gmv+OaO074hedBIVZ2M7EPmUdG5zY8yx+Ex3mK7
9JwF7RUnZ5YmiXh8LPad8w8UxYxeaTjJgSC/P9xqzpb7/8bNtJH9sgsnmquFSpGFS/we2edVkhK1
f2dmcxMHWwP6nBqngWNQI6vpJquVl/fL6Vz9N/mrTY45AXKZVK12duDEF+9C0epB986dBisLNka6
wr+h/H6ef93+sMQHCtXVu859pMZs655me0gQ4Ecw5wu6O+EwEqxq8T0kCPAzXtpLSosWmprfBQ5k
c6JZnEKHBBO5ZKQLoqYTy2oLerYlU8JFdrzYrQCGNoieh9+FA/NMUvywV/Ic0+9+jEK9oPYV6dv6
WH9hEsd3U7WPVOE7xv0SBo+g3o0yidksRZrCu/28gA9zM7nH4X9wCIeK6WSPgRwXoGsFHaiWti0b
DP77Z2FMy7wHIbl0pxlDbevl8S4jnFotj0Hkqy6i2QQzbsmiSTw/rLfHJC6WdxtVK+tg6gPI1vvh
NBMcsCSurDvRF6Ku2b118mqz+2Wbt0yLSqsAv+0g6Bdr5X918hpxjl+R7kRbliIJ5Mi5hO41xYL3
0OtuSBCrUFelyuCfXdg8nOcWA9GNAsbQ+cpM9Cz8aqvKXa6RKyae6nep90awFKqRMC27B69118Aq
lN+eicFFj472rZDqxcLCYFUuakbpGt2Gdsh+rdtaAg4dvYCSpa2RCTaDoa9qWvjxxVr23g0q7RqM
DBQHTnuUs0xbBwg3dmEjimmOQExh0aqgWVf1sl6I87hH/RFNo3xNiCDkL/jjq2vVPC6aWVS9W8I9
6odiNvTRUoyFVLAlaUjyC3Wsdz8/zaFF+siB7vN4wKlZHWsesfcgQ31bYf7pEcbk/8MtaxRtIe+N
1TuIh2E6IJBrFQzJio9vHPHeyG0S0JnTqZ9ZSILy0ycrtGUNZEs/IzFlDGdkOPUXZCuczbbEmOwY
9PPhu9TOsfCGkACVUve5jiwuejlSvKV5MMg2C4VZYHgGd97WNFdv4YLzftxLWH3MAk0JpmdSVYO7
rWMkqbgROxzSjq4Ymn4blifGsJgCoZ6LOni667ri/+uAog1w5nJMruryIAKxwa3TCvxf/am7jgKA
0zMehQiyDRAhAO9Qu2zfjm/qUBEYOsUuFcRZ7pLmTUuSHA3VNONCbtUdN/Z9+zG+BopN+s7BedvK
q8WI8kY3FX1RpH6bKnnjqOJdvW5ELNFLtpJMVB512g4PYvd+fxEFmRXwU2+L1GtA391Dn2sUItXF
dolQ1PFgnsBiMxvwOcOQBlRiLtcxbxPt3O4C3mW0SUqfbhEGThTlBNctu2EEFeNLgRGoa1ExUOyi
Jd4mJDa2IUgma7VRZhwlJ1anXUis7n61hwItNcp+0xUQAK2GbSMakQmQlz4REVP23agMQnUtR4XX
sSQFgyq+U/PYIweQ5hA8k2uX7hTMcI1KDFX4XudtbHaOoyDe3yPZGoial7MWPRqIimcj787AN/sQ
9vy5Z1LVtq6lUuzAacG+VbKT54Wsoq7g7E+O/ISHGZBDWmXDI9MvtM6RvSa6sib7Tw7KPBZlmSBN
ZicXf2vMY4c4py1k3zMLUSQ74cUXpFDhB5AsOmdBGVL89abO1WppTxsvi71LrpSG4RqgVm9aJc9l
ooBDDu9WdBGE/jV/88z9GMPf+/lIAm7+a1TVl6v7veQMb162TFGdMXFyZqCqrd172eo5E7L0soas
UcOeqHwNSbdT/9UQiSubls1a5Q1hAe1wc1OMLuoowCGJfsSDTXZ/i3Kr1zR0L/kuyo9WqvJCTFkx
qjtIJLutn5SQvd+S8MD9Y42OMVwSyd7GXLvn2gZvL9KlVCWmzAqCj/VMKcRmzhz6Xo0bpS3MkuYp
UobWHf2lz6Kp/ZEzD8sJfF3BeEJH+VmZq/B4/WgrynzoH+iUB6Llzw6LALpwShG21/UVgZ9ZvYru
bqBCubr0fErNR/sW1mwnq5tl3MIcs+Ht+EGFvjrWGnZoLNGgVyh5FQsUwxGuBSgSYR9b84AiWYTC
K9m3wYpr5y/ZIqGPk0xW3C/F+/mzNJxNR4io77lWRe3SV3eyxY0k882OvCQmQ3UfEUBPZNZOVQ/5
7zbnSFIrfm8P2HiZNwkuZsKdNczTAnh/Q5c3ffozvWPR500PVd4W+qf6jBut3NFZWpfXKqeMHvqo
gHlLApm870kN/lRqoHs49EbFaNpJuTuxGfLGs5OCO6dWIiGtoYRheYnodQlx2iiyw/e6dAj7oZSW
7hQS+DtCTepaSayvG4kPjdXqUK5ZXs1wNFKW6TNiosk3Au3lnyTmeAb3/jAlXUIZKGgxB6bvGedC
/i+ygFhhvsWhuU9ul8QWYynALMcKASlfj8tO9DRhgMNSvoB9NjXRFq6zpDWGF+pspjeVl3s72/o3
XlY0Rc0tERNMj6DdmYFshqjHLFkm9gi97jUl4saMSJr3H+0QQhuJGI2wHwjprREByRbJtx0hSHGy
4DwBoQhnpTeMF5CZ+hlkwAxNI1u5gGyCc0mg8SUTnYWtml8rguUlAPfTTAEJTrsb4sQ4vfpsedPc
0JcihraJkBorSvaRZgP56HDHJ8NqmIKNE7t1T23rBB0n/MUhfvsQ5KkZT/ezbrR7hWuVajDikts2
aODYl/zVW49xEHxIqyGpkFuDmrq0LIL1LLANT0m5Gfrq/uDkWY9ZbZHZKwB0eLVJr00z1EqTYaXV
zyeDNsHGaWIKYZfHz/5iIQlSTpazu/WfRTqNpv4F2/U/D7VI5yKYEHNrci0XJ2HGdSqtH28udsiy
0fM766XrxVin1uGlJM+l7qBxS+WfiyeSEd7Cw7P5+8Dc0wmoK7Y0+M+c6zyJDHpQNZneGzwEyI90
uyo5BShaX7VP+/iD6qIOeJUAn8btTt2BeQlgV5vnRha9SN4QMixh8g/3hAtYDAsuI7OlcJ3StoER
4dNjfumdkr5RpTkaWTZEkWJeS0CbAHKTIl7kfH3W3oMHuegzUtF4Le6o0e1z0zuDB7Aa/5vtvTKY
UIx/bsTmXVP6m6XytF0dcmfTAPtlcrmp5sa3uEPB4W97QTY4u2dWxDT8qvW0Jeyp2zK9NzvTl+nz
qQe8D3AKRFmPsXwyGKvobUqZCxdPGk4qb9yD9tp7bpV+cORMltqU1LONVIN2kiJ63CrZid0E7LOS
HNNbzHhdCo0uIZAZFpD32yrPHWhBtU/klKlvPIBB9qULZPezlt9j0rvuYJBwzHIV60GFWzsztxXQ
330R85957CVxjK6Tyj8lwGVzKe0Iws54SXo0znCkO+7RRoW1SeUl/gDpKwuoqjMx26P/O/RtBdJx
sqZmbiDqJGaA4LRZ0f1wTTDDt5ZAHKEzg4m/RX8a7Xzc/hlsm2RsK7BgDZgh5jx2mCakXBIIraPi
VH+dUaCJV2s5fYjDVEJh9YeRAl+a5SINoa9I7wlNd68K4Lyjkt3tYx5/9kQwEZTokxz0/9Phi/1G
ymKIT1/Pj4CYDMHuYWwJzVmMzxgSNov+TBKGQtq+SU6tGpKnKJUMxCDHLQYiSIRTxKkyowTjbPUN
7lVKi5D8cYgrq4IufoqG1fwB8gTuJh2loSmdvZOFHK6YP2j81QBTrXRysmxkjf8yyc3MeXQBbXhX
OYSGyQjEp41J9ZsWDzINQE18YD5PSPdkvNs5T6A8czRA5JNb8lSZUxjYwa+9PFf689dFE4x0un4q
rGO571PY8iPaTmVzyyhMRteednSJnlpADt/30+VOXSFqsbdDWYSNc8ThNWjxvv0WhQVKQArgcY+q
TNWqfB0bUEsHycfgEg2cxHz1OsFxFLh5ZlthCUA7lKtscXE9LDLVP0c8x7QgvhDKVoWzlhbfsu+P
1/mRcIDh5p4I45RdAynTPaVRMONjASOc+0jL+gzGPRfyBOD6/OQlXR42H6xTyrnH3CvDXBoWZgRw
GA3TT76Hu96XwqTohuxC+7oqfFnsNCS3wmKYl+SOuLA7bRKwoLZ7YSwNfoeIbjgbe9/VVAUc/+4S
0J7Zxf9d0kJHueVM7+j7UD2CG7ltB77ebeQcFVKsWNmfJzEd92NYZ2iXprsyBjvGyv/BmWoSmWaf
KsJxfbCN7Vg0VwOwQp0A7OS3PvzUXDFk9kKsiM0lrhADE5KG0W3iu/Seldr6VjOxlBBQpIeQwyZQ
IkpHNbYZrQk6GLEXd27sVWWHDBUTNrUA3TT/D6GlpH9lzXxNzz/4E0W3gS+YqTHaco17t7UQ8cSu
eB5igxsLVd1iYXs9wtraiuMKo2eRwgUV8c8SLfpWoYaOfZYApp1clRNMWEzp5hW8+Yd4ZPDKx547
nG/MhmOpJh05QLKD8AwmcMGUQNIeQ4ay1fEVTDCTUByDSYtOrfLnnJJQqOnSGH08fma3FHKU/fx5
OrPxiW6DWuwREU6kPhnF7PmDrYveBBHnrP/zaE2RCwucYzJF4Bx3qfAVeYSKDoa3XjI2kQo24YJs
tGU+rGENuYzDyAWfGcndwg5QM+8FA23iXot2d0qW3SGB7q7gdAxUGoyrDCXp821HYoR+dsP8m7vq
8cWTBLwuvNvcJ8B/ZEGsgUOpvG1ME10J9PmKoYhIvSiW4JdkBCtlPSbWEFJ37kLpy1fPeWi14/f4
z923W1jMzKxJLzH/6cHVTyaeoa5sBm4XGGBhM+DMSg//cdE2Iil78HtetKEG977voE3reSjaCMW3
K4QNwBWoehGhEACV+SvzfGDUMjRl9hRYwxPWmCN9iE+ivcI/Y80cpRlZVLzG3jB4n9izXw0WBDXq
/pO91rsNeUMcZh2S0Hgw6Sl3ykNiaGeoLNyrE1k47qyN0CPtYmhoENS6ntTpVxn+k7f6rrgV+SKz
puZ/5FE/IkbUsSdVXwbjHiHezGMk/iXlX61E6xL/Hp0lmPZ30Qo5Cm5HQzyJS4ExjRglsWtEpIHj
M19+uw9WpYZbLNdNxQSjlTJ0momjO9FsMijX4xA/TEJqIPw1T17pXP/zHRPFDlX+atC81+Abx9+9
vRuCQu1VBWt+zKCMV+LdMgivMwaoSpgtRYqPGvYFK4XS4Th02RUZcAnxVuYpNrzO6yKWhG+uBXBo
R6LAeKs72ZVKPzVSSproYEO6BHDgbxWy2dCP5jC8Nua5QF19IET9BL84CmSjb2s5F44x6JlNR9Wy
KEFua6UQIvCDTVn2nFIpTezk0HsparHyL4P9Na0kMIFuNETvLndY3+RVIs7k4k43FJ43rRWafNsB
Q7nbzzFwVTemrylEju3IW78SAH/it4JurpZhVz4q1dOaw051IOAF2vKSg6tXGx1rGnwUfGw1vcTa
cLrR9DPnb96V5OOHfFR/Q6cMnatrCndKIjon5pG/0u3AdF9EXzMSBqi5J4vCf4Znq/UFtwukPppp
9K/JoblgYJ/UJRh5qxAn+oAijlVFubvH8Ms5R0ieN/Zz2Tl3KRgPqPzYCWDkOsrVQtR3akZ9xuH0
kFPsRps5pp4AqYcQ/Cuu9frLvma97iOU0wIB4N4dPGMSGY5eLxhao7Da/nBzv8cJYdxiTX4agt9b
Gq7jIajaaTgcbs9PGuT0/3aaGrIvxaL7Mn9iS37hqqgHUYZQ9K1kC03duRcpeSsnS7I0sRhULR9b
ezPoK3z+8RoEcbDsEgu7BrtbRaGtz7LN2Xogk4d0oVc+vsXMwXgvyTYh8B5p/j/WbFYOmh6xmeNh
4Gljn/2AQuMV7phaHRKgvmle4Xb2ldd37vC2xiCqT2jpIfvilDRpj3yMsgbIUTk5vGdRcvxhNnvf
JNV4EbFgnjK+T7/PC7g0bidyHLq/Euow8AKe+wpwLVh9Vah8V6AybW+qgr9pH4g8y+CSTnoGpVIz
8IxzeXuZZ1h3b+ahFBzq5Xu21md8rDas9idXOTn+Rznb5vjkJekL4dbyg9UbuoDf3Cx+w5Qrfdrm
XbuwBPNav9rLnkIs6jfZyvOxDOJ9p9B9hO7xZLdSBUrlAwwr/SSZD3PshAPYn93SfbK4ky/NSyGe
yNfoTFoYEfKumFUDwPtetnOa5yFSACvSXXUDZim9/Sc/ioPaJvNKOYZhnARAN8zQxNT4wGcHFmUS
HzMXcFu9rUPKvJMIn27aBX9BGcpWv/bLGCt5kCnQl/qLl+Ypl2rhY+Iy5F4GFVh5wuRYiKaptV/o
bWh8m5M3gYr7pLMJ/YxYEdRZRJ74VyGR+wZDLiklIirIdt38Q9sWqU2bzBSXRmfZzepzQLG8PjSo
7XWnZtpWX4KlFzFNQSy47YISN9XvRS/1/lZYizbmOZfyJ2UqVVokrNgiLPoybbGt+Iowr38J8QEz
PMhs/8FsP2OfUGIWb37zMHjxj262DP0nIi5OR1ycrEqX8qiEgs2P2C4pZrFu8b8zvW9y+9IqogwP
r6pdipoJPj1dm+N2kiI1a0tJtFeOy6eGNmmK6YjjLiyXG3G04u7ubRLke/OFSAcPxTKsn7OQb2JS
CoX34fbZzM+/pofeRxQfliNu2xZa/zDOgpIzxRuyNPrItdTBPCP+avwbI00HUOgq7VEMlaE+JVqJ
oMWtposQnVZHnImBtVZCidsBOL8XOqF43WwXKsAwEd3sA+KN3rDVj8o9JSh0VRXfKOPGUNZlTecl
84SG9SNA/wJBCxGghDH2rxKmyQHupqnpptJAID3hCTDT3lNCbLzFQX8DV2Lag9G03I61xcBSo7mU
kiXCYN1j8qWGLgZ95iN0liLVJolibakV2rMgQelmPS7dffFtSri0psEvdnzGW1OFmHAMf8Z/zBpp
88TEgf8Xg9TSJDtCCGxXDxFJh6aQi1vYitC9f/ooEpvNMiT3U5NSGKBbeNwnTtpuH1PL/pxgOWXX
pDFXprrYYJSPVUxx6qLXCHtxs+MsnUsRZJ2zf2nwrFqqVSk2EgODa+JEmlCIZpn1RyulN51y/dst
tt0bS+t7qw8JBEN1+0e/2CLAZ99V32+wj5sYEWFTiv58NcS+64txam9nafbSOlW8mx0V7cajcR1w
6CPdU7YhNxJCgo7gOepKT6q/xfGEYFHiLKQ0ShYsI8qPaXO1xsqLP+Z0msl8WG7HWlXOQLNEKYJ1
kDc7BqpTD+vm00lWP/7wN8N2jkTCw4MlVEAI5hwPS6FinKkry7STvaUyDKEisq1d05M621hQTh3G
T3oVuEPDygH2JUC2txm3pOrD8ItSpr+8/MTsOxkdN5vE11pZkpmX1wFc2XgcXxaqqOrT8vQyLrcd
nYzDMIOnA8qQpUgm3VRiTRH9Cx17ftfp7LbWGdZoYPg/TQzFSo3xNKBFnPiuMZJF9jd20tKRB1hR
EfdWY4bqw+1P57chjAYElhLX+81EVa5Zu4v+dFCSMeS4Uo8pomUzgmUbLjA/RWo4+9qIBNIonks7
Y79WOwmwsEupNxKfejACkKDxp/e+ZwUQaI3oOEkAsgqchBcxIk1pKP4AUD+Uz6Z6y5W4zYDSKS8j
IbnSp/MoawX73t67yvozkucooC9AXzMBzYzlZY0oHSP7IOh/Ya7MBUGnRpFEOK/dwPDXiQfenJS1
9e+XwkKpkMI9Zqn1JpbgfxTxoN2EnZ9d29pOQaJu6w1K+zDWhRAZYmFTm2u+7vg8sWWLkLRQ5Eoj
t2yPVVGqw4J4nkuwd5NYd0XLmRZ3O1kg3/G3k3LxKgyweieq7Cn7E+2Y9bTHs1kMilpegPuME/yI
VqjzvDn7zwVpuN5XY1fCtP7MSnXcuKyEbXMyBdDc1haqVRJXM8hXvAfpyixKdCQBeD5cYLsfJF1R
M51StBrgrF1geWOWI+1MPkTmauzO8r5zJHLUkuml0mwD71oZ4CpKphjp+srpmz/k7J0+O63P4J3s
d4etoPZ7xeV2G3olpL5bgpYRqmpHQovamCuRCK2OtSF7o9KFL/blslfbBMt8NiYPm+TnLc9Jqdza
FB6cRLZoo3iDSb3g86I1FtNgIH5DQGIYjkbBCPqlN4FyPi0IDVhSWgd6tr8nU6cAvT61ZGp9vv1P
i7TWxScezmZBEcQqowOS+eZX+rbPJPdMvrzHH0NQaEEiXRq+S2Q/OGc+jvUXdtQX8CRqVSa+Ou6k
nZ5Y0xpxpJbvJVJVzWtJQkvnwUUMLcpm84JhzzG+DS5DVsirXLjot8mnlz0i7JP6geYm4mpjoKIT
gOdL0dbEZgQFf0+dPfrUkQ0k9stvctvMlqR2TM9C+Yh9pgK1RnQfn5BdvCX/c5nbQP+xYN2/o0Uk
rZu9RUL4JaRdotekFxluyKrc+1Np306qrO/wC8jbCaPbgA4ktLy/2pVN6zZ8mhvrFOCcmoe8GR/B
/Td6wJYH3ETHaWL3qgQB1yfQ8qESY/iJ3xIN43CiPJnqssnpGePCa/C3/mtv5QR5nnLujaAlANN9
pqxX2fQLhf5CqdBkEKZQy+ZxqDLBBc7yX+0gdTGuLGlVHJId0gDz2s7Y21uWLnjh3G3NIFhVm16A
Hs8F8J45q9WgvKFkitclRncktzuOWjnORWGVBCUdYPnAPbV0+4ST1iW9ypwZqk7hktTI6wxj76GE
ftTT1W+nWn3eaWjaBSsVsly7OavRt0+8UmCt/wIZV+udgUv5xI1thQkXtS5P7RVXE2ZN7SgAnLRv
GJJuHy5nfDUnQvnuXBdjREGxC5Ij9Qk+vHapr/wZfLn58fIbDKTNNtNp3ifG1Rqc2Tv7EXYKBw8D
cLs80V6eiUoZRtM/D6kdeqLNZWzyYCQlz32S8us3CVgudMvduFZRdDMymDhwdKHonh1+tzf5p6aM
4gPWIQJgaeifRwQr0UzsPdSryMEmuLsHHiMmMD9sDac5hTDWvT0ENR6PiC5y0+1Wf3mJ7fpNdA9F
dTAKqGWST9sluZc/NVGHGVn86twc4C9NTQQgYL1HVCJbfbCJsoyfY0avGDY95LXLvmiYM3Q3bXNO
Mcw8nEbm48cs+ZvHLPpxmUcq4j6ko4RpjuPZaZ74EDng1LkxNpDllepV0D4MeLM5dPqUPFMZI6Jx
t7ziJJtIkrLFrQ2bdNKcSHfPPSnE76dYGFzFw0VK1zbyhTXMYwmvXySHMlb48oYAQyL56NmyOu8O
mIX0p3LAvXmScdr5B6GrPsfuP+bxFO2H94xHTDEGBuHfnkI921kCLcX8pIIchH/loJc9fP7paOhS
H3ehuAmJiWBJoqBGR/0fEW6onSkgYQf+H7DPr07q69CCEb6IDB0pzIy3A47PMfuEG/Uz3MMjxy2A
CewYMSjL488/wTi8UottaZuQCxvsKbyMmzPx2xxtfCgL30peDLxhJ5FuZk/6VjZa3Xd2IwULgm0w
hLA0HvyoZ5nVoIjy4OU82Av0jgF2lqsNIjyqbUAM7B11Ir7cVMse/z8kbdpg2CbXE8BJYs2I08AO
VUwdej3MtoHJd8nEdOxxlnhnRTrj5AEvj2FV+j8jx+eNPtXOL50By8H5Dmm1xBHYsE+2JycatiEt
Z2mE4tloeN1N5tlkJYb7NnBdsuWZqxfY8mG78enljhx6AEPYW1gZB8u43P6lZgVL9DzQrG5/Toox
54cmT8Lyqa4AyjwnL3TBEO7ogsn9LfB6RqaAOHiq/A8KDwwhamAXxR5uYDwvz2VjuZUDhrm50N4p
p9Ho2CQviJxKYb96t+H8gwbQrEBEn8PN7YGl+NFQXqvY1y7WHK/JZ4DJqnk5E5UNEIl9tbnd5uOG
1pjHH6uy8oL7bwisXE9HQwElf2bshe8QJIk0mkt23NNoZr+3+YnPBCn7otOptEHWITcKnFP8I9zr
KaIiUgYAsoe2/L2xDSPyRymkOu7NveKB2blaR6aOVdjxRZtvPyZopnqdBGAztIqWQEFG9V63g8Fp
fChacfFFiOlP7iCZq5BI76UMxYZaWEOyb5h0tOFPBPKom2EZ1RaqY47BVjpAwGdJEVLnd31JX3LR
0U+PkLadV0OdmNHNYiaZB7EaSrtNbqi/zvt3HQN0grz5JTlZtxS5kpxLsHPOC3ESIL9/h2jhq9nC
LWmJgZaSeopjbYDU/bTAjNc//xf3sAse/xurNQBb52Qmb/bI+ex0CuT9nFBcKfOzvAR6JrXBtb3/
AGZyX7k/RSgdRa74JeNs1CuztgVCol3LzroD+UaS9Koym2On/zulXcnc5Hq5jbefkt62P58Zf8Cm
fauZnXG53CmCR2P0Zwc1yTw38xu3tmqdMBwSxJvbnPEP6d/AOaVDfZNI6iw906fzZdIUhyFV+1rU
VTM3fSITl1DPwDw39JxLq38TiHxZ27JGHoEh8KuJ+/msbE/xgtM71pN82NtZOcNpH+3E2Larc3JF
V8BJ338dnmQbVO++hSysi/VKIQV3W4JGNCFn0YO0ghFgACh2oMJ4MfHcfaH+wo4fRqkK6HLIF3s7
MdNN+AHXjZM/jjlfro4OMYKutOfejpDpf+U67g8+feHPPviwUQ7BmkWxkdjYQFR/60ZZRdtZYEo2
ht+xDWBonm5evAAGo1SMVxkluBQ7HF4mRoP+DYAKvRV4FXxhHvmDFDZae9atYzQPoKMqbCI3Ds8R
LHOcfY4ZOFSzRxZGHBF8TaaaLAy4W4wBucApZYqoJm9o6KsZl4iiGG5RLekxbxlV8NeOaYsrFae2
PNdPbDCahuPnMwG64wMetJmqZrrtkf78+qp9uAMVpmtF4a6zxeAC/VAgb7cb9acEeaiTQ9lYtGKA
wJ3T4nqhf67lYi444slywvZbzHgGeiS70Y1soM5qsRxOzvetC/zpTeW8ER9AlsCFWuLzTRlON3d1
yyM+8/sizp6EVzAkJv0KQcOk8MVPLXzp05BvCab3vLAPqe1Gy8YHHzSEL59hIOUHasOOQ8G5F07f
hrq0/XAMqIktCcMp0tg6ORM4uLKT6nki/omy4CzAl6DeaisK1wzOzJOTMby6B6ARqCKOlCcIhU70
EkqpkgUttgj9H8zav5iA/h6PJ0sDWEib7Lxgi52A+sAs8dcOeWBbwuILCeToxLVEG591e7oKBaB5
nskL4EMrZjN4Gszt/lMommWP/9siPjFWGelPzEIjojbhwUgYVgeOCWQBZ4wumtDefu01iQMJDm/H
CxCBneYeGd4FdBSm31cOClxXKL6oL/P5vVuDi8jxGqgnaETh2jIXXQR4zndGCztVsEBkG93V6jIp
FL0N9LOIeEvSRDYXW1IVNofasmUMztaTdPN//iTXH9yZo+U7Y59SXvQ/JCWte/GAU3J+wvG2Jpzy
KyoteRyk/9gKF9Lvy+VOfPiXhuy4NpbvJ1crDBXgG3tC20MICOeLEraoAdKmGg6s/aAN0c/3utEs
jNuEghw7PS3rFvg92yJuG9ols2xkfj0PWb5MzyCbYIQITugQVok2Txznnbvp4P5ApkqArKOZNR5A
YHqc43KL+0LK5VLv0IcbAyyjAot6YFn7hMhtafmC3HSRdamu3Ry//UiJ70cC/e+ucNzdc+5rfqvL
YSKRUU6gAZZsLxhE4tji+JLGmur7MXQRMQc/uHcAYatBvDnmzqbaGBrlnQh0Xuler4U4TAYv3GHM
uOhpeXZMqe1gQrGttzT/zwKrSAz5qcB+xzD3IJlxvuEtUTKihkCfto3yFpWBdlWBZ5HuUkJSd10D
duU6hjPift8Z+gTrHAiUv9HeAfds7gfP6vD+lLQrY7raVuoA8dDIc5zRlDP/MhapvNegu+jt0ERD
0EaXPhhgkjt3xa4INgmmmot7EXY4l3ehCz/54WqgWmPMbhkxBcVjtl4pbLPS8jPatqvJcW/Vqn3Z
jITyXv0D+zQ7kXw+zGWCqr9s9aoy6KPYesnIMROUWW7AsAF/0HEPbRqAMrKOfvXkaHla9jobUTXk
/Ltal22njsUWCn1SOkzFitmrpnpGlZIgLehfBegWxIGMrw6plIB6iyh39mjuEczzzxqGd71cyHCv
RXUdbrkgd6JLPCO2reCYIUdZIB8lmTFsa1MCBRkZkisDmXbbLuictmZcKHHDZUZnHnLQJAAJkq2o
BP4zxkycGhHuM5xmC9XZIuGbRiaW0JfLC49Hcz8o5sGobJFcrq4sFsk+cABFinnOipMIPUQYKklm
cD3SFUEfzVbEhOkd/WXHyfl6hGBUdmU4Xw+/uFoz249mzY5enLtNbvavjzK9By1Rn3N3NoebS0Om
tN0di1+AuT5bwhekQjjCCahAd2HZcQu/FbTJWOAbFYx++u4TuXsKmYm9+NMWKk8jDhGGOc5L4Bvt
6lDWTOoR15Uc49o/m+BJu5DygOFaMyF1ZxMv4wbBzzHN354PfRN4RHzcvUxtsvFTC/6SGRRvAKvo
UlnzIcia5vU9bYi1gwxr0NkmExumap3+NGZlX4TLt67/ORfuGInh3HQ6B86soOOrBr7m1JPlvkOh
GakHM008av23UmtvGXjT+Q1OIMkeG643qtNzPg10p1ahNEwVJgjl28i8cnw6cx0M6kYMJHVO6x2W
8gWD7r/CS2dTCvvSL9bEvNgxI4MT8qyQvAHoXk9wMQDx6SlMhP/vLzJImjPw/F/SqZjfX7GKbV59
Yryqdx0QJ1y+UdNtWtE2wo+xXx9ljwCF7pQVi9oy/W6M7gCVmV33zrdM4r42EY8c6Q9iLeNg/6qO
l0GUZ7ppDUvYNzstJZ9N3b+yh77rWmRgCExa1ndCnQKfrcBLO3qQw9Dg0rYvulCKD6h5FcS/4Kuk
v1DG71BnH2WFJc5nxbCam/TNkuPgnc1O23VbAIQVV5FnONYY4BBhGTqYXmvx8LhtKKFx/XNVvzPd
LMODEAjPBnxjO3P8CEqXMtPrIlDsJcOaIpImARyvQWz00njs45j3IKm5ecy5DMA8i6EaXSKYHjWF
uxIM0WSMpT4MDhaa9A3dhw1piFTjUiEyjuG8iKLKq/iWMy0pOS6Q5/OUVJi1fplzTG2BhHFzQDM9
Pnl/ap8JebvxceF/1nUsAt/tu+oprq8YqgPIpueYCKOaaH4W1rX1LagT3dil7gDr44VVEa9EzQBx
e3ii56EKzOWMNMFT79/0x4Jthu7KUIP6wiD8bRDHfpp7fg8Yi1PfJcoYvVui/MB9bTXUNJZiYfY2
nAujNpfczyWiZwOdq9j+W+F/NNCh2HCr8jiTwk3+Rcwt9hvHAU3t0H4Z3MKu7YnuXeyNR1NOzCSo
i4Q5/7t0waL0IwLcCzaFIs2DO8vFkO1zI1Or8Q3TtlURJ7oPzsmW5K+/husoN3ZSTz9Rj8BdPbeP
I72E/swa9CTg/lxUMWQAz5xj2T7GwDwzCpSO7ds9iSCjydhkZR9Tupqm5LG5xhE6T9/XrZ/UmUs8
K1jBZXkfPi8C+lrgRqGAzt34KhNJ48ComveeCWvgsDBCKR2fSx2dqNT3QsSAc07yO9v9YqahdX9P
wdZnvgohfuHAx3+MDKkkHkqxlns1nafpe1Se9uY39Mdu6F6uHKjHqXyXVfn3DRyRLt9SzsK//QDA
oltKro8fZcwvn/nHaJSU5P7tk7r1y2MFVioRjGwMMfIL1ynWKA/cNhgc4trsWMxMGNWwONAP2BBt
xTMw/E+5I7sTDkMeRfjYDWrSbDTVTIA4gCRlT9coLfSeEbPNbuOdeHCed7HJgGwW2cc54pHDPQz7
LkCOWvRnTUAejCN1ohkGaqDxvOaJiftbvRb3xCkYdH6mg1KDGfDLE9Ge5WR9AvP5LJFjfMkG1gNg
xhtQyxA2iviXzxPHeNgc2H5BLAOIcsemp/FUX8qSdzsRtOss2RFCDjEA4gZkUIAvG18SbbZSVe5O
YT0rcHtcV2wvwGPK8xRgBOh2Mbpwlwsbvtjjewj+cZRiBKpkFT3MUaryy9s4pytk7342nZ44nn0K
/DdX90YlvwoTQwmHHKwJwUT3D0o6Ys4ALV/vlWBkUe3M/0dkanZJrTsHnoHMbe5gv1QttroDmXFB
3pZVOWlX/d6OEJuNi6EBSfCbv4kpVCuop3GjbkzbPUoZXuugJqvDjiDtQdtiPfzyFBM0hnCvweBu
31oGhP/a0Lwygob2fe+kYr/8wKLxy/9PYeano4tUJQrUw4RDcuUJgp1wz9OQkiDOCN3R16Nz420T
CTtw6zs8k9iNoABCV6gwdKmYPlcCdV51G0bwtaJKKviWhN36f2a75I0nqvKHSvnKst6nvi3CsTUV
yEsXsRuW4zuvp0+rZhao/xJuIIMSkT31lFZh2zXNAnh5UvR5yFxbow48OGzQQJnbgWqdeGUbudKm
nzrVIOCuCKTJU8L6Zm5Dujg+7lgljnu4ZD6nnJNKzXMfe5tzZ7Nkxdpp4EcoLCFVe5kncGHqhdYW
XyTsqlbbB0298w6BpOxJ1CvynzPASRNgvavDETFZV7ZF+/Lx8HRjfMyt0feqFGKa7Yy9FwwVdJU8
9dxSL+lO2xoTHu0JFOMhhG55lwsvzcPBCA+xYcWLwrrC9mQaqRqYAcbEkVLW01ivbtuge0GfxbNQ
8B46aGdDQOg4k+tDF31+jaHSk88YaT1S2D0MTIrYAukINnwHHPdTMC2bt6vlPZTKR8aBGTXxXpXp
qcVVvEPXWt6WeRfuTdQpliRiTXemjm7eaJMHq8IbI366ZmC7Q0fW+nh0IfCiJb4MoG9ebeOH50KG
DPI8/QkxxXutEYQdv5uLt4jp9M4iHJ6rVafGs1WGzqoBNOC2Dra7xIIW0zMi0WVDFvCJw+7wk2kq
k/MFDRUNG9HNIFhfzjyi3nOowcRfttOcKhAo0ZliUsnsVL+Gpw1ZM2ktrQxOHwHeBJJDVXhH2O8D
IATwsnBKh7BUQprVHfsUtpr7z7LBwPQue44JxxZtHLDREiJpa+xfwf00YnKbZEiXLDLmtlT6mlbI
6aB20+9Lnh7BsaUfsfesEZiirXrLgZEu5/MyUfse2xfHWexA3IIXTRUGLpytO9kndaBcVRxRuOZJ
AkhWKLTvA/nmmPK9ZYtcVDox1uuiIB5sFQ14XGB2akGXXLvbwXNJ7b+9YTxN9ZIGYZU3VeXRfHN4
NVJOnSAJTBgQItpIcWAksjef6bkF0Bc6kKh1Enp0BOlgGb8WHc+pJDjlsVRux7hDD/GkDsAWgJJE
Dg0ZkNP3JzwcYMPYI/VHIcdJFJJW+hon2U6WRf+W6ipIhUbx+OOJc4YdrylMpvFh+4AzlPUl3bne
CcfV44gUu7/ByqGMGDbqmZ/+heVDcdX8Aa5Mf+1TQU7IIlhDdDWdPJbQ0LNkfiqEjKHocyv1x/N9
8cZ2ZBabp0/25GZkl+G3bhcUL+jFXAxBEhZvXUxZ45bIC8yRfK0lgyvoqK0ASYhcPZMXfZ9liBS5
x8i3szDscVHXBmk3vUiiVDTXdxM32ZsSMXrFmkRFMzswlaq6ufglgoB4K8zhI37CoL+D6xVg4KWN
WVwppgAvq70uan2g0l+QhBirCE/dzVuuXr/LC5UthoxmBGKLF370OIfhV38KWHSMuC77jNh7o6IZ
sXBatzxs5wT14MwEz49oKUXC0myqYJwu0s6wQlNDPYufPZ0fwW9zact2pd8y7s2mz/selpZBzdE0
YaAsKM8xN5k4aRuhADqJ1QQ3ChA3ZbjVv3dccsBmA6bH1sSUzKpAveb/iGgYDtpTiUOAx5Aba+zZ
bYwRnHpby4XmlyDww23mF8gJSEmqIxy5N5QXrbwc6EsH32J8E9EMxuX8d2hSZQ+Dorg69vJgKCsy
ZdkwneTBY77k9xn+ARuuPxp752CFJuG3eRJAg4V3P0U3izjvl5L4F3l+hCIyvzs7rTEaA9sG5e5t
KGi8LrKiT1Dvm7mJtAiO63m5xCG62ITw68ZM/7HGKD7+HbHIAgQX35RSG9bvrW2YzwJFtvmXE2IO
SN328eAeZ1HzBP8sBCeb0hU8FHN+3XDcNatMJJPQkDB2SqOof+O8tyMyFZAZVZXPoIzI89THrNCB
8duPL9DZROZ7N84jWo9IGTORDkp8XRXVk0sK/Z1udmXCuH/I4aUlAQiQzHtyekpHCvDR5dRSsGSU
jAVMoL3GWex+nOvl0rvkHFEQ0Efeiznb8uqidC478yfr5LWKYJULtg0DaNl7YQ+EFYno7EbTCf/P
DhYAxLK0zXFLwNUuNhEQnEe9DwcUSvDR7Gh+EDpJNqzlJT6fPeMEpQ4LsHGj1jtaFa5FezUNZOFI
ekSMLHiD86XKH8Pc1Qi0kFU3pFlLtvhFTCcDeR4bd5mKVoqOUPzis+iwHlsahTIHIqug6c7zEE/k
jA4MI+Drj7iRRBjsNEBqKGJahq6oaB1c2xKXrYgbmz5VUlucnmBKZUlTrBWnnBQ+tMChgCx1Rkg+
Ww5CzVey0hUXks5DvCB5utf5SqS5Dq5CO6jxQxE2iTEBIDrOqaSl/BB0hXFP3lDg+/ty77tAbgQf
L81XodPmJ+4jWR64g+gIBKOaEbsvBgQwRA2fzRWnpWifXQkuFb3F0G0FA8QEBkGIW4FJEnaxYxp+
fk0d47UdoU3lsVOzLawMwm3ppJUFJntfBDpEDRTF1E+vwLzg7K2FOLBYXcbaB9Os8CsivVOk17IG
I3tHzu9d4oZl3spikseDoioVCFEia4CTRr+7bq6a0Wgu4yq/EzDMyFd4Pjj5tNau5BdwCQ2ste2X
/CbIl1L21sfzW/qjsMKU+V73jUlfNy+oGrWQStapAoJ/B/j3mV0Bmo4UUtW3ByOrGG/YW7Pibsxg
AiEfIa+au3r4sSGFNqZAWSkahgkFbH7MvI5ayfRfoPqmATgmtq8AdtlKuBRMmz0jvJOJW8NL8T76
znYPtuZ6EpqNLd9V5ux+1/kKc5wClsdKHod55HO0Hy4cabO64EXRy6y/c1FM8ZKNPA5ONdEYJByw
qoayXU5fMBPZQCAEeFUz30MHLcSmDcekuUuUqi7sQFMZGzMHfYEa2MqX1lwchAjJyC5CRV5j2Vli
5FTmOotJ3GfmEonOJRsXtHASk6Qk/JGruljK7RC/uzdscPHgEhQFROnOMunyVDOxIro/BfdbSDq5
LCnzAb5udktmmcDQIbh+SV9/oeLfSYyrv5Bn8/DvRE6946XBE/kQ8La3DSI1Z42iMBCipbpKp7bX
cmAnFCok+AyGFZvGNHFgjo3ofMHSgliW1mQNtbhJV8isCiKmfsr/Gg3i7z/UV/KAjqoa3BWClztU
y2Sw82+XDWI/yXEDTM4TVFhIZnp08LydsI1T6lxZMXLJdPz6R7ZtUTKuP0r59z9g2nZHz29V5dNX
bspCPiY5mxC8SYc3HOw79JlT+m7Epv5CLFEAwuTF+U4G1G0HcrbZ005z+NbcWriS5SyqWrw/A0Nn
7Pftz45ESskpvioZtaZGbWAp/j2l0XTC9/6URlqroHSqj7SHcxFxoI2JnE/Rxz8kwivzHlBed/sN
FIMncMtOikJ0xcEJCuITCIeGhW0CuDWBhKJaYiaknuoJVot9QLzxQiH60gYhvQD9+AAlkDrw1Iw9
xfPjvb4wYzG1RAm5yWcbILweGscggdcRjjUM/sux8vfYWa/lhRX6Qoj72pKAdw/ZfBQWZAKSMKZo
omyCDgODcZuzkgKDgVTAmJnXxaAf0ndlAkGRVuac670usXNBeOkhZ4p4nS+18szYonhGPZMa3mIO
inQ2Ky1cdlZ3o73kIy3TORdC3tmVae0y1YY1hGp0FFup47sO9IQvxoE7U9vdkn5Ow1yIzKv/JLxf
R310Drg0QlTeUrrQ97q8xw4aPqbs40dqWDQKEwZFfMtGW4UMA2tlFANitahPN0pTuLBJ1oTzoLPU
R+obTmHgV/j9ET5hvn/zaTBwN7ARUo3yjc7EzC/JenjK94mjigLEf2lGtvSKvUCIzzm4B9ndLuQw
Y/86czPnFiTNpJFQPJESPlpSKgpgEoypR+Fy+eglbqWvPh1hz2bBD7k2dMcu/yjd3BzFmwZKaseZ
OLzxGPqlG1NfOHAIr5kY3FPZzPXuooE/nKnmvg2Berfxovjg/NO6bKctJhWBjmakc0sCbkWjD5Fd
pyTySBiyWVltMYfm3B+hB4qZB4NTrx9xHL5sTl41RfV5mOPH/C1lFeXOtMLOpgG1o33hx01TV2Zb
n/+FeGH3cqKrU5x9e2HQY0Lq9NeLlFiIIRKLySzwDcRz4oODTO9pUxL7acBy1RRv947mJBYPRkcJ
tVYukNDxHmmyZhxRzlr/iWZ5i0O0m7KxytiOgLSbyPM3b/TeJoFkF1Tx6y567zCz6QE+b7BrnCy/
8tHmAh5dOtmc9XoSnef++FezxWIn/ILptkztC96mVAJ7Leu+twd/AoVTvmjJY6ZQYbJE5LCK8Y84
GxcyNF2Giw9mXVGveqP/v1c7j/q2EjE3rsQ4prZ69jUY4YtdcAQtlaQcI6VqWzxV6n4Dm2ioo9Lj
AsD6/v1K8KlY0M8UAJe+ldxHHBhRxXFpQ/F3r1WxyNR7GvNqK6S2EV+0I+uelZQAR67uISs5NB45
dIBx+gl4UphYcf/5wma3pYsh+cFubOrT13Bw0sqZsPWZthhZjshq8Ay/eHMosxhG5S+qAwJsuf7K
+T16SyB1V0ZSjNIeV5l+JbS9bIgXgFWP/5KSdaI2YtCkFO4QoQLpIWpaNyHVK7klqU3UKf44VUy/
jSiQFfRJ6MaeOs8ypSEOPAa44Jv5tg1B6CJ7kWabXl7Zm5sOaAnncKfYZyhFAzy0dZDFp01jYhyF
blG95MxXrMErWg5rFIKN5t4R/I5TI8maQcwTMW5/Ibsl4+BdcAK6iktTNzagYstSFS0wDHrJelO1
Pv1ExE/mgOg/LkEwYVcZsuAVkGN1Zr6AIGnwrTtw7r8eArzpTGURdpJ1pbwEpy2xqoGxyO/cYM70
MekdfxaK4H/1x0nIU7+y4cuGfXhUOPiE1iiYc0OzfTGviR9bMF047zRVPFWVPTX90K5FZAZZAKaM
UbBlLMWfsTk83TFj353nwUbLftjHV0w1pkIKy2RGRAWCOIN0ep3wsLzGXxLMy41HtMpvMif6jh0B
X4TIpador5TNhy/ZjXWd1Fc79QiaPvJN72FNLxydQxvUm3OhDa2kvmLlOZhAA7BmDN50BTd6iSsY
jccfqCgYpp+UPomuCxCqGuguCef4zeO0cNONcBc9oZgEkZ9l1s9KxLgQKRoRB3ImANa6d9Dg6war
dQyhxQLYbG/yerUkT0C3HsXPo1pdVKyLNEWNBERYHvoArfgw/0lE3XO2c8j6MJ4jCjUp9XVtfGFq
49c+bAN9CexfPxriqoJj9cHqhw9sOjrGrcMb+cwcozV7VcXZu7cpmbntTat8ErElVreOwUenHqk1
k5gvSRbAhGm23iI7w8nsdSTk0pYxdcryiiI0hsGZ7i15OPsouAXGpJG/EziUFxvdF+MIoIYhIRFT
mEGIzZeFVSoNrxx83mvmcb7CiSIrQ3uUafTmvBVtDtVJNHboOOnhbLVmsw+ZehOY2a6fS4m5PdiA
OLsDzKN/QmPUJl1TWwjB9RVIsTqeKXgDpZ+b5sKMTmd0NpE6IefOM+dMGjSdn+ARoeN9HhguF2aT
muFvy8GRFniHrLKUPwYHfkGHHWryN9DEffXrU84Bit1xnsps8ZibzVz9uiPSGkrIPlMFDnIydZ/T
D4WMIkviNWHYBtoTNKTZfJdacWG0sg67WZPhjjD0hCsE86izWGKq1VOj3ZMYPs7rHGUTlYXBxNS1
BjPD19KJUd9ORS8NFcO2sg7nZTNhQZTGc+NZyDIIO3q89VGvc9OUdUgXRTSs8TVoau+Kx7Syvnfm
62QmeCtH4CSrEATfQAZyxwaq7CWWN36DywFiX/Xbl6YeKRaMdGs7ZZ2F6N2oJ5Qe6/Y31mBGs+bo
nntISUO9FJVGqfGIyN3XCCiNu474uzPFBangnWqu4g/Y5ZivXZK6T3/AHFThq4dmxOqLe+LhDMGX
2AHSIQ0UQzXtrabcgfJ8UxlTpeFkS5hB2McPqmEGzrnTAqFAnxjjcZ/QlrKyH0RNMGG2s2RecoWy
gbqkHvD3cBj9wghhMvrt3LkFtlY2KtRMBsA3kML/rSDZgB976YQKl7RV5H2DJQDSGxqz/3+4mWqp
DCi84UCfKyCehOa4Mf2lm8lR6v6QS/JWT40xrfnyynDlDd+AduM6gVnHPcNnM7ThySLc5gRgR+ip
cq0T89vUo/oP3Xs5/uvwUs9nXwugvsP9vhlWtBIMZ2fThc7ZtbVocRDT8K8/Z7Vfd7X2kVGPV1Or
BmmLFmAC4HyMiR3jLuA3ePRsPmGfO9+LdBzl6Yh+lSzldJhfDInNSfEVHtonXcZiu8228JFNnuKf
tnQVob2gowhMTOp9qjJKg8WepK7NChSRUbUtT9ioF6jICSMwbBC0lBAsgJffgMyMGm8gYnplpOs1
aVBtOcjt2JTKI6Q+Bs7Q7kkMkFoJDmFhgTLN3ULAKl4d+k0OL8VXB4XMm68zSMoRXSAi3ZPIPuY0
KYMwjhBG1A6o8WHcyV9QqgkIWRCCiiLBqjPoAXrISjtl7urp9GZZ6PJnpFMGoOqbzrGdvZAJQ9o8
HysNQ1Z0XldYubtfllxLjwGukRnyLTrWioqsvkQ3jIbeUTby5gHSLTl4JkYpnAmfEq5qXBKgGpG+
yf0tzUWu7eHEO/dlInn/g5ef2Bl5VZwwbyYjcwIjc97syWDtTDKQSSDYRyRcAIIzi906+YHFWQrG
hjH1/73+3x0/45Ka/WJtC+Y+p2jqKMJnqDzFjhu37mGDu5BYy62jUQ/3qsepVJmY8Fbqgc0WaeYZ
ZjQbAw4Wd8onYCtGlk+z1zYGV2T+AjwS7pMPkRohGwCPSpSgKmtqSxuqVOs1Ir8GStP4jP347QZO
BYliO7No1/+288YT4xkWn5HJ3hbvYJq5/yDpVIiwCTHhn26xBu8+FTH4RUe7ZoOAFQS9WY0pjjY0
DwtrC02ujRwKS7W7wJLBuufX+n9/PcoJpQWmVoLhjGQK4+sA2QR3WOgFCdu/TTg5AcfLa5kUwvUq
QFhZ+wK41vGjL6NqEG40MMvhjLvz/o4Dn8ujjtJnY5KQ2HnGSogDiQ8sw7S7M82pmvm5QRPUaZUN
CBlZ5bvsjyueqf0/Tw6kD5TwuI0ceLZoy5o50kRKnafDU7h9Ahl1K+MybzpAboutaIJehppD95Di
M3wGLrDJEPnepDPfl4SQg25onBxnTo6CQYpkNhy3u//X0zDkkOOW38td7ZACqckRmxcSGFX9JSMS
asr4XiwfWh4lpzAcy8h4mR/WHKOtKBn0D3CCjX0MIJqncr8m5Q5+iD0gq+ENmsnBuKBtjOovZhAB
OU98UiRgQg9eE1agah4umEjE4w54aEX3zdYxS6tAl7mDfN2ccLpSDHBygWhM+j9izgV0KGpjWRxm
m4U+6u9/QR8UOy+VOaqwvO5PRVN6X0rUOi7WudxHhPgcFafWF0CZWPq+1AosFHbXon7yBDDOYZY6
i/k+vnh6vKAHIzRExGSNX/6vS6xS3amT3ZCTRs7FDgkkty2Qz6pJBKVNbGdT+xbuaMFqzwNYDRi2
U0fF0nVvB/dy2m+F67SLBb4au1HiONPuf8/PPye8oxdmg8hcgInt6MAqfZzBgd/n2uO/RJcyHV7Q
4JsGNKsX9bQASnhPjQ1vVQiQKHdIVGEfvmxa/+Mz6ZFUBxkKv/oCcvjSd1MF7wmpJG7mAVycFURL
v6G8pW/FPEg0jobA8GjNwHcQv31abCD8S2WDwZnszIWbsJau7TTwJC4n+hOliWXKyHNyAkBAlg7q
8+HkLBWg3Zu56VzwMkm7cZU6VnFbiaonCYg9ZU4vCLPvFZG2zQ0TuFbVCnzVLHb46qLxhANaZfpY
N9BHH7OMTWXjtyf19LDEu6qdxn5ptERjdFrvFGNTAEMwTEZ4Q/I94f3ZcT4XcYHPjCWCVH01QBX7
IfTO1uxxZ1it6e0Ws/voUXu5TVV8KYCz8CEZRXZZRUwGk2xnk92AO2LacGakrp+awQ4nYd5hqDdy
xKKVogJN9IGQpnfKmhgv9LYKyZiwfpEEwptiyCaBETyCyPN02+jVn+KmrYUFltkGr/ZmPu24+UgH
A6A1l/zTEsBtpSsKUM6Lk3F0THptqKVIxAyFuTHtqxcYSDhLkVSxJ6S+/fQgk+37Lby8UUBN0lgl
71HEWrGJ41Ditz9B32AWG3ohlbEwB+MSf+zQeJKi1SCqHjLaHw3jMCg5uC4yA5+ttLbKEMpq3ZEX
xyk61xWeZZX6geRGe8zcp+5U4ZGvjz3bgHzaG78NMNxZecOaACbwLe5a5yRtzG9FWjhStjAfGf4S
bHtgypEzgY+im1yeQyDeP6y4RC0iH3bLv03C/UUlwt3vHk/3penWETsqGLK0PFNEogXvMaDg5/RV
O7JIAyVZcWV9cEPdI1ljbLa4ekwc2M3r8DvipQ7HfdDUuZpPwGaQ0WPtvc5fSlSRPAx/C9awh99H
f89bhXC/g36vbNGoBU3ITM27byOUdBvnsobtUaZIjs0JtSnYyhlUl3vHmdMOEhazS9w65cPNGXOP
7be6s3HyhaVae7bPeXlzd19rFEGTc/v1gUxKLXdMiguHDayp9tsLZ/69M1g0UIybKymWmjyEZMiS
9PKWllw3+CxOcw77qc+V8yz4JHZ4NWxaHqaE0+nvqhsGrfaHYKsy4qlAL+sApUPNuugM/Tw4SIiG
hh4nV0OGHG53hWO+/Zbkxk5L9GHv0mkDv8Sn4BfsmrPG0x10TcSarbdxYo8VsF9a9HYj4r+NIdcw
C/OT4MZR0i+Da6ih4snrJAmcHWuD1D79aI6QMQdkcp2OEb7mGhDwGarktkcZKv2eImAY1owTmwAS
N9KEYAVDZ07Jh/bM/MX3bjTXe0WD+NxFeAJ+1Rua3Cg4A0GPnBtuzbVWJlBe23lV0sfSUcTB60jf
cFPnqyiGutPuXAjas8ye3KCcAT4GI7M/za3HuSYrMN899STVy0vbfly83FGWFyC4gw1jIwFP02Y/
V18nQw99QlblWPBmZFOmSw4hQ4vsRdkbURvOMORxaI8GTFi/Cs5XBjCwrmNtxGc0Awu8C+9OtKAs
0UGgt9ZYjeal73Z3W3UMhqkv26Y9cCNhflLGYRdGZ9vdddnTvZYnsGBduzVnhAnf3MBddgG7HlhJ
D4Qewh42O/RmSk0Mh5uKTGfGd2FZssC1SBmWr9HiUMzRscAFkBMQYs6VOxZx16c5fJlcxL9zG5Ds
Z8iEB4c4xiak1+oajQ+Ngi4eGaCcrdBkGeX7RGOAKxCkT9BYpU7ZnG9y5EWnlNdv7xLfyS5dqdQj
tif1EWHsPAlpF9eohFOVzskPNiHxWMPaylQnwaK9vDN0nXMBFg4WSvakFQaHfAGl8AzD36jwiUuW
AKeDk/kmkhwOLbTe3nmp3oedkPwsZ83Ugh6Sq4cX/aDFKX8z6xdMkJZYTwJROAFaBkXoMZ3UYMok
HBqMneeMSuvUAByfQrCYeHawo3sDCPjpGootdIvHk5slx+b+Xjbb6O7qXMKq/qQA0TQWWrMLQW0l
8OsYV5Gyeesgew6Sgi+EWCx3/tycdKJ5tSo7zGqNx6+H/gCCNsO7rFtQu0nQJISdfBI0nwU8fXnL
NG5KN/2DyYM0gtEVUDZ+OQ2lbYC+vvyq3u5XdxwmTh4OucxAq2zzmH7Pslu861GcvpvyMvhXLhjE
pQaNQA/EyRxm8O1ULp3s2B5+2phMHoAtBC/nQUzXVynpVPh3NyLtBrs0A5XrLBELHyYivsJs4aBK
6A0odqEUS1CvLdmrOnfA6qi/NMCHVIibS3oEUqKd+AZt1nks1BP6RGUQmLmkt6vynRiH29zHNBDh
RJy4PkLni9Hw+TtJft+XHWqk4Aczx5aYNAC+4FubI8dGQMtI65NSmbheYTRmWs3abvcyK5c8gnRy
RgLmKXETX+821Ctth3GGCXws92vIPaMgyiJ1cpssqnYU4l+fE59rx9alHv4+FXVfFSh1Ns1ydc0P
XFW8GVCmkjvAjI+IRxHRkJ4Do+LdqiMBy4I1m5f3uCilHdfp6fyuFIA/5KZcwDmHR/umDPaTFif5
TnNcu+BnSYT1ILh9s2VFwTefEyX/0jlUMEw/QRrRve22PaBkaxx/xDUlHgj0yoIK3Q/RkyjWzKbX
eXkfYrAASsBvAqsWtvMKmYLLIsrt2Kzzcb46H/JOIcPv8tHjMRcDC8K6HYUqdi3fdPki0DIF8HWo
oTaeBGJNn/Qu2Ok9ywJhjZ9zDwMhSa7r80OGKHpINy4ZApFLZd18v1IGYL6ZBLyo2pd2sj9v29gx
hkDL37qx8E9qzoV43mFzCajecbUijBBi9ONs8IrNhekva+Di7hclhxyVYBeHy9hJ4QL7GCQgB3hw
FwiYsNNSncliSO5wznHx77IZOptpN0gfOsLyUIMW3hOUn3gWXQXWhQhw1193mqa1HicuSz+kI4u0
1YiB7HVMlOzAIIx/N7iP+3TQouJl1oRonMUiyNzQq/NipQqE4rFzUDQXbbzBx9Z5sLumRjKOcfma
XSD29N4DUI7Kb2FlSA+VKoOaM392ExEs+mwzRDTq3aC6DGe5R20oOpA9nPZVi8fCItrwepI2P5Ea
2tZBtldFQDXGcWdy8ZgzoajaR4cdp0bF2xfHascpJXoQ4jzMAMoQAwU1QcTW2TozFhiKemHFRZII
ddye5eTWAgHEYpE0B9hjBxdjxrz1VId/wstw4Tr7gjjbeLCSzAc+82hNRtVXRR59LfZMmVWE1ULM
2Q1PtbNsqeZAoixgRNHN+r498Sg6D+ye5MYDWESH90+pbtV/Z3CvLJSaRcEa40vOPlrY+GLFL/HY
mZjeWC1+VxyAcYxHASDRV26uA1sTOUVwx6GW2DBRq+DWNfPtpyDZ4dNeo6I4+Rz/1llEVPf79Txt
/Qn47J+p1BEhAhK27e+wmcYgH56CLcwxOpYJVerGZTrc8CU0LE7nHGH0dF9F46UJihOYCm8RY5J0
vCz1h4psgiBSqFNIUzlti90hD+ZjGnswyCg4/LUXQMG1/CLu9nINOGUxheH1fNgQqm3TlLk6HVnj
bvl1li1JlblyKY/lz9OxhI87LFaX51J/FUDaAhQhezZBjkssoAL72W2IPV8RU8yEVTqzRmdldRJX
MGfkwVjosBvy3ts4WWUfXqGJDXjpk1BZ9ANosQyNyLznXhacqoGiS2DDQE7v6VFQw7Nh8g0/v7Bw
g0ZC63Vrwn4jlCCnTKIUSQ5yykW5AntdG9u7ltQwF1olhJZLqB0CzXvZCsiqlkCHLMGtV3qJw2n9
9QKhU9xfwrRWa8cN4tzom8gkAbr7OE+TCLKyfsahVHamSHYcSsrvHVy3miECtZuMifWIfF6CTZ1P
RUwm+TFVD8c1ylP3638M7ihHd8TAazrLSMhUoMvQ3afZzFpMkgVAvLsG3kulv0cvbWYCYfx51+V2
k04YYbaYoI4KHu4tu8+5ZKbXnsc5rABt5EYARBI1n19574O5IF6GdC7Z/D1ltEATI6eRGRNHsj0c
kZnoYJ6ugqFCcG2YWYl9HoGUxhmN/e0GhgL8aASubdubnx8FlLvW//NYm9emCooWg6BMvfqcvPlu
uTeCQYDOcGEwLJkJinXXu3n3pV4cKX5YNd8v7chlDepNihkxplm2p4mO6uDaA0xyhIhYn/FaH/zP
oQXNv+iYYxmEBXfwGeWfEu8LwjH04pnrN/8jSZ467TgBgAjA/aFWQG45SGmM/EL9MSjGPSks8bUy
riPy+pzLN0xPxVsn5jwqoHd0mOV5RAKhhE1xZHShPvIM0D4g2hKQ4apzrHEZlVhU/7LUW6iB9AUJ
M3kytGxSY5bPub0mq2sZLgUb+VQZNyzTpsLGHqRJuY0jVjuSddeJ/Qj4/zXLdbaqLU+x33ZP77Xl
stBU5IR5bWtnW9xqESz1hQUP2lzkrVD1R726uMJGi08g+qzMyDGE1B4YR717iJpHZZGqjx5GRvF5
THwsaeLiUkrM+JPnPB6BTcSfjDleRAjyMxvMkGo3IfH7YOCFW9guSz/8DobQZMD5x7TR3d0hVQ7E
fnVObOFwtPil2tfpVFI2EKcNFQK6fTDJLOFaOkDzIDB/4DfDEyPNCxnj6TiJzGAT+R84N9oC/f7Y
699fGnLlcQ9XTjblcH1W+Er8uNiG0VYXO4WLE+f5MLeGHMDo9UU5948GZVM2D5+XLHLOXW9KbUAX
4+e2cajIGiwAo/5rCn9v0OL3IFFp77Ya+1EpBY4eKOLTfhDW1n7RNSMtM20DkCqen1KoOalwU+XL
tuxKCx9yQFdVCOOBioZsSFMVt3pgFtkPKRCcVEmEnzmS/vSN614vgeRWNsR1gT1PWWtNxigmXxVf
9BeuiBEU+pCfox/gZrCGMKGPlmDC7eBu+iDe87rGKclULYtP+3Luv7XSwBjLn4YBrQYV5dKxUlsz
0S+koyssf8Odo1VoU2aMXV3S7WrhBiwUkmP00bIbFT2NpDSVJXHioL8ZoPrHKeN3MJyXDE++Ndcv
zLN/DsnEqOFwvJa6AErsGpgYalYIHURleAZBFZ+S7a/wRC7qQ92AWNgTI2eQCcYE0KPYEIDxWFu4
1Ei86iIi71jZeqwGsoSauLBWznfAHyxldZNdWeI9vm1kHy1FmZnjOV0p51AR0cxFQH3qPMGQxGCh
8+Fqn50WRyyMOqqLD7s13oVyp9KIuJpsCbJ+QqcWrYjj7F1v6ZrJBr+3JWPRNq4kNL4Rs8rkUryx
rb+90af8C7u3RwQg9N0unOV3HBK9Uqa6ZPtdRogfTY2kuibbzqAEDsV0QWoAnt+TVfLPLI+1jnS1
sKcQUGLACskUX1Eax0K1wFD347NNIZXhR2yss9xzOjCB/72RGTmIoqQK5+MhpxVQc+tUc+ZS6vKP
l1LChZaWEEh+2AbtCKiB6vY/FQlQref2O9JtVvOuev/+TGEZRKNr7pFTIbR4jgXhiWEuL4IQ6Omk
Rh93YkgR22cA7kWClPRJKSz4kDEjv79O6UiXF+ElS29cmI8V7rGs/2itr+oqG2uvhSP+dG3NGKK3
lPhN+K+a7517Fhhp7/PtLA2hmpnc4orCCd+CH7czEcnqqY9CDUiT43/UJSVWrNUhtrKfov0HY1XO
BN4aMs/n5TaHKjXcF+RKBShAdmi0A5Rw/+CH0ukF+uK/75ZUJSzJZVB2dORJNGFyOLahgVJqHA4n
GsYaguw2mfrfu87vJzNTeHIhXh9rY5e/DM9jM/LeAGNKB0X7LrD3kZ8B7aNu55GJsjnCIKz9p4fL
XabJnHCcYGl9NLFyQQXv8YI21WWAW+HPQP/Rprf1thUSlXdlMTDKuTc5MYPhXbLb4brshhup3nM5
pGGCTqDKl/JammLLoa6o6nqnsfL+aGT32Rrue3Zb8dB3OFFSIgwVaIzelPbEhJmhRMYq29r4u0t+
qS6O9S2zmJczWACbdgbh+y5p7u4e74PlrCcDy96BrLZ6SY/IVmV3YLAbwqAp9TskM81KiAEIxGIs
SCveKgl/oAeUdy5Qo/TAr376AsU0/6S68JwowY3ROwsQKt/0uZIytgOusBv1sp8GxthLp+v4T6TW
sUxcmCRHZ0xlLvreZ8Rvhp642pWslQ/4/IYSoT0+qmu2+pVTZ7kBkkQR7v+JJkI3QDITCjNLU/UH
vBaMkGXVz5LsaivrCuGJXxbtSf5cVbw6Bta/+ms9BVkX/Dpk4rp63p8NCmGVsCWOsKvUruG3PSc+
R+NZxYMFvPcF6uX13WBk3O+/susIhpwEN7yhB5R8Ce/0yXFhJoNvvxj72gQpeZc4y4nKAchtuCc1
mtiU64YeQSTh69QjzsEsIh0dFfjCmuviZ2/OgAfRpcFZ3MPwwkC3Hn/18xT5NgPscDL9KGnkzt3s
ywFXAIrEGX9oVT/2gs/UZf1LtRTxKkCZN5Cipsy/zs71PgLQb/9yEwqTkvRT6IIZw9NSm1qQE2af
MFClEBBNCVdDIKvf7o32YuYg6sGoCmKz6DaY9JDrcIMBo0oT7tNS1FpjA5c20C1N5BC3fh3HWQQO
OXXIhlZLU1HPBeUNDYWmxXiR58yle4wTZkD60MCApl0Vxtuk+bh2Q0gpIctkoq//FhhRyTvMEqgC
+GRHCkh7h1rLcakU+iShUdTMfpasvXgLI1Dz28Uzx6vOlapUaA+kHeBFxCpMB9+QhkMXTq3Dfgs9
KWjTh3/gZZtRWQpHOwXXAIjbSYMhGmxLcQYJHpS2TcnYVlz7UU/4Iav87rMJPWA18rJJTO/Co41Z
c/UimVBRk40c0eMpF3BLVD3vKgkOevNj4iobjBcW7Op9fIK4SlmXms7GIodQbo/yAzgzfFbPcWOE
WWGFaxAM1NAn1/ZODW0fibK2/gCqu+PvE1ROWCTX+Eco07RbgXcbwFP8ia5ls6wcZ3FkcYYTyi4N
AdUgAiG3vjCwwc5jQEsmHEmzSAmRoVt49eSoTq/jWJEHAa5uSrJN6P6LPWSWHwyU0dnw4U8QTU4B
Fdk5BEVzQxRgD7zKNEwmhi1ku41kq7B9PYdnP4CaOWi0tH9L7gT+U9uSMo+iK8MCAtK8zyaCWmGd
op291ZCMr8dDt+4QLPscCx3T8sil2gc4RSYnjDYEnzh0rlbdJ9d3r52agxMKzQTAW1hbcoPCKcfu
7rpTQejBzsQw58JUDWW7PLeeSI5Zc0zOnWNYaHl7vKjqh9gWWqO6dE+TVn3ICA+h0tt3yA7jkKtb
tki6biMlX9cgXF2oCkaHn1fcwdRytIW2JWDtlioMKD1sVAmYxlhNBHHA81QGRYg54bUvR9574tY0
U1uTCNxhZBMgnd3vmSdS/JSp9rj9Glw67WyRwwc2y+iOGbivVOMezm6EEf4lvYD16c0N6oWo3hh2
fU6JuWI66o0a8mJHOf50PD7aP80fpVH9E0D+gFiyUksp4izbcFBbSD4d0YP8fUteiD1OCbx47+Kh
zX9UNdpaM0j2c4g7n14L0tQLo2rvbfZBn47xnJV6EEI9hnPer+H04EDII8iT+UQI4XClX3+5s66r
2Uuw3pnoWPuLc09eO1Xg+FZUBFBFRBI1qNaf7zwsRMqWU6MdvjvyPet4yUJWH+gcIJeuir0ZC5Y3
1HFJI3LoBRBea0FXz9bJqiaK5azW4bQ6J2WzeXOY9k9a1/sjccfUgsDVJCz7rtwt1DCRg9JJQqby
aqNUA3aXpwGIpAHfy1EJzBdlGubz30MppkZptBAkfV98vxJJJ8KN4YixEycLuuTg7Hq60umilSN1
JEzLd4ZeKXF6maW6KM64HEHjJtpEOTZ9zrZD/nCUj8t4zZFIjBv8xwEnypQ65hTwkIIVrT7y2COc
Yz4FaKAAo6O1opNF8TUUm5DSqJCn2lE6Jri2RB9rbc1ru1r1oD7I6ne22Pz1U5B6f/x1W/c0GF6t
wvjlc705yi+KGkVKOVL0J8lhrxUxqfjyPWmRayck9U1zkjANy6KDuiprouobnByiaMht/03UldWF
rTuYeFPTQxEhZG0DwToh3aTaKW1wWuQnGcariOcyHin9MvdeVWIq3hyev/D/HpqFhf+Loz3YwffR
8SjLnLi/Wg8hx2bHGUhAbA6PxB2iYu5EDIrblfg1/4QnEuxtg0ZheUFBzcIjzkehtfFeBJLKn0OY
in2HCvMI8QJOpMYiqE9t6DdM9gXj1bANxA0LBKOULaGRihVcknxjRipQMkisFWrfHE69dPPJL0WL
wiB4aMfzfkPEkwYQUz8AExBqmHfOeyt4FoVeRDIyEMS2tP7fHd8WzqcgfsCDwJ6zv2BbFLwQqgEz
/Fc65oKx0cdxbiclDdPPM+SZhtkcP3bbBXHgyuZTW3RZhekWLX/19SIKIihUVZxCR75+OEAPIeYv
dvwxM3HIFvDLdocWO8C9vCPpx6o7atpf51XIReWe8h1tuAoax0L4Dck9VSglDow+Hthqs6XCJK2I
+Qtt/lP2Am0JmXDbwxb9qj5i4pqu7pXe10zbD6YZs+uPyoZSQvv+t2lUVIoTf8gSlyQgYh61PJrO
7JFvsKfan2WN9xXBFbuqEmlvCWCb2ArHgYCfPGGbCFANMPmMmDCQu5tMLryDN7F8nwxHLIVx45ho
rbf5nTSb4ztlEZrjIgTYEZul1Y2FyIOyxwNYLgtvduOC/Cc7+59D0mlQx5PAfnab0Fz6uFIv7KX7
PHdmo5RvGCTk069sbKxgneMVnXSKudi61JU0Dz3q+41U+0Eyj5kgReNT5bJsnerlDEqEbI/y4ASS
LgmfRmQPXMbkQ3zke68qF6cf7wwoFKgLBtRdfnLtfgrxbQssf5ciA8NKsEghPzT3vj+AWhGZbXaj
oKIbnPA7fvPwnVBmZatdksxh6bcFx1VB7P6zN+jVbRlTmBPYZVt9s4928pn3lMkv7qCmbNGgc9RZ
XH7srDV+RfXBBuqkzFPU8aSOxiUnU8YkOWhMNKNs38zX6yZKJxPRGxK1WB4kcalspPreP+/QqQsY
dbjecTtL4Y3Q3lKaX1sn93ysAqNigQWMLWvNR/w8qAegKpUqITVhbAZQ0qK8s2tmI4zNUgqRPZM/
vn2MxQixCRicuKBgo/v7a6WrE4o6WpoDH37u9SYvIgRGqmHY2adzUGMmuY9R4PqHjdfsi7zbQg4k
iRrCAOqGuYEQt5LH2sZNMYrKBlQl85gqjfVmd0tOL4r9anS4FPRPWtHCqKaKOjrL8GRtKtVLvrA/
Eyi8VP3UelJeTAc39yxr93YOPnp67Kn1nk+XRODsvfjxAIEySXxvRB5s3Lo+TltGl9h4z0n9Nxpi
2tRWMJQb72OrAgcGT8Lmgeky8bad+edpcpnVyEiy+POgmT5eS49KTwkrAVQ7aYxZ3Eoso5v2Ip1x
14qsU5kVHhKOd2IxQp8X1kbXSw/255F0w087Gf7gVz+ChKESIxOXP8m3mYlqXeHkBkTz4vGhX1aB
Szm3kjpu/CoYJ5pyy3AQt0gpxg7Zs74C4PiqebXZAM8ciP2vMAjOPS1TrgS0uDGKNit5TYjzP3ZH
IHu6uvfAby/G0XVgVNCHzO66tC0bqJxN5onxbBQWQbvfYkE0G6LH/14rsmIHe0TpYYDoLOxJXXpm
Ii9JQXvm8O8/ssaAxR6F5tkgabhpK/qndURoyUvssIeYlnV3bta4ZZWESWQEGkDqNx/RZEP9gKWE
3QV5TnUzayjjrGFkVu5PYviV1CH07jfdVphA60e5e5FuvgJaf5DuQVo3dyKI7hPTO6oPtBwjDyf4
5CHHyE2j45iKzWEAimAMbgBkewd6/LzPFr/dYhpOz4TeH6gtUEg+wUJLUCcmr9x0oQOKRW1Um9To
FcgyO9GJzPHw6h4Sb4XyY53bCTGLDVVgjNUu+74VXIHFRjq6K3ZCFjg72GGqoSCaAmoX/AEbQUo8
7n/t/yZu8pME2HkMC1oGECYj/L07uucoZFS00S+zCBXm0fvmFLHQhF11+QZs4tlChRxSpfF4Vfht
ImAzBQZfd1y/DK2sECDPjG6zLJYJVyoQLDDYaEtbif8BvTAWKv3Gaq6tb4zlXSSy5yVDhxptdSmh
itPcXhUz4Z9Rekzq0XbztK6mOuECM4kynxRd1ygjsrGI1k084qlY0ZDZ1HtA5qNA54p4QQfsqo6i
0wN7hABT+Lx2uID8rrKQwWkKVDHP6uTCd9Gz2rdDpBldWICJXSABzeTA0E4usBOCkGFQjoExN8Sp
qV5itFc0Bh10ED3sRxVdmhy+msLmAE2EIPWMsvEZtcKvAffErUaE2vJEjGuj5SgeWfQTvnbFEYVV
zMQpHwMt9w5f9piZwt9/Jqigh2PsqDifNDw6186E9Oy2Y1YQrCOsj6Ny+ij7iQ523HAT/VPWOo8B
DLwx/o19r3x7YhNJA3jbgzam2b71XSkACmUuNpEucp6PeT9YU3zeVOFF2qfwYRauiHP3NsMdK6lv
yxj16C/+FJQBdv/k7KZ7smZBQnBGHFhnywBNafeUFchkQR0OKzQAKvm67aPD1Dju67f+hgbiH6yO
olst6OqnWBUZRSxJhd9DDjkF0KMNgm7oWG8GQF74MB5qIYmyR+PoyP5B16x3fZ0FunvlFayS+ynE
pN8ipyvGkP6uIyGQi1D75+N0BwyCd2drNYL07keqXsccV4WU3FQc4nktjON7rPlxM4GV4QT/5jvz
T84P1+gpxBPCsqa5I/MOcZgUqSSGM4wlDDVEfbfCpyCr6Ed+6faaJ7uYSZbKlBaNGl5Sob6mc2Uc
SQN9u70icXKiY1u4+MpQB1/7qFCZpTjOGGgIgVmWymbyxL4RjopJK3Z7NpSN+GxSGxjyPivN8Oyd
ht+/eB86D0xjVxXvVaqpEQAVd2YvEKyUcyEqSVXbd/baiDtRaLcS3ccgjxU+xDnsPj/KwCDXfm3e
y8b6yE1S0xMyLFKE2200GSduzzzLALvy+7v65kQbrx9xRuvgw3C12uAfZtZFlou79igSoKaOXSHT
ZSB+4iooz4IfxtAee5p7bkGDaSYt1KcjuSnMdfML9yWajKbaLla1cjsJykzTURN/LEqo5dVmKs6l
cGpS00V9n6jO9vYusCeKgaSvkVz8M1+y1aaqwoWrXUCpf9wPQOXaEzID9dKF6QoKeH1TRRhw1wKQ
WcP+0sPj8h+veG3prO63BgX7NOoqPxX1yqvvp+R+l0wbhNR6103sAH6mil6yGd4Tt3utgtZLOQ+t
qlRY9hpUj7DViUegBEc3IVYKU4+dRHBK/d/g6GnOaxln/958xhTmNq/cROwqClI7roSVT8Wsj6m9
ADQ+rpRX4+BzWLFXQ6CNbSro6njFcJiQ4HT3puwNZK/CzNoR2DPKbJCoi0c6ZbWwTs/FwysGCcY9
BuGv4x4aHDI6TJXHDXoUbVypEgXR9rMni1wUu2NB221Uz6bm0FXSFEZpbr1Ja+wLcwaAFfuRPm9H
v7GnSzZZ34X2Y7TLPBxWHTvEyIRkxm17QwxAGbQ3bEl5mRcEZ94OAUnESAIdRhmIsF9ZZJ9YTx01
+R2QRTCkqPi1C1LBPS3CfQQBZO9Pd3J4dVUFxgoLynFWoHxVUWDbMYnGYG6oluK3i4ayfZQ9+jy+
WtAdgPZL3xdrUvmzCq6HSj6r1vQKH9G4loQv+Ces53GrnmI9zVQ8YJ7g42uf1fD4qxeNekipXvRp
Gsvyv9NGDJyGDNFQGc9FVaGPBFviyZOTdStjtdTQ+moXUZJaNugQ72jStoMXwxWNLHWYugpEGP32
OW/+Hr+orA+UO8NQz0bq6bQfXVx+xAN8mKwdagex3MZKUGeC7HATxykFGHc6BSVn1uA9O17eSYtv
juL2WoFgkMCpoSJx70FvSvHnb54skvT4ekAAeNqK0lwqjwAwv/vLJoiv71FwTVN87V+1tYiG6E95
cIGGEm3y2EANdFc/WA/2JYH2G3rJSga5Fs7lUMcN6JU7TzetEed8VhqyliufkPOh9sc8NfjtDHQy
vu2L342NpBW9dDIkK7d9fKZKNCnEkVR1ib3tgQewIiewPwu0sdTLPsk1cxjpaktSrcG1t934oquh
eohpwKB5dg1/A8rgSjEl2tKIqvMLfg3WKz9lFQr5A3wHdRGwk5Ka2l6eRlXmzFLi4l1ebMnNLyf9
ofiNwsRuhfMMrcV/tYccYZsUtvp1K5yOuyb4m7oMbES+kOiRtuk58iZ2XnOAISbaK6AsAY/ns0DJ
2O9husHZ5hFH/TRu136Iktx7hyRMVq8xF5wW35arLpqJuViy7CaJWuXk6sbFFBFap4S1L9LY6tcY
6wEAeknXaNHmk5YCSHWgxpcFDKYw5Ekn4GoUUBVJq5axvsz/eQWnwEEkBqNGPDVjADIx2BtFuUed
5WnIgNItUXRK3fpL9wEobv6BTiM0moMoj7N76DrdOr4JeSY9/4eYWpl2JRya17iGCE1sEWvGLASS
ko774N+9om/BiRh0kUE3UJMsHPhAo7n+RmDYAR+IxlZbl6MTFGL+jZBmZfM+nONHsrMH53BYs4fH
UE5wboho/MKatjggRir7wbasa6+ech4NCE35tmlVfhCkN1O9FgiplsJxIyVtZPELVCZsZLst3kJM
Llq66QuJpS9XkkXzYcuCcD+NB6DgJ8+t26hqa8gRlDiiekxLErxQVPkkCNz5e7SE6GkOfoJejEk4
hglaozFzIsc++VUDjgjo2Cf0TnoQR1jOttnJH7Fje/DNLuHMjVXyBwKzHi9bGc2//DDWhGYyZFIj
pN4D2AQlUJKwAn3ltoJZEYFffdsO9LSw4lLzazTf8MMW1TtZbV3DMWSfK/bFLPbs9FEOImFQxo0P
TIE1WG9Ohs3+w3ofprDy5Ubfd4chw3+IrlJeoly8Jtw7Cys8mvtCOEri70ikdAduPjo3/OXRnO/C
qGzgpQq8Av9CfhmYtsowHPoXasD+Ay6ibFn6PetZgWNgcVv7Tg8vhxT4g7Ra6DZnE/PgfHsQbPtk
Wf11TZVyQHcSpp9eZcWVe+6c1OuEMTYZHbUAn02BGMEvSYJcObQLS0as1ZynQv7yO23ChUaqM/l0
p7DJXTTvTcYfDrt4mkCsaV0Qdlh9xjdcQyYmuO/iX6WMn+Lf2ifp9G7tsqQZy5MusjxsvBiaEcrE
ztI+c7mOO2QurlcQ943i2vJMH5PnMpSkcxtk2OEYyDPjAngPqByQwcullqMERujW3bYdykuebowG
bQljj4SlvZ30oOs+x9gXBx+P9Cj3YCc43QEfdIkAH+vRbKdpYNX8osIuQaP0LJkqszB6aBIe7Bi8
gbWiFfAEcQa3rp/BbsD3KA9TDgT35/wuldZ1YLR6ewL4fln1hxH3MXa2irqB4a9I/PsswDyGmVxP
B3HzgDTAGGZ1yeCJgQrxPiz/okQywvgCMNRJompmgecqneEnscC3gNqeoZUsZ5JlF+FvOfJkGMCa
gsTGrcIEOgHfctFSP+6sUSTzifQWTlLQQh5wXD7vn7TN0RW6xxAVkdZcTqMAO2TZuTkDE0ILZeab
y9Vsf23vlPy+SGem/rhhZhRKmdO/yRaAw1/DhSTdkBIk+NoJMagIrfE0phojzAbL2Yps/yCma2Ir
AnjxDZsQIrSYtqEt0a36l2lH8KFmZAGL0EyAOH0myIqcdAA1cQyR3fRzuxwFRyf4SNlMoPQELcM7
2rxXUXOYgxlAWvuOLNiiOgv2ZgR2padKQfht6tHzYlZk/U/mBDmCGGLlBiOS7Wo4/+32lrAfkQ1P
5bJAHWtt/K586Nv1DtacW0S6LEjIRExCtP4Cyz1vFFJKY1yRS9jnhJL71p7jF+Ktb0W7EvXTr9fu
gXWDAPVnuUVZ4H0Jw1pquNst7N7F7L4SL+iQaEVkv3RhB1QP6pJ65fwCExZq1puFONZbwZ0UYniI
YXaa5SiV55laWMiGG89MsBtixt+xnyHA76Sdy3zgVG5uaPQo+im6SlZ7/5/7UUbrR7HDrVe4ly6U
i3/xeASTZNNSQCtES2grdM1ZqjBLbdAIYWOuqXwOcOuDopgLw34n3HQTRAvJfH0a0cDPlSOHYAmu
MnxCUkvjekwoBjaXGaJ+6fBdKF3K5aqqE1TG9/alyY7scMEC2PBv/IHUUXZtL+whIjRO9Gd8q7YH
/TGs1xDcfVKnzXVJhAZxC98s1+Uh8o5u4lxYwz0X/lpN1ZMjeEFh++D6fLuflnpXPZ3XmRGBzICH
68sT/lCEZOZQcBi5Fs4VIsOihCW2FCgersBmlQV2aYfB8I0mn9DjUBTYb39CrIg5Ovx0yIC08WTn
DhZJLNvAmLBPnQIJeOliVusVMxibCvPzMDkgt5YfXh64Pifl9UoPhsy++pnqtru4N7F0ekBD57OQ
g6Hln8VaRu1Wvjc2qvEwAJSMCPb5RHyn+t3wvarRt8RdW9Z429FoOSAoUCh2PjUONjJVt/pMZAZl
pz7vXwaFZrTLuUgrJxyCVTwv50IMl1bfO02PlvVAfNoggqo4NofnHAJ70u39yBjLgit7geVIFDE/
MLtRzDc7b9A19+6OaIhJbv+K7RHHP30LowzU4gAPEJlNi3UU40SMmv47Wwx9EjSFdNafULly+EQ/
2C4O1qcpBYHdR3I763i/DNu2yAHnRxYfFMTdpCTlP1MZvem7fvNHMhSV8VnqqPuw0jIm2ZB1LZTm
oLyq9hvgRoafP+zMfKv6KFcacfWtqpPOFCRCpU2LNIMhdOQFIWM2qTamuomkGK/KJoZKGuFDjzo0
9xaUnnQP62GnEU64E/6O57U/XFXdwB5DTOPESXDzwqm9f1IlYaRCUZyDAuOtvlJjFwuAU7SYyLyp
fZidCsbrGhteKYbxgvaiIpnT1+tXGJyPAPY2QF2bCLy9ZsKZ8FTr9/yslp/WHadQx8MuyGSlOMUj
ou8ZfOdPYJKVc9+9kX2AbtHni7IJSl4JrTjYJAxpI8uysHvf4tV/AEV28BBKOIA3P5b0sHpx1omY
XSBvIG9Vu9fKYyDWghTklT8xvjJgzAaanRxvvypYTzb93LmnAChsdjBz10drBF0/G6yxgMaP4XhA
QHlzvwB0GCth9epsbk/dQMGkaQU4hjTdVzNr9wpgd0XWbr/A7obxElkDCm1nfODmcLCV4KCUcBu+
CNnv1e+qvRAI4IGmBuYlSl7VtHDANT5734E+cgPGaeXlz0znv2wM3ppkb15Ap/CLlU9I/ZG9xryL
+u0V81EKJ/UU2IFjlxAb8X+KBPTG8IyN34cq+RmqumE0NqPyhrOAlTpTEeFaGba3WWlD69PB/Bfk
1HnVG74tkFXPnfqmAaw3CJgivFw72RZzRle/xSEkvO0MaJSwxGPz17kxO24ed8Z0qBzgBWaubuli
6atc9PftUFOSrKbCzHcgXoBnrqySQQXBjzGuBUv7mzms8/OwHpRboy9lrAyoM6U85bNMGWV0v5mz
Hj2EM7F4Yk9IFfdg9ccYE5d1jv2roQ2A/85InYbISRs/Kx6SGZDrFYbWka4fQuEvmNMgXGj3lKfD
X6NDBFLwPJc86uuq+2MPw6mtWvrn2V8ccQm0DGf5PVrbiX8CVrS+t165EXpUKJOZEFnQC1T/dFk9
fMUevgCn2F+f9l230MBCMyAqhywDa62NjzPC7+zDsZD0bSF/GiqURXKEAHh9caY9Jz2mdLBUC5DF
5B6+reFYIevQGeR4muOfRWRnSmyoRpCseFGA28x8v/TwKrcxUMc7h5bqeSzFDgoeNiJz1pNyXnQw
jrvvtUR+WRUC4Q3KZ8kJai3GLf53rWQD1az+bSs1PMKHk/K9W1DE3+2P3PpoTahou0A5PKb0is+v
2EzJIl6CMgmzEh/el+UcTL2Mj4/hXcVgXuKfiKdbNL4WNnpOi+5LTGwzjkLqELbwkTDA0pCMC8O9
3MPZ8Gqce8H0Jod9kds3m1+Etvy5eMJGXkIA1hnHT0xOk2959/87Lakwh4IRfRxl+FcxjNUbd8qQ
AlalLMX25odm8zr+iMZMsMMjaCbWC6fkxvIY0lc6LMtlAb+MMNS1g/0xyMjU/nxd7rSDE3GFMMSg
tYij9dFTcO/JggNKwhx6+se+3z1aaPCVItbVtaHfJEhWxFCYhc7iVhHTnqI1tcaqCDC/5ZODD7po
56buK27rFxEgtAdKDsYVir9OxIBMPKZgz6rSie7ojVlvuAqwVhdtRiSpuErnVATodDxrA8nz/+iv
5N21EAGYRLbHJ8FBa5TOJ+V1Aa8Op/c1two87ILbrPZSJtdcoXSYm8f9v+QkYu8o/u327jhsyVGE
BYvycbUoLCIhOZDvyILP95gTostBe7KxdhISoHeWSRGPV8cxMLjVp8XDaUTbF6nIF/1LUvss3Hb+
DsxIcnzBYeGARw6YHy4qfr5kT6B/tqp8hv9zyXOupzYiHmIUXnZ2rjII2RFlD1j/Z0pk6jad/Fgp
71wngOQ+sIIJsDDpvztiertFb7bsHInZVT1wUJN3otgWF+twU8JTM/kbE3AllH0AQ7yNTOm3xCmR
oe6pSZvqbh2ehFvZiCSWz9JHByT1cz4WWEupHBXj3+KxPZVp19avQJMdkjroUro9z0CCnXOP307z
NLRE3IV7Ul/OaH2gmhPvn4vSHjYPjAPEbgiXlSNx+Ir0TvAXJ5EeYS1wYQ7R/LwGAm/Hig3xOkn9
zGK6cy3A7YCd3KacnD4HT3T9gv1Y1ovZNTPOhlwbZfwjMMwm4zxMRlsLiKWDh9YBD9GE67T5ZvyM
ZM5VrZFULY0B+lOaIqk14cCZIt2gCwU4/l0cWVym2SFDJDRKsBZ+a2IkQXpuj7sJ3S8DCBZ81jdP
jRvxIh7TlubkPAmDYHr9Wypy4oiSlampKQ5mgJBkGY74wN2NnoT7m2uUqlpCg3vz5Nd0OMq4OK7Q
JCG/p6Rlnn1uUHOmCj6rCX8sq9d1qMVwvz4OpNmZNFnZvZuf729qodOYlDfA0EI1wutBUE8dmpGk
PAScNDx4ec3j8llOdKdN5f+5eTwFD/IRExaugu70VQIErLaU2oRm9OcSJ9JOBw9JU/BEYj0qNP1M
zXrd+eBb1Hv9UZardkjCy7ZRUiqafnYQcJRlpY722M5ObK8NKB03oNENIVG21QTGBMOBZbzi9VtL
Fa/w4x8FOzNqwoeuTWGhKCT412oL02ZPQ7Lv3Mf3Ihw8hdYGHEowyF2tkssHpg+tNLejpgbpmijc
Cli6JpEOeu9YJL+WfRzhRGAodkpKumSfQPruX1s+HxvvjQJ/M120cqiKabzmv0qj7Jtvvs+f0qdu
rD2/Xhyil4dgLBlBNimhj81w+NaGuR6wazM89jAb13OctiRakl1+cDWe2Fo3RYIeapoBdbpnW0Io
Rlni6oJhJHw9WLBny5b7GtaXG5hZ/vwLDB1MUsQYPyRX1GzILxXXICAS6v9ML1F1zyQHOPllvCr4
AEGOLY5i4hsy+byq8nSCEC3hu8tunALClY7tmgk0Td8WXa/FaXCzR3oV725TkxVa7vR9Wr+kVGpB
nNmwKniJ0kq9s8FvhJh2gu0XqSEyClVoTRHyqRD2DwDCrZMuGfVSkY1aYQRAngmrw8E5L6ZB6NHi
RsG6WembgOdXnxtpmjtPYVDrEZE8djRieC5Xv8ScBHeV7+vyfn/vEh+yiE212hQpd87/DRiWBEyt
xgGD+hISUHD4klI1E2e/hzep2Dx/ADqEY5sz9ywpLI1h4q7daWT7KncK+jCGjifujkIZOjYQXE9T
cIkWTvDww2qMZpGXdST3wHW0L/0OaL4MnW4dj+FcmkcTgSx/Ur9hmjI6ZownfEx0pSWZQdZJevhY
p+mXeFD57Hyb+gVUa3tPebbU6v2SPUeo8Mwcau+36tNtPMPTXlN4bGzIn+4oNLznzS5Odr4qnF9t
Zhi4C108eIGt9AfsIALTA1J3scwAyw9fvVSbsnC0jE+UHW7fAtc9kjlVhK53FOI/uzFwET0tJU7X
fvbGSxP8Yne0cBnpCWam57LRZx+eaC2ztFjIj+ufUJh5heVz5C4p2d8ZOYZ4rckQ91WuoEFS6iTL
MVLmffll4M4jPHoPUH0kqv74fVS9BSwbfHP4AJq55EWSM090Zd95P9KQS8V8zdt3Y0hcfgGQDOvT
/cgG7ODoqSiabqsd19YZyU1YxJ3Y7omQQWG/1ZM5Z1f+NDyw9Kx2W57dzLFH7fu/eJRX1G+f8C5c
tK9ze/SgzhzQn9fv757IxZeOqIpox/HrqBUDPOX/EqItcDBzbxGPUET0W/i6LxWfJZSSqFZKmL9p
snAPnD+BhqLq0CNx37Qgw0bZTGTnGZRLxV1LvlEowMZyhhDK4yWXtOyiSNtjzP9nFIatdPPYrLIT
BqAxSASI7ISJV3gaFjDLCA81To2zu3+gaFNSK9y0LW84ot23EaR3gPE1k9av5itbGKQYPAicWFvE
3CZdz4qrt+UqupTCoW9PVneS1QQKiSZK3UyeaGvwLEuh1Q1IAO5lQbN9F6ztty0Jc3y1jZqX4F7h
wEQKI/xg78RSwSY6tryA2XC85bssLy4/4OHNyhlWOGUnoJXBydJ0piBijCgxuK0xBjGL+3ki0PWx
BVEI6eJmziMwZPIUY9t8tgD+zEdB1X2wZE6qEK22vk25zjAI+DakDggY60ehGuTpBBUc65pOERUD
4g7baGSz4vm6MTUTT2ArHSDtFAFwkpNtJU5T4bRQWuMBcniU3lw09fufYRSmPzGY7jyf3kb5PfGr
77dyigBEEUNpMBWj+PXqKUjoh0DChyO04yh6ZabWOgrmWtEzHBcUV8tHN2Qz/wR8twV93nKWiLAD
aZLv3dmYoYdA2awaAcOxsA/nCaN4rxdASHrHcITxFgBD/0hF/xNdsL+18+r/udnEMSF/hphESkrx
fBsvPBe4sS2yxU7yShvlTvNgCRQtPadtWsj1L2Ets7Uo7plOWm14iqwJcC5HI/jn54oKHnXcIrUV
oG+Qd6IjWDAzbvVBbA8mNyOEK4Ls0X2eByfznun7i1kOHqAeXjqAGyaVURfmqA+9Vbhpkl6BxTne
aPtFIZAWFQ0r5LuZSSmnViuGV0Y9Z8+CXyWzaCteL3nJmD74Qtf3R9uQaQfspTClt8zKbybINMLv
VqvOJTt4Ir52tfLpbDmWuIJVv6+JpGVUE8GEgcuJnZPEealrVRaTsXAmfpTjIkNixjSX5Zu4o7Ys
bjM6Mu5uKhqWZk/rUqe/k9KcC8jCwI7hL0x8VXRmzX5iGoPljlV+MuTGq6lvsyThJo2bVqFOUAJF
4mo+jXaY4tNAAmJwITboz4ppUUJkysqDRAEtIeg3JJ2VBpMjqBMqWyBL9Laoj+4N5JzRLIcyK4kE
xwz+JV4YnQhUM4wPnXzrl14tgnLwCbz6RKRn9E1t3MXpEKe0mnjvmZcWNsdR7FegiwjOxCv0ciJp
1R8Omgu7UTOZYhihJMRrNO027hFmFZ5f1cKQtmL/y86dR0tKK9i44heZiF2oejrMkFWzO1abIag0
K691J3wjHKdulGsly9xxROB/X9GhGSXqW7CPcUFOCexoOGt6YbuXsIlvrl3lm2xsMtDbivPi99sd
gFXpmufjanyDKQw6YeGrncmUqhhV7kqFc1oDb/CrZ2VD16en5e1jhSD12qwxfiIUP/cvBHkRRNER
jGjTqfDVnEqNQVDVnzUCMbq+DstsWuDRwsalye7XxcX4PtWzKjsGKOfR6SkS/l2UP53CgpfzGdJG
gpf0EaWJNRP8qsIhGzZ5t12aJzohRI9mo22QHVqXCm1bXMJXQv8RVseKzQ5vCLM7YVkzkiXMmHbP
+gydXJlEVd3jcEqfslynDTVphC/yKAZWJLOdi2Hp9kIGVvesL84ByFebAksAPPVlYHvl+VHaL9XE
mnyaXTsiCKcSpqgEKG79rqrj0cqr+JYuaghab6/b0DWcTBamAntklJDpLcT6zBe4uIpm/5KbT1Fn
q0FYZIwI8yz7ctkBktqZRGefXSGvARF+aDoTmk7LaLuE1ZeXBbPjPuyQlkkLLpPmYQHzTSajJPCG
1u9zxUcwR+MEtLXUDqYSMNN3Zvh4rN5lWtmG6RTn8WL3hnQrtysw7BfXaCtWz0psfHN5DsRL3Afd
NImBJVD5uusiuKTKY65oXb8UBgiqjjiFOf+BBQ38rTnOVJxym8bXwEQKD9vHtYbEXJIDw78FAHBW
pnZbOoBhZJNb2D4t2QE6vjBj36xdHwKbUD4olC8DULnRc5cGjiUPuizmAYt1TDbZBzRvunHgTsC4
cftLce1rWBV61ORzvmsr2/ilKX60f1V002oxRa1CWiOxXfKkgvP7hqmbCB0LEkV8a7q7Qfb9gzOg
/cMkwlIRgD5N9voRvT1rQ1yH1axrZfiDIYZ9g/XfK26Dc9lDcqnmMr/m4aAMf6SL0vrxfswC4/9l
v47tZzX4Uf5JL5I6vkLKEGXTzAxBDja1EjQ/bt3rcH/g3mDvoidT4jMGA0nUw9ObGU1lPvz4ndKC
X9JqJoMqfhhV74OKKY0geQo49hWY/G5+ittVEca+cXv/draEdufaLUOgCrgqnrg+nJNLWaxn412X
10U1pH8fg4jvqdyVXNKYOg7JV7/U9CvcMP0Det0GFArBUFY8OHL+IHiby6jzX/678wajKpIp4ckQ
0uq9Fe3DbVLiTxY8wxuzcsb369E6GgvDaoJdwR8FuwDYrB826XKDcj/w/uo/m2kLkRdoolIiEjBR
q7H2hV04TKvwf0bluLqQK6VntIekc/G0GMoUriaoqNVQ5U5V5iNtvIdxgFL/+ilSmVhUUQ6pJetY
4kgAWYSckUGWoxjJlDVoe78JIDuY1jassmlOkHbwIS31msXrx/VOJiw1MANTdndTS2uqpAhUw837
DXJSnpcPTn0qNKsxt9ueW3QMaa7rITjUa7i/CpuNxk1gKLNj4TG3EBV96ra3ekl2Ju1xURam05Fn
DkZ9aKeHNBPrD+akbCOP1urck8x9GuI4oBYlGQLU3uS5sXwdxWwk1UCDOhzKoxk0u8dy3THpCML2
iBN2ZaLS/+qwCn7Sv1A0blVuIRBSkpJ3WtMlG7LWW730wnb57REm0Gq/VGOEn94rZjRL95Jcx8Cb
W1WSTFDSzolKXwRowdLCwHJKmWe92OyhW7kQXFnjOp8TWd9YfF2ofXsxpKJaYCjGTdMZ7R814RDa
G12oarKt+OqDJKDnciD5Ap/BG3KbRTVlWKOYmSK9CHLbLmFE9cVNoBFmR2PtL7gm5U+0jcxm04qV
oXeU5VUWFH7BBs22vjaGsjgHuPlIIR62EzN0K/NUZ7pCu/bEcoXqIHPVkn4RsECzFLfM4qbKTL53
tCihNgrZohSSqDp4nGGazfNNbU4Wt8izO0amseDP3rBX6k3UF1Ff6hL7o2M1K8ImZZ5E+VEsZsMj
eiB7WrGE3Yvi6yoJ7ou5SDNNwkyIoUX0ZfL82TpqF7v524Phz0dJIIXmy6tV4yipZyunpGvD0mp/
N4Agn2v7ePJIfoDYHC+kUTJggumLv1PCWqQBc9Aj0QHujlyyTpRwTufI0kz56hWIol2GpoBzIfE+
P6riFlBIb1FfWLV5L3J0dJlksey6tbgdvfkMZNaxczRFCGnXqJddOra0OwZkyYRDP6nlDnNyCrAk
Da1XVojQcVnWNcgl0tAw9x/dGl9Q//lyYUzQBpS+xYfI2GZ54vrn5hdEyIk+iid/6DPgkv/HT8MT
6t23Bbl3DSNbBDuljrsHHhO+qxQUMIGGlEZDo74hbb+szbzJF8LpeYUQL9D3FTpB7blNTHf0sAHk
Zmz6laB8QnoEM17oaVz3jj42l25p7VSCCPZWPz0VI9wWbVsjrm+QZg8Qtl0zjsj61oBXqeuPb6Zu
UiVW7hoCh/UK5ELUwocbmRbWpJUQM7IasGOtvlN8PTvN5mu4KsXRYHNUZw4nFL3zNF28rJhBd8AA
a5OvSegpsk5/D/dtmC2jXeph9Bh19DPrnCPm+sJ/z8rX9MH0uTXJdix9dSgY+CnGHE65g+/3ExTc
MRiOLvcqdywi/9G7hDkXKOOh75pk3QoBcUjL+dso1A1OkVZWxOON6YGODSgM5Dsl3EDHzUywsTla
mWy6oMmiPVNkkUxpvRLnQmoYHc2QE1nTMhdgnxyf9CHidkgifinCLphiw5DnyeAo9vfpySKu1R5M
0DE4f8QkcUMGgQPcWbW9R7W/7khM2Q8qvX3kaZxqH+ks402Amhxp+aRFhTarShWO5wYoas9LOchy
p3q/9tU4ueFfzCORWQTpVVzbiXIA0cOXEPlrSiY8oVtkBhL2gB/XuqKHqSkuoQd5tudFriJPJswp
QVOJFekIFhKSbEDpRCTGSRX1OgDC3UPy0zBLU3R3+E9aeWrd72hQgs5RIpTIAH9+D5/t/+NEscuC
0lh07DvUm4+eFqYmHlXoX4wEs6p1lbBagw2vtqus3r3sbaUdPHUiw0jotIvMWMM/AI3WQDbWRPry
EthDPdHa9B0UDuYda303yji9ClOaskFoaJPl9s36/gAuQ+gFLFxn8+nurGRUdck8EFnZrgv7VkCe
Tq7VbTQX972ErfGgVLGk/ssUU633eq80RMwv5YpwGyxJOj6DTggOqpEiGTQ+Mw7AjFQdNiYmyUaZ
cH5Ni1c9AOBx5a+KH4/B+18epTiiPr5FiGouiFBcwWJ6N9+b7BO+B+XLGeotqVrLQU6PV7j21j3A
lSkVQBgtTyNBdkvy4TLW7+QhmZih5xRmSfUudo1GuyYl2tG88g5pg7Ey2pKZPQNLjf+C14hwegYf
4RwZX1ZHIb9hqYFrWTuzfXfxgZboPiuWkHOf3GKJMXG23GB1I1sVZrX8juLb7cWuZt1uLIrQ7KYa
y+F4vizNafSUTW/zJE3P9otKYU/uyDT1a0nXPqH/6tU/wBQB4GtXH+6Z+9b5ZJCYTOX9xJGu8x0w
bTRdVVFwvCqxPyRrSGlWddtW6xkm2VK+DZ8VSXX64CUKGWcSONyI2QaxXtmzWDxDB0Q32QiMFPNf
kwc+cKWeYQ3MEda3Kc2lNgcp13giaMr/3zWiDfSi+Tl6tD6ZYi1162e+GvxZ4JDHGV/9joTFpkZ1
OUzyeMUK0NTxJtGXaq7REEc3bLLZDn/B5LhMSQk+lcwvAe/LakWyRIju2DieHFNn2OyYlCZnSls/
ICYyxyKJdX1blvOmBaLI7XjGphNTLbBv+EiF+htckZAHto67iZfc27EWtq6P9PuG7NIW4Trwx01K
NFYcHPiXSfcgAVTah0wROrxd0Oy2oX3ZsJKnjk8nUKBwjnCLgxlgoRYl3DXJvjZ6TFbiXXBj5fOU
Vt/MkPXnxwYEroA0QuZauGR2fCu2QKkuV3lJNR484FDR5UtkkF5eZmBGreV5GAydtiWiopM4hSiM
gl4/PfNbbNy7DO4xSuebLa7PVWZKFX/4OLDADdGhpON5YfeTPJuAVb70xZrMaHZnotNVda/TKq3A
LIFwYp5Iqfo38t8vVxrtpUdbGOYfV18qfqxO+Y0xsbxzjv8FPReGNHeP4V5Vz/c3lx1OozasxZ/a
NjB/iuSGWn2acL3ryVs8Q4218iK+ZydoNrREzKVl9R8fArUigs73uAr2iNlyZFjoy8xFPWan0YhJ
EVqXK2wvmlEhQSo8mdcYFxyEyr4/34a0d5tmXLqQoFbZtxp/Vwsy63H+M36TUWz5qv9QJE70KSkE
HyD8HbcJN+GN9iN1HmBYjTNKUGzRraNUQmGyNoKyqxgy7QEikWI2VrDaXDOM83iYFqGN6NtDbuW8
uvRi8j1LOIOco5oMiJeq5pNoX3p5lid819cZrQZpPuD6dG/lfSOP+VgMq1mjYI5Hx3SmlkXTMBEY
ZQkDnLh1B+OJxj3rmVEmwJT41zsrLnwby3jYGBPozMEV7HJHK4jwanpDJqFU9rcBjguaukzguYxJ
buZr0df0esdQej67b9SIGenK1bGDiQaKgTecs21bcC4ETbE+ylIr340EiY7p7NzV7E6TqJEGBpoG
KHtBjq00ihSYKc0Gpn9H8qolvbaANz9PKrPbWV/afCjb5JYuqKiWZwetCPWZsBoANZK2OgYDqT7Z
DfrwDKihFqmXl9Em1H29tFtZJmoAK57Ar+Sd594nMx9A1kgvF6k3UonsV3RD/GHRKF7nafIe25jc
FtdQMGjyNz0Cnn06yBDw/e70O60jnKP75upFmr4ceQVrlAbPX6gnJFEX9uXqxZAjTXoNkc2oPyzH
+irAPOLUdDz1We5D6I/E88hcPFDhc2HtFxElvnv3x5cx92/O1F9D5Uj2wBUNiC0deMdvQXOXv4qf
SyoeIhf7/1OXfH7FhXl5OSotNCxqpMlComa/02FVhiOaZlTERHi5GHU5RM3+s3BC7Si2JZUQd7Qn
HC7FnhXohsiQDgga8ImJoS5tDGY1wAS2xL/V4YcUypGyCDs+hKfcK+P6AW+q1I4V8WYS7IgxBtOM
Shn0xxjDX9BvFXTb7LRoDAH98dUWoztgzul3rmN5sCMEtVm8jTVDV5fc5jMDM8s6275K2KjjO3iL
/aC1co+HuXxwRY4x7MT850HR9LNKeHzGCP6drxu7rDOfYb/Sh9fAAuACAYCvFNIzYEC8+xeH3rqI
C2L8fpSg/mwkX6NNGRwJKthlLxZFHAUsmo6l4xKyFkEnfuXoMB7hkalnvY2OFyisuJm5kDf4QQFZ
DM8211DjQxhmZdT1BKy1XF8wcQT68/j/PBrQLvZHRWEbsYX1UgSx4XNpzrPxtcrW6MZoeajXbiE9
r41xHLcArOVbdkT2N1PepinUnh9SnmDuv9/tyGdLhQW/V5smAdb6QOK5ecHS9FX0rXbfY2oS+qa5
vHF+OQjm65o5fMD2PjjTqVFOTgc9aYWtsxXOzlZenlhtH0PDQeaDddXogzMllPHkFFf0FWQ75838
bm/JinjkrEiHBF32oKcyZ+EAaVS5iQSdC2ELObKXuf+2bG0YL4v7nhnKHAfZBxynBLH5ae51ATNO
s4gdw3s1LXc1wKke9wCI+JAS72BR0sLFH6oWpmWKvAlzkteFfqsDsNdFDcS2z+ya3tAwv/YQTO0D
WadXAqCHU2u/BT6YOgEGC6kPbdLxqm3/WPDRdWt/AxycMmvD3R4LR9Sldhq8iGnNzewfBPdTuhZL
euwUb/Xdb3xJWswIIIwV57rqkGSg0Q5OO0YQ2gh406XcXZD3VpZbhqbr+SZ0wOjiNp7owLR+5YHZ
+0aph0bbSkCo3GCGXWgmks6o31FMZ6uiAvYxCMxHZYlVwzbPCFjy6trimX9Fafwzo1soPdwHmCat
qC7IDGLHBBwJQbyd1zGAoWmAhPCU/2k5Vq+1ccYvX4uaxt+fAGGVidq8TlMu+26Rt8CCAnBSog6V
7lmRX5JGtZeq5VwicOl2ez6OrYp21csTicKW5zdIx7v3Sj8jrRb0l9KnJB2AM2ZdFKw6l54KmJF9
BU7cFKWa5RKFWQYZlFQi8993xx6xuJS4D3H2HHxt9LgOJwEXIbDcuf6ApUsfz0wMONALMDDxpe9F
DjrNQdQsDjZxbiBoboaqRlx3bnAEF5X33vLzeopFPKfLs9VXIXbfQfMfkQa5ewZMqo9obWmushFs
vGY8M+YQ6PIrCS8cC1ccxCBId4WHVFwPhJENWjRF9/HHyNr8ZHOxSRf+3qkUasWa++AfVfjUgbs7
8h4PrfGa27w4adkGtpZwIDwYy1zC71X4XYbc64klDG4sSxavlKANRHixgNflDmfVgGSg/lyL5xoo
fAxsUZfmU5yTPUeEwj2NneI/SQs3Ib6fivV4BogsafcsExPZtyPFCpf0L/MIyVa3geEVuSowrytn
7vhHwj4yhEAods3sQeHKjIvlYVMmNqhqrAvN0jclYjAX+LHC1HyoPaJUTDY0SWM+OPg7lbEttnWd
TQii31G/L7N4jcTYj7lWb2zBPMzZl9K1Tt/i2ajPZNjrG0/YlAUTweIxjwRSN9H9MUeNVV5odNzL
dP+svB3CmzxGAU2lU2CfBC10f7/26SJEqUw9qFeAGrObOOVaq0PDjW3fHibJWpNEA4xgOv+j7kz4
R88KQJ6BlKE3eYRID32xVKZ1NvL10YMxzNU39xOpfoS5hEbM0c0eli0O+cHngs3F+n3z2RqHg68x
Hq+NiQo6SfOJ3WMJzY40L9tRd1wDJI/9W+Sqb/9MbtxXd0chzoIH3n3lpgHKgpVnjvYF7lNz9agT
ukHLrsuylRKLHFumV3EF6CscJnfOmDA7YVtm7tQJPIb792QS3CE4pXqlzlWiPlbL2SQfMUhgQlZT
P6d7REUc/oM73bDEmF3B7cILO73ZTzmXsZ3WroivYL+XMIkRpIScF6oFDWxWvH3i3o5SVJE0fUd2
zFiWvy5MUra0Ivrg37pMq/SfL5l/EFBQPToP3bJpCaFaWHlt20H8roq4lOGy9661s9vQ8gQQ93LD
neBQ1twD6Kq3ztUKNFTl7v0kVbOQcNhxIJZjH6GOU5df4srJsJfdz2STfSOu+gzExkU0Hi7TAUBJ
H8+Gaeg2LXJjTgYPi0CxTjA4fhfWtB63H8h67duDUpOKQSH1YOSJeRIteY3vVZdVuaQVjo5ux9/p
O5/lRAdwAArIWzVwTrNbGP94eevdA5DkA3ouOrhGh9+Utte8AvJK6GBAl37rfO6KIP/LgyBN0Coc
hLUJ5x9/2Rxk98KWQusBkgjIxAtwa5Wuhh76Gr4ye/I2RXARTr192D8eK7S/seexTOuZKC5y1egy
7wt4yJUBQ7EzZpZpYWvpjOhieTyzry5QLBXS4Ep+cKudRtwuG2WxMSJCPXG3/huyv2VJ9ZZkwxHu
cJMTs3sU6vu62Q45jGPRhp1BH/byuKiGn3iCqzA41PY1Qm7zKH46eVhEsFEwfQ9lsjZIzM70k2aG
r6vSVuhUMdFB72GUBL6PFdotnb1BaHmprqzcEvseHYWqUXmG2a8rBEqwu+xG2rokOi0DMKAuraFe
z8TKV1Ijy3w0yenbdahwg1JjHWfhWUvlALGmTB4efBszRB0CXHhoiYcik91fqCCTcN8VU17e9Fme
MEaTVjyBo5F6eOmtGarRLV2UqUZ2k4bBAur7LuozTS2/3qg/aIZNb4wN3qscFqkYpvMlHEKx+QkO
GoVehFPLU6v89ZCFjEelx8QEfyWTwjEhzNvD8icQXzBheANap+uxbyccWf13WRgIbmEDz/kTaLdF
CKM30NcOa2ayvtyyaREQrrzVcWxMxlbhcO8YApOumsid2MK1LKo48k+Z0/xElZS0opoBuSygeMsD
3ZO4LmF9CTnvHPeiJRyEMIpTheo4ZkKNF0jr/LlPJHcIW+HJwOx/fOQPEvlFNrHiZrs7tn+LjBcU
oNBcX1UURMSoKODFx4dMYJ35EpRlYV/EcGpbTpSeJA0QAJyRjretYRH3LJcerXQXz1dhhUfZkt4L
Ge1sHWi1Ejn4CPthKUhRdMayBn3QPaTo8NJ6xOravWXP5iBav0BA/fISrIdQ3x264e9N5TPNuRr0
HxNiYhD1a8H/HoPA0znBrZwtT98Zm1aTIK9zAY1b43X7xaKSY70KcT88RCe1m0vWtkfp/vje6F/U
vgS7knHGMpjpPQGIJqE/V2XCdIm0dZYyEhZisrTr/5KZ7OqTo3eLUumC/NU5+pcu7RHba5d5D5gw
xBPEKKhFo1vE0gKNif6CaIPMT0WG6d6dpDjWK/hEA/El3uBlkTpgSzgQSZ0OYL6jTB2B2u838KqZ
OZTbXYcpVa1t6G1k37e7knLCA4WM/olFwJ4NtmvKglYXIj8letwHp8PGg4JFocdm0L7E1mvbQerW
yZAPPkUpZTP0BWSf9o5wq/U2UQqEHkGXN33GW0L3x0UhiMEoE1osFJs4O2B07Zlk0hI1m7wkMMSu
6k1akPVrCaa8zF3pxBFY+uywTNu/7uXmrWZKRMGf5a4kvsZY4T23L3BUVlHsSzJnuYJ+I10W+LKb
41kPrq07JLfCwZdSe4BgdwL5vHZUVgOaW6oyPAziJFmjBwSeI6GmmsZXfgfsn0GEL0llwMRcjQwv
URCNE4HKwJyH8HG1CCjf7cdyvH+Y3Yc1XkMINAnNxBEjnnOSyC0piDpDTW1u0CsuL8dvVwO0uKPR
JjS+yRZ13t+pHhF06ZJL2QHQfwr6uSkwJ7A5Brz1kalQDwpO7cACZ8ZzMWw4AeNaGca1q9tNQPft
8X2poJmnUUphSsG+ytOEX5JFgd7tafvd9/bnB669CyqSnSmtu7hy3HmGKW6Zpid48E741zwnMZlu
3+uoHdNYOMtDJX7la58noL8OwVYr9veNFhBW1CDoEhkxgT8PmaXTvmvo5ZC/09Zy2+PRgBGtUhuq
5tXLzy/Pm3d3lN6SiV7epFDzBqd9/BNQkT4hd6vLstBBcULrW/aKCmuxrJkYNa+9xOQ5kPQxIduP
jU/uGZJ24tuakyC3H+0pB4Fns3AGKd8+cuHXfzqnmDuUnbu+5x3Hy5qXdN4B1kvl/FyWOpm1scgI
OujoLIYRNscZ0mG5F/2IjNtJ4AwxRjQbdTrKUNdAwLGKlBa+gYiK9CoBz1jjBUQyfvMa8vQvEH6Q
PYPwpQFGsR1GjPMZri7J4Mj026EHWX1NOkqJUcB65Mw/tIyA3E7Pa4JOq5J5oBgCYXM7QKkwJDsd
Edv6k2R8sH1xfuD2YB0WdcABAOgD3g+6njNsqwlASGvtOgiTWZF4wcYrCrRJW9ChRMEMlzEwx23l
id5K59ctC/Ke6OZhKsxUBXSbrX4mTBQOniiUC7e5tNQErNnCWHDuU63BR8rgAhiCXsi/pcfLeGuC
PKpjTbl6Y8vXKo3a199ido3pGBbDkuMNvIWtT4+Mpow+0BwpgFSStdspToDf+6/FXoBTxsF0Dr4R
ROsn8TcTrpWmJbMDaQ/IV7ASoW6T75Tr4+dtXCox0of5Z2acNCq+eQnpgKE8oOusebuvMIPGyF/X
Vk9w8UeA/AF0uAql6UtOGg8JUPXyJnHseredIBLOoSJv61wbmgcS6ZjYj/pBDZg2ppFkLugweDyE
EUQbfef9xyojDut+klrr+4j/hiDIZHYcM7NFQQ9evKEE0wex1N6JqSMP5uCbtZuyFH5LCGOJ3s/7
lly80R5FBDcDPLssTNBW1pfdBhO1vo4dvArVuP7dazWxUjjFIWwU3EUqwvr0Npqpl0ehjNKTFldN
Gr38jEKLdWoXgYOBKsiBN7eBpxT8+jzOuilAdZQOJn+ZZbXvqbvfcgNrFjDx9zYDu2cqAlAZs/no
2qaE0noacLOU2+jNe2lGSCeijcfTd40D8qDd2aVOrLlUQwwgevw31Dx/ygG32Q9TEl6zI69ZFon4
L6DuSJ5NStoyLkcuoTi7fEe+gEpgirEUCHtLxADsjYU8HI79npvv0OW30PMUFRh4Vo+ApytutEdi
Jzv1rqXaEdzxCzDOu10UDbuPruRUy+5H0m77JEWSGcoaBztTjAbAnHa8VCXzKNTgFlyxVWeNEub7
4iZjKl+cGRtIKPh7LqSUk+lx8t8ZMpQXRSFIPV9tSEPNTz1yUzUKVRE7dD2SXZV9d32JgxKzEysQ
fYX7bfnopEetHXzIYTeumcVuZQnbHYF4Hy5m/Rjkf71g0ROhn4z4NySZsnXqys08dI++uHkRu3C4
2o+EcwKyZxzyrq0mzktt39CAi56KYzspdOsiqLRhC507flG0kcqCkMJ1Dwrge/BcB6SjeZSYrE7t
m3ToqSIZFxxO4yQLbEZ/IjkCPpfivWTOCbLTMjyAuuBd2jBL88rsogGDsTlPobsBYhwAwNlkOhkS
4SwmQMEa21PPirHl1CDONzHWbSpFmqe5dNyNaHIItqloWVJBTplL2Q2fS9zdLjP67kshkYN5Q687
FJ1Jc7sUrdLIFBsvCEbOccEVsw08XbIRDtdDCwn8S7Ra5/Tdik9bZycrcxSb1FMmNid7bIAMsyOA
eqTlGw12lCBT2tlz9X8yocSfsZsvGt1feCNvIcumBugHwhF4KJVulbmBV7drENe9pSkWmkkPk6w+
4ISfoLJW5nlA8c7CIf1facwuJML1b8//t8oiEaLDzr7D7E60MRoBf492nGug7UUNnB/DmF83rh6m
l/DFoQQ/v3PX5n8+YD1gZzVra8rw6AlejabRRXlniE+OSx7GbHdYu05x/N5p5lyseEqtAbvvaFLe
V7V8JZ1/j/5mVkk6zYwqPX3jmri2W1xpYFPv2QxUu8D9MDW88uPUvISir4RocyXcClEqHaw6N1Pa
PTmpouN8h6OUW0bNwD5x9rSNzalLO8rm3tVaGn4huIUwgIKxzR4x/enz+InfxkmvqVNsRTVBBwWH
igHuYHX1XE9KOtfPersuTTOTTFm6ttTvy15s1ChXCEMFEBQBmQyFqnQvJGe+9HtGijWoasOHS17n
fhWMy/2JuGV7e6hTg3apUWhg0M9PDoY5V71STfVgljTEWv/ne953W7WvKR1YoyzltWySpNya9bFc
IZv2Duf7Bhit4ZqV4M2jXzKRlNILkG3xHapd9V4ucPNzh2+fhljPMACRGZfzoO9/2Cvl0KVf3Vm4
puVCc/50xL0BVpSEVkz+L1UgeD3amUUOmCoEmM7Lls5Cf2DsXoMEnfeBCre3zaaSGxXuAQDXXUeD
afX3mksOtmUHQagoeSQAdRE6jghYcZ4MV+ObRGDdfYU7o0hqnwTtzd0dp3v+ULz0EdvgJI5L28u3
LYK84mf2M7SzArrWIor4W3lOMyHbnU6kSRNQ6fX4JXB6xhyrCV37A6RXPkjRVXxFh4yqO3FzcjsJ
qhPq0h8Ju/0pPKganSQVs+JF3nDHMoXy3JLbx42TaLXlMCc5CFc6eEOuKUa8yz4lZCEEZO0n9kDv
iSS0HTAcqCuNDmf3exJT3WwKMa5T2h6B/Qq+c/z5gSdTymWG/LgLfFFP9c+ahEqmWKeXq13+WWwJ
9bWpzYdzuAIlPtvnqWc69jIo2cGQjmPBPUmD21mF2om3gHWjCRnu5J13JeyGe0plLvameVc9EQO4
iRr/P9aWrAQ5wR967AE07ndVirpruHywfgu10iuvLlbibC7anMVGexxQa4a59tytgcjpboV2mY4j
EUIXtsfg3FlKa+IuPFajqhlmPKxqPJJ8j+QF29UyMdeFSN9Hq/WPr3cjhWKzQWxCprpHOhDeLTdr
GufdDFaKJg0M/p8G6c+nCmww7ItBvJEXvBthukn+wugGWAEglUupH1A7F75gTSWR0/r8RM/nUmGj
3NuZgxl8sf6KSLqevb1a+Gssr7/5R/gGVbTHUjXliewSjqg+VmIOFAlwP0joSGscSAYMRbb6ecxi
GiADxJPcqQH4R0yHnXeGKWOdybZjuEwoYSiAEGd/W/hLH+CdSTwkpHwqNPkBsNbZxq/4Ug7ikA0Y
+dvl/6tj7DHoJDuy0EkTTGpWMsnNzbRbNJIAAPpux9cV5gN5S5xHAGJu0BGQu8lcNl39sgDyReYW
6Q/RsHUJwjpM0kNIhoD702/PtX2Ry2iCL1AJpe7AvlGL7MUjMRspyoGkpFxHo6Wf/XTXqdqArqrJ
llD9nGtmAQICf3urhQ2GlryyhfVo+1YJgD/MMnRxq/kBpIoaPkex8zUlWwNAf1nfN8Eq8IBhGdsv
DKaXExaULCOeQSfr2QUZS8uBs4c6/n2JI+Ux2XicTDI2k4PQjVu5K8rG6EywgeLqywyUCWUGokKm
ByBPPTIWd7t445EoOkL+4kxDdMUiFjbj8H7AXY+virfnmZgoUk3jf1hX29IWIrmDbsE0Lwz+ikOs
B3d/p2vyIUhWkW8L3eQ+wnzRtB6UZaYesQbdJnzawCE48Iq5LSLpCje1Ge3qlq7Itojy5Iw1o9Vd
yyHJlMuO8OKzSOfkRJ4xxRotHfFJaobu4+o6oBIEtB5UwuKjbagginPBkw2/oEtZ7jxFE1lm+Mhr
cKA2mK2FinBntv3JBW79BZ1tB88KygP+4xIeEmIi2M9go1EA5cxcPF6K7r8dV8ktTuf/I0EFeata
GQLlE2Y5JUeRoyUImOlXcuk/lYk5jaSiqSZD8tiHkqMtS51XTwHvb6TaKNei6yfuaQ6lG6QU0nnh
VnARDKwGqIqVqFnh3xg3I6U+wEzaMZkyT8plh/bWjL8tHMK8sWZR6KPuOZl4h2JYJ84nxx9Km84M
TaepEXvS8gH7CJkPdfIIbUoYm5HCoPY+aW9fCz0db7Jjr3SOdSoepvtSYtzpGbLEPd26bBd9XogQ
B50+Wz+jOnGkv83vRnBsOgc7jMwGwY8UUimyCSVU+7jarZKON5Is8VPqx3G5a2ByF5gBAOEl3tHU
fYnAZojCgNrkexWeI+S3YsheDp4ImbaB148m7qSJmUOb+U1Z3dSINttdLw5Sx8r/n9vFVZOEpa5c
yVO7scFLiF48yCtihTVt9/PR3zUAOeO9ZQ4seDy6vfOdgQ28RphqW+JweGRaIM/Ynj1pRc+Sghqk
xx6MvkzwZRaIz9JyyhDQAZGtrPmT3egJ0VgM0bjtoOxurDKTwC8Nb3dPtxlU3B0x+nCL+xC9ds+c
p6a8rrXgz6uLk2tdZ+XLUpO0cWoOZb6bvAH4gzT3uhWMYXNQmOsYxHd1gbeQ1czvprBiFXcTaKnB
UrGG0ZYcbYaTjyUdN40qVIAiM4Vin0GTRPLh8LAPS4bov7bVRBlEGVcZMyZWfkzwcEhSEyqQ82L1
mJ+Teckdhx4Q9m4c6upXG3CNJjp3u4baelXQJLDEScrdT4tcMMpINWoVZF073xRM/BxLW2duJ0cO
7Ofoey166BE4QzT8yWLdy6C7gE4WFkgyv7SKDmRGfl7bW+ip/RKxD/srYFv0HOLKnT4CgIDhxl6k
wpBOzx3fcg9EDL8W1jE53D0umECbwqrDE2ic3cIolBTUcD2sySquIYAo2lrU+mJFBe2j5oIxDAf9
q0bwnFp6tkYNDdsh8zKGylMfkLWV4LOWSStG/RbgOySFK/78az3rtL9g0F/58MJLjO/CWPTy5a/5
ljrOl9tHYi+i7c6Y4R7JENFn/bl38CHLqsGampU3DoQtsTkafst+L5IpL/b4G6MLRal7Ci5Jf6yQ
UAvAvv4qLP4fJx0GFCgfvqigRnrcqFgSzXLSOPll7hBJ4CU3WrYThi1lEGy/jGyeDAarSLhZWxUJ
Z4r3MwObDkks4yoQC1rxzHmwXCYki0UtgyjmOxr2/OmKzoxfXO0Vnol8ZmLl2b3vRAx7RLCvCWSW
skJMzT0/VXoq+y/VUhSDs3eXVS/q/X5DIAq7DrfAKhibfvvPnNVy/MZ7bVIxHN4BO28ubtVXEKQt
IiZuCRMP0u6+YMzDwBORC1kEV7eVbhWupbG9zOTCeaDVEjTWLahb3288ERv5X/iK1ECA6zqAnsUO
HWUOnIq7z9kcGD1lrXva+2gCGzJ/6eQglJP0GX+OXxViETXIkRHvtCv3DSDUHgwg/9cpztW2wpYO
1noeoLI+o5Kg/45dGGVOVl/3zyF1V21UAdLef8ad+Vs7m71j21l+eO1cyUYpa8+JDQoWsONj++CH
HmhGDrniUuc+A3lWjIU1tFTbMdGkNSWkIoxZWTL9UWGNPwE1wsdtj+9gwHA2QtO1EtfCZgNJIFBQ
sJaHz7GwOKtB+xMEZmtePBZCasYT32uHzXCZWqS7eX0jSy7lgxqOAtuyIsXf5yf+KxKmqLG8jmrS
+V14aRVW8ngFFiFny4AjXqW0ql+81cO+P+66aZSYqtmLJEJyRNMKyBbZKhvcGCio4+5Pee4iM+vQ
gR3O1YphOmXN766bJ+9aetOt+nSxW5+5frM1HkkdaJV8h4O14dzGkqz0KBKY6zKGu1rWf0KEsGL/
6PfZTDhjW7L5cDmbtAJHN8+7XdSSJgMM779BhiCgGJ2IHS6+YEaszBFp8/C+WA8ycG9FV4fswEBm
gV7PJflFCKdJGLc+47tnyGVK0gYLcC9fXtmbMNeZOETPk+SG5r/RGpeDe51qk8QM09WD03I8U0/s
2uIBDiLXcN4KwCvalb1Z6/FYHnhZAcSKCJW/o4ev5ECwS2eL2VEan2zCIrezU/ofCGBoOdlSUd+v
1cMPw+CAvdgrM/OXDgSV0n7r8XtpMZTYdPpnKYhx5XN80j1TS2h6zNVZY0OjyLwsqYvubxdYDT3+
mvKW9onoUmoJcE1MFGav96aZ4ZN+sQbIB7cPiozE914blmLUmLezR/Ze4yKz31c16L4JUZk7LHEN
9OjtrhiVSRAduMIoyt3Qae62BfudzkUktwFKp+Ayz6uWfwsPwsuccjYPwod6LG/rPlolI/0mNqgB
nJZidKJ7+G8CElPmehCsVGjf/J+XB0Ecc4JKQsbERUW2/7Hj5fBXoQtq+zJs/TmQvfMWjN5CF+4i
Qt6/6j77FGsDphLf+4cI0z+AxCo2vwNIyvYpvdj7GCDivbsWXA0hndvF9qTUBk2yJSWIbn7ufKmT
LucX9KN5AzIA3gLOdA+5ffadxdTTJPdxd6ZlIKj22hFrEgpeviCtUziI/gyUEfJZ525poMDhYW8+
bEwY3lhRdkHOhWa8BdNKHv4N00PNVAUsooeR6sNhu7KWMrJ7VgCuNimv5XxG3uQCoqiEfyqPnVaf
3C8e3wRFf2aHnHnbcZvPbfcm+6rD3irTLUD8ZJENkf1r0Fr8vFmIfKg+Zq1vStsdtAVZry4X+pCf
JCto1BBxvK/wdKvyHuo4J0+PJ+S+jx0mgZeByhSS8wMh1S+m2uz7GK0gEb68RbKswxE6h7k1OKNc
0eV8pKXC4fSufPONBG24EH6mDSjvFcqxc0SmwUiIFFI/RcAhMyr6Er+zJhanFq0QlCpnx4Wjlw0m
2ST8Uw9IHrLlc8iSVPWgWVGdpgmxW2mWynOjSNBWbmS+dC2ggsHR1MbkGZssv02yfO8FAwu0SXaJ
+pLsvQpk40FeV50EubEmz956pYDKX0pkp9x2r3Lyb2a5JH+iNYaciWdRy9E0edUcK3icct+3P/+3
khsdgO68HzqeB83FHwViMogUt3JBxFVAuNt8mEBQM2wB/n1Ukz2R6oHqEepCvXQa/y+En4n0W6je
ho9Rrw5O5x4Fhqjfut3V22reXsv5U7Q0p/ddxtAW+tyRycRyaj+gPRxQVoRGTNYwZrgCEsHvswRb
6GgaZ5Zw/zELvPFLNATWq16glSskUfu+Yv4+HdWIwFjc+83E+ab1JleNy1uzhC2zy2nbnD/T29Kq
HBdfPuisnmm/qRP/j05MziKBhxkd+vzvg8EGoUVUVzjVhhRpzWJhgmyikkrJTo4H3YBmbGEd/rtO
xwo0wjR8iTNV1vmDvGSZpgiz5BvKAx7/R0BjqLNBZ9gA1LKq9xbN1mVQqZNTc04HTRlcCrctn/TK
949ABNccz668Vzxd0bYIkE7lHbetBhXxJp4Vf1+ppe09PrHVyT9VBPCoyc1Ws7XZi1qqgTQJFWzF
sklXFxPhewgcSWtTiaUMIJq/7AR+oDRfEIolazqsmfbgpsDqJcsUrIYBnog1pQK50uLXOvEAdEMi
5ZW5kZzSi8rE1QX/o6tVG7bLHi+aNlKQah8l5ELpxz5LRfwse+gXPQcQpSvwv5gy01FVwiEj9H5C
Et4X+55Kbotln3ficDMd3Xs3L4+xcpCCRUsS9mTvDeYH6ukZMeUqrmcBxR6hlJQtbuQo1ikYRwFy
p3xNH++Mf+H3MQ8oEMlK6b7y+4f92WBnic6bD2hsG81DfDvRdgKlnT0o4zpt/LP/oCDYXoLzygIC
ZtoCNgj9TA8OAIsmZO3z+kGp+QgIxa3h+kg9A6Z3Aqan7Bga/vSlYJpqVGOoJq4FDfIq3o1D8HH0
HoYzF9sViSNZmS+67miLsfAup2882IqbiIN021G4DOqTpDGI5z3fSNcy6mI7IFFT4BVcn2EV4M5w
oh5oPGKbmyQ4fWw7DJbJZiG4mRmQ45doEmLtOfbV7j9d4Np8YIaJdPEP9Ecx4SCq9a0AmPnIhK1F
5zruKF4kjsekSO/QZ40m7kKxnVCK5W3qixgwtDlEqRt59Zli1nx6wG5O+/DhTF0MmyabL2eAj2FC
DgK4IirYc2AdzegG+3jtDCLrMjGzm+ZQ5u1hsfspdUHpn+r/uvy0GPBHPKUTH2dqC+8PNEB9gc1w
8RAwkrK/h7g+eCoX4tjupuy5fEe+JDRCuwWDq7ch0YBblMg6Fp6E6UWryuJ2QZO8ZsN62X0Er05c
azK4nWb7L1cXvgwhdox4fCjU0C4ifklgq15xS+O2geK9F6dCzM2d0FsTfYG1bVy56SgatQtpD4RU
Qo0/yxxal4jhyyY6EZVFWIsh2qu2LGHeLdLAWOUsd+u2MeCUJKadkNtK/xDa/+bsXP9SvvLHuzuE
qzFWlt40t6gJ99EFTg7MbAcb+vMAQe1/RhrHd0+jh8SVt9Hp/NW+ab1LglsG92nGJW6OEGOjlpQk
PcD8D6AVAolWHdSzX/oUeevmxd/HNTGpRTSFzts1XaKtDK9CtaaoFT2RsLK2tNX1XIqQxhrwMCi9
VF6ZsiewaEVikrHNpgU2psIN2Nr4G2vd9EFl1JksRuDv0H2wGtMj5IsjLwz2ENuhCFQsePiREhN/
L5yDQwZIO15NKPplBfh0ouex7YA6bObhcddzjqIgjBtDEqxmg+unB2dB++zZnuD/UHd5FzUdeYZT
Rrwul4bN3Tj7KfLXingHtzNZvC6usQXbJPN6pTwLiNpmbmLSBEyEH1uK7B+QlVoyyX3bbEWmVzoh
R8dUY6D75LE72jUmjEVa/UNmjStF2yKoI19fE2aKmaI1YDmia+beO0oky7o+IzBnEAhoVWSK3LVi
6xfQHD3uBMwZAi4sBajYso/Tlxk+aWmg71YIlNoFTnUpwL69LUzUzbybBK50Fm/867kz1RZ3stA7
Sa5tYLt4LIHErp8i9WRE60XOcb9ujKY1g4J3OVgK4s44m+3VVU/HSzU0/bI3a8G2RmlzwGtjhkQY
Ju394+hkqobMZ3QHEqqDEqOOk+ngJiTRvqIxQjlkKvKOCDYPbEIsgaROVFQ9RxaFSdg8uJmIAK9D
s0lOui9VVuPrvXahy6igWadYXeUy2QPZLhvCMXP25Gm80N/vqim2uFFJNZpyLrMNGI4EwzipJkuO
YRVnFFBE/rdI5cn1dD7/Ui7Rr0FDLgjXLjxGBGy3Qdvgv88/M2kHA114Q3ys66eGDPPXHgpZuoqD
HGW8pcYsNxiM5dmkFIW6QZqscLAazj5XJRhSDygTgr/6vLqfMmlG2abvP3idnmt66HnCG0BaV9HQ
Olyl3CaTn84Ncrh6mBuusH7jhatvLvDVOVhcW6G4OXFqQNaAxqVzcX+f+SndyrRPrYPXfytbcLTX
ya2/eT70TyMrYOnlq53O8q6x7fM/JMJA+qUbwjheVbXWSP/zDJHJKw8bbkxxDGmoRO2QgGB22X0h
W3xXKqCZureWOXuIPot+KjAOTAoKrbzQ89QoV5jA8jmSMER5pDNyqnIDYdsDnUhfcLuQa/q+/QV4
UFZRKOstXgubkaf+eaHMHLR8Qx1q2BgzoJwhQM6PXWcf/DiIqVsUGprgdSfKx63KfQ5T1gYFPVUy
Xb6b2qA5cfKl7bXoL5mpRjRAMLaval5efqmXM75dVkcRHdj/eQ0IqblkFUiKV4ESOzAXPpngxkJc
ODAbwOutoWKm7yiqUgqrERe/34pVuWzMaJAqhqU2Z9Ab7vp8WNDZI0RxJZN/lh8p9R4yjEbmzM4B
AbtUHREVckNEAI8rH2EWY+ro2DwcMRGVVy8td+RC1shBOEig/acaf79mZkMpAKZBt5W6p/0L7G6w
GaHmcOGwxTW7XLJnjzbk794etiU4RcUTg0zaFoZxuIccMb/pb8nF2FX8nWhmzctogLOQT6vACbYn
aDvXbJGMKoqrw5/94WOPza3Vj+1OWLtHcnugc6tL393vsSYpcEPAh3tEkPnzjI01xuDGJsvFoEWr
xHN6QLfPQwP3fYVGBTSVbTUlAiQnXleB2/xNTQ2MtpH9rFE2ARhF4jAAAow8/Oo0+kItnyEC3ixu
7WeGylGI0GZnzpJ5F+cQSS8uCRATN+TDaA17HpBswFSJTSpmSqmahbsb9qr4k1T4j5gprM2Ipids
kHBcxak5V9w0n8ZUS9hNj/ETsz34urwIhCvfs+uH+D8G1+dxALzewOjE/Vd7vVuaSi62djNMmsmi
gwN8hHFusO9D7NdGii1U59J8uT7WZ5yhsIArPRpRQ1+1028FKiOuHtrWyIDoNfxPxIgM/7pdSIpt
/xozVDDjmgTAlb0GzQamCVVPLtAsDJAvLSh7qN38FszbbOjMo7AN1/w2QlcAPMyVf2CA2TORORxk
dS3BZprW9+DornwNOCcw7iSaZZIP1g9AiJDxZrzo6WOBd8dd50nXLBOLVkK/usvIcFIeUY83sWlu
G++JwszKXRWImlQZStQ52RaxXdaBZG/CFUK8FeqsJwhNUuCbt2FDFMkfiFKnY5OrGfKlX53pRpYX
rOX86UB4FnrFjxBFWs/ZMmOWR9Aodruer2jf8sLlC8YKBbOSi6fBO29Ujw5v3vJ+V/5P62psa+8U
LqlDwiACJXGZA3YtKlHWRKdi1Kzo3y9ysKq6jR5j8C+BsvmHMza2wl0tP4IT2Hgsy/q3WTm4KLZL
p5Enl03Pq8kgRyTxpvWWMqOVxC0U/5pY1wy1ws69YkC2EHZu63ekSRY2+oiAf9Mguzqp4FT2b1bH
e50qlR1hVEpZg+FcMDIFkwDRws9QsxNPpKPvINWgAWk+/H2EftiUoEiKw/WOsXqDZvGupBfn5fh0
muj1Ynkw32HPogSMuHzitpXcPdJRqfK6xOCSmkj2U/87F5KdZIaXfiZNn6QjWP0NgJ96Kszi2cPS
GTSdg66VYEcY+1PMwbMP5LgD2nQOH3QQ/UuPGfe1ZZNfXMyU2DCpQQj53C64nSwXIOcX2qI8ohte
z3/hQop0m6Tk8NvX69J6mLP/UboKuklr7VqEhGKhggMoZB9eqo0z9IGNtW+qXrfKwl39yy5bcTtF
+RhIGpP7Vo2HKMvS2fcs5dhIrkzf9wd7MAE7VAV/iPovriZZLEb/OYvSOsUB72UH0EJnv4R2pbHm
MowBsskD7pch8OWRi/pR6DNX/8D7fwSMzJbmP0bOGN5O5CZmtxzB+ASK0xZcBM/wjb6mRC/oZ1qe
FvOs2jZ44JkmqIpoCGjk8m5wtb955+ymp6GqWLSUN/w/vQ8HZav1DWkirxej3DFnQTBfPVlFSTWM
LK7Lv14iQaKnISJe9rfDf2nRjWjbP3JkThZuf443BmowafBhMCFCodAv1qTwI9gt2AX12oFYQhyp
A9TNyosp9R/MsDZ7Ccnk71LE9xw8Slrs73DxCtFWuTMZhtGU+hR5/0dOwwKeBqqhEUpQ4pQkmSII
9iXHHaXPau0Fn+Jc5xo0ZDeFeItYdSgITf0XTEeckYyN6qDuR4Qv87jL7kXxtJwYLUNgZ8jNtPpb
o8bQvKkGFmGZCi5GV2kOu1yyeUkGWtao24MagFyaJ8ibJPcG8So/kLUkWutO9isJ8j6UQP3byGR8
FYHd/m0dKRrd0eZTTptz2/ahUn5jUrp1kiKBBAv5olY0WlnkhYux4vWPzfskhqqD9oKnDkQ4TETX
1ArC+XJxFp01Yq6jiqhfBUgySUhbDG0rrFeIq6HD4evn/fLHM+E8Yi/dhbXzLvcwuR4jKy6l/5Ki
xkV8xBIYkye2Obq+qMItLcNm6APuILNOZzPTqQC3h3WIxSsuosxSrVJqT32Cp2Hgbae1guY5v1dH
3ocyAUKunLA9PanCH+9+h+NSOw2VM01/HQll8NlwRq3FTPJv3sjUOA5Ua3V/Q6q8wk5WVziSIOWM
fzWLEMSZFN+f9TrIK32eboDWCzOGdE4SUdr5fwj/Z/yhmztasXzx0Z7RWCLB4uu7JD7zX6R9V5N+
e7MGOphL+Yef1LprpV3xg7tNMtL81joK7/O4V/MwWJERlFhApdsmRGAFulLtuceg3vflVqixzvK2
hB0eZCiVhwnf4j6BqoKYywBRYPtfu280wnYddhZOCSU1iLjyast+OMNR4fCrcOMxy5xqjgX5Il+p
OtTKIx4OKb+H8jCyLNLqCmB01Ixkd/ODoTELi1u+Fb8w07w8jXvhrmoI8EOBZ/DCajm/X8VJDjxm
5WufHSK9mNEsJXUqqp/XtYTSV4rkxeg9RDwLLXFUB32VhaZV2PDgMjZH2E6RMX49zEdoWn2cTlWW
9tabwyodpaFIdhojnXUYr0dm8FBWo6dATmShUyYHRwdBOf52qW6MDJdY6K2FfTGZUlLB8rqqIpu0
nH/hHMcLEXEMFuZishtSmcQmScyw+ejGk7uOmGkv6dc9AjtXWnhJSrMtCCoGOP2BmrCatTDtOiux
8XbMSav2PP+yml5eSHX6oPrZnG13jWlIuEEfzJyRUawTdXn/wcYvIBtbWFVTBXBMiVkXw+Du6prA
JBYEGPumqSFVMLPn/ClObhoGIqJO/ai+7wOpf5winMAnGcQCYWcJ16RSnz25Zu926yeep/IoTS7z
OumDbskxy78E4FBofu5meqNSHQ2IPwc4PLfPJ1oIyoSgfL83cvkOUXDPUSI1iydgwz/oQ4VK1lf1
QYD+t7bkGAls98kOP8ESgV30Yv03KFOKK4bUiS6GVqHeAJ5eBQeOcEIYbTPZ19ykcf3KjxZTkCW2
HI7C3ykrrWrlapg//iIPQrmwD4Hutqg/OSuQPSAJGnNOTG4R/pDpahjDkLionn8fkXj49oAaL7JO
g53cSyPzN6OG6k2J18pYTfHZWw/QsmebYcgr4UCy+Q58oO6cCwAvDCT7qmIQsnbnT3DRPdD964fQ
3gK8NKNI44fXoLXvcyalriQuOTQp1QrjILzBT7JG9+Lsy+ZYNmCADbHhyrZeGLvf3H+/+VK/aw9P
BLVBuOKEMp519GtLxyTH0DSw5VLDJDofzRMWmiOv0RGL8DaSbl5TpwOcrlVNKBE0A5xUGCRFVrU6
QcUuVM7vbgwj/V6SWThgsFRb566Iya3ZW6z5E9hqLrJOr/b3XNWHjZORFbWlX49h8HA8fmAbeBC5
YIYri7/F+07oWeu8c8wL2an5ouIeiHfkBfPT/pr8NkPeMkOVs+tw+3iqXz8HiJFfAR0O51gzQCLM
SSsSM/vpVFUQ4Yh/QJXYvnXHNS273XrMz5Nm46n9Jth6mL1pz8n0b6UXZXEuPDLHI6kaeTs0JIAZ
gxVR+wFucSO5a2myXkV6rVzCBi3TS+0w8A1nc9rQl/nJzDgy1GR/M/8IPnYna6wPZW8tKBndasGg
tFgpFKn0hbeYsDQkt4iGbsxJSxqySFvXoE1cGKRinEvTf2M7EDzo3bGx/LlWrR4RODowmSEaXB1L
Wj3n3XvlX5TTdMAH8uKFGTZE4sf5tEopNkszbtBCXG5+NN8teox4Iw0GFp/0ZCTcVPkhinwmkLvO
CuTlxK6RqA8G8awXO/zs4Qn22KBBehykMcv7kGJpdUH6H/ImW0pmYCvr0YFsQklYBO1ps8eZO0kp
bSCQkIWX/vUUXQ7dTNIWSTWzIPqVxhblwy3QqNt8KJ5cO5cG666hUKJPt/Xz6JJeIaa8JonFqjOc
HBA23bJ9TflZSA1LTdTDtobsKTxMHPrm01cbBodaMn0JIBYB4YVjkuBTzL0ARpFKsekXK6X8BYxh
jCVuVB60sla+n6/siJNdkRH7IGT4zG+sKBQNk8nto9+jx9z+7SVhhQzPiXNzgC/gvE8MgbMZmPOS
+LR1aXF1xfGQqaViTS8djHkg/iAE5zM/55g1CmrsDrb6BIhH5zguyx/biYqe0BRT6pdzsOxzwXIt
ROgmEST213VYm+bD0cs0mr3Kip4ujAzRw/4pIvPcozwHzx03+YSwIr2dkMw8InPi49iB4FVO+P4I
UVfsk3RG0N1S/UbJwB+YQCB3ggGJypNieM3dyxVgNjjLvugey2S+MVsT8IoMi0ZMquFnEMhnEmsq
oN6yB+EMh2gME0XvNR2bdBNCKfXSyqikMk7uE/J7d5HquUYT7mU0J2t18AEn5BXpbtao0YFZ0aAT
nemRS8eLh3SSItFNlQ58PKMAwUk9YKbrBGU+EL3fg7sEcciDR4ejF4WdR+8BndCEThXtzOr/xMEA
U40ORS8Rab6bwCEdNwcIw2RpG/Z9VG6i+OD/NWISU/rfaOF5wzWDrQtBoUFLdBWywK5/heYh3TsL
WmCw4bwNVe+3VbOvgifJXTk/lDpqg2nfA7el+Aw7K8AYkKeVFHJZqbZ3y53nCLW9JNpMKbM1NgRs
tCjW7tp/kPseYQUbAxkPDYVqdC/FB6lb91HtkrzaBvcl6YTYhYlYZ+sQCXoFatxXAhlu1MUAdWCv
Ivi1wu0c6xoHRZWbp8cVIpC8bewfJ+g5hU9eHcwl+ePBfxzV6+tJwBiMxWV21lfMOrVJ2gY7Kkwc
EoNVMeGWYerCgLmR4+spjDorBgc+4J1m4qhAKhZWfPalXJZh+Gkq+2VeZ2h8vyMYMQpA9gZ0NtQQ
7mGEr6LW40JIVucg0Gezb9Md+FO6W8HCJ6Ny+vnsH3E/X59kXYPg/2qmAc9xJo+bXkANHnP39Gt4
MTFtB0mFlWDTK1HRgjih8b95E/As+LOSmWd02OE6Sq9neA+17QtWXQNoPC1W3pW0OEhvShCdhjsv
Ut8L138R8RrCjbjDa0lttIaNimakXmz1kseHOv7+ZgERcCROlBw76sZCKZlPANBLi23C/02uUM4U
w8UpZ+FWE/fJodZd1dvS6gg41ZszKKmQaBsSWX5cNqBL44KLIxD2daTMrmGHb6TtS+TQguEuMwoD
PDjKPVdARohYMi2lyvuRy0DLKK+m+I0l9aZCCCEg9gAWAUUk8/mGihaE+FfEuLKp6kkjDOPe08wB
Dz1Vhf/2sX8K04mk8i2uM7hyHYp4xLt0wXJXm1QGAz0Cb20R8icNmF4c3qXfrfO3OKksubauPz6E
F7PRWVW8vhFhEEBQ58XJqmUlyW/cUHu/pp42Jy62hoN3fg4O0PfsN6Ab8GQO9yDX8mdM5N17pxej
JVVOgGXlfx+tRn82Mz/1lsbPDYNLh/Hc9KNK43vWeBzqlfzrv92piE+3CwIF7E1oSGYYUX0oIASN
GzF3UmfEWwPst4L8C1lpPobVOkVqCtpDJXsNmNEPla/Is3jieN5fCfeMKl2IbEHhMKN7WREgiS7A
H/szyFxSLi1nOMWwEldUOQgILByjyexNQVnJ4t7xblcK7UOzWqADdO6iTiP37HTb53AZv4nAy4V0
tpU4S5haU4pXdjlqTHLXGIq+GU8cal9faKEAyV4UqOb1DjbrCZSv8LBtRmt7tzoiHcZ2BE00maoN
XC34JlGEwdtfInrRGG4BRIF1pyC536Vw+jxbSL0U1Vx778EkQXf15fjcZnzHLk1W0pCbvlVNZ6Mm
FbuaQYiE8CHDtC+UHem7IjOQG9CPA/H83jqiIm07QWGWITagyCxNLeXDRXzS8EjJxicCQ/zjb1E+
4k6E+UaEFCpr2VZbl1Qo/0rANBXIxSOxFV4rnVnE7Ry8aDM01HdWU9gDGn6in3JPrpxpBb+bUjWj
/7AbYnpPjmfKw6+KBvzKmcdNwaWK1EzM5+z1GPMQZRY01ghj39bfUGWB5BkKI4QkaSWfNXLYD/9r
yqlJPf9mzScxyX+Iouz5uamG+6T5AK3wWtQZNrs0MsFf9cTJT4LvXiNnvqQ4LI2JqYFvIQwjAqWX
02+Zayk2uymFRDujhKyUXcPGRauNbOZYl+jdEbhU4EtuN2bn7BAdnBLC6hxNU8ubITxKdYOQLNqP
AqlPF7oDctmiGfr72PceS3wqMcmGmUipMBQALbToyFgnW5+ym+afTc+/GPxKAxTRF+IsfCM+yLqu
uEjWVKa+rci9XxXqK+N4CR8oGMMj5HCPl6fdOdSS9jMzByKuqiGutnp6VEZ8yYoHywptSa1IRQPy
ZSnd5asVE76GeOWLAKgf5aehUxWQOB67zicuMiluD5ZdWHFCHy5TQ/ZRWgQRE7elDBgAyouZamxa
3fn0Ve69MGd99wnE58FSxtsY4SHVPRe+BrjKiDZqHMksV37zzr5eMipkpbzh5737N/yzOFOlpkEL
69P34tUYxTYdIPy/r0JOkuWCxF8M2/CSKFAk1R72IE/ZV1/7LIdviW+S1LC99t7y2Xovpr3ur0Av
1sZ5u0Q2E7q34pqcZQZ+2pCGo1f7Lh8DwKieGF7gfrAH/o+qjSByNGURPUZOL083AbuuzjvDoxn6
nnGqjbhnu0cyx5xE429nOTFc+KLKRn3w6O4XFRnkYN3lMwtUJ4cah0X9gk2iIXkmT9HdYK0jDZKI
arijixhBPpgPfuRhAjrTDFMuYAyFHmZytETRpp56AcGs7mBtWfQp7x7KBWgJ+Wr81rRKM0aOHngx
Hoxaxfwxh/hKDbyMse476vRcopupfqpreQIh4HXo1BMwH+HXGCHk4CqueEijlPVd4b52UJlf6B0i
z6M03bcDLmWF/rNmCWEhrxN1xfvpybDLZOVHX3Cyftc9hHY1ZxHgMnGTjG6cfpUB5DH6mtJBkIYy
rK5at9HUqfiRM1C/nS1P8NTNzPuIdLH4JLytZboQnVctlqmQNghE29Px/rAIZYjCIv7zufUoIwQo
A4Px7DWFoKfUuedJOidCHKXbmMJAcdHZieUMOgmhV60vhWdZUfGQzoFeP8Q4F3GkcAngDAyeiOTc
SrfQdRFKDr0C3Q/dXf2e7GACba60ipFXOofApvOZ4XD5POqAVk/gj5c3PvsJLjUcO0ShxzLtLfoA
C0aHlOL2RbCngJQgpCSIwfuEOqp14y3EUvohm44LJdRYeRublPDSdH7odyw6esoq+4VSCe+MFHha
BgcWzRk50ZuLkErK90vUrNZr+fu5YPRtKBPBxRCYcEcDKC5h0V1sHcUUMiWt5MGVf9Lk+ZBBDhTL
yb3gfKHm0P7towjEwj2qgY+nosGBo7L7y6riJzfmywuYAQ/CzbR0VZvYDC5nikqnBC/tCJsGkqx4
q1Tk3lt5rDiIahjW79FyVvlIHeh9+KzRvCcoslliFUs30WMXyjqCo2f65Wkm8q2VuL9yim80vpJ0
buOjeJQZi+0lAE6Cpwcc0W7P+fIQCLmmwqSaSzQjTRg9hNyLzMvmstIZMCckc3K805S+8/1HwX77
fjzUhkKlrDeK+hHRvNHYy8LMOomyEfusYAUhwSFeaF6p5Iogzlu5xBdWubE6lrTj3953arvFS76A
6nJcCKz2usCHNBp+oagFtC9R/vtev/41WZmooKADySJ6AMewiuOWcIdHfhoIVU1blXCjq+YQqKb/
MK6uHKvcYizjxW3Q2UUWaBYIrHAjkHNjrYKe3jlRR+NfXkE6NJcmLkLtmN13gJ1pBFaQj04BaMdt
BDXVyPrKbiuU3fkvyK7TRXiGcyw5qW93/wJZW5+fpv/KQ2/98vVxN8tUAcaLfOw1wceqpaDr00kt
bKg0VzqT+hRilehAbPuq4QWIXuHl3MQVtF+QSKu3LoqmyVIOBD9NH8Nf/bdav1zDzc8jTYyIeM9m
myLAoitgQbU3k7xW9ZMKGJmL0aFoNppKnfQrH+PI/4FzeMUXKz3/GlHrESBI5HO4/yRybr9rz/tu
ICyQY4kweruU7/+1ZGwZg4LDszRtgT3Bu+bR9VjnM5Je2FxeT+fci4KtG6X9Zlk0kBcooodXCqBP
8wL3q17wlPOrOeUgQaCWUEl7mgUy+N26oz0fyY4pApewyMl6FxzQ90I39TPBdQv1cpqgTwedbLMI
Jp9rtxejj+1H5lcQgtXea7ONuIE4taZCkm2I4x34v1DlQnQgejbaWl+TEiOCl5V1eFZWGb3k8umK
w5uRMbxQwTihjqFHBzFYboT/kC+UoMz9iX4Cex8ODLNOn/fqzaPtlNpGK/qzotC9aJW+zEj17/gr
OXcWlWazcTyvkPYU+Qzoa4A6Pjguxs+SZ2VL1TuQ/WUUDZP1H1cgymm+fn1zy7JyJPop0bWFRT0p
bMwwQituTJMW2R4sXV2jiEEAfdOQlUDpqBZuJ3PEvosZj3mn0eSpnyT/Xh4Uh6kcYEuOAcEe0e5l
SzUX+gzR+XqonbVGbncoMI0WotSIdNsPC+2mfVs80I7/D32eeUyIzwaWCylWe8yfacegZWzR4GtX
yx9CDg17VbeYwZ13buie2GSHJacQBjbjrlmIVlOd/5TB2rYV7NHjZZ7GCMO0GnP7dxX7T3hpKPCw
8YQts4klXAb/L4Gn6uSVC7axZELT4OK0KTnZH/cJn7JHVEar6GbKnhtiJWAutTvEYU6wPi8P/7BC
wR6zOyRAMrnIRHG64AYWvoxfcT9CDrmKLSaamG/RxzFTl9wIAe2pa3ARsuu4g4KLlyw+7/hA45ey
06OCUKKlGy4J90RoLNn6Uxt9xB0rl9YSYb1gviuGMFzRDj7btanj1est9um7h77/MtgmQ6Pcs1LX
I/4yAKUnIoatkLFlgyHchW+JQbP+6QpW0hcwT710Pt8y7Z+cI5nBybB/m+aW3H6SBQAvq0nq0zdO
j7cC4jbvwkxD2yrvhh2TvRLDWdXkx9FqMFg2142sXphXS1ySkYtZMyEnLvytR2aYTnts+KBG4Wsu
iXqPb1MtJnG1y6zgqGITqqDrKd2tMHPmcbVaB3oqDPp+QMCUiCJ1jVrzsyBZ639cGAbdq6tF8qDr
oblkqNgBRJXGtaXEYD7pAnOamNMw8MCfy+VmrtfaNP3JN2s2gLEmWF2n8V/EL5cpr1/sgxZguG84
h8g0EdWZMdCaOBI+DzRnBiNQm9rFrkd58t7oc88yeClNWWFFOp13gWZa6B4+glbHcHPX+GXKM7Vz
QlfHrDzH3JSxatJerVdydHmAciZtxr5Jx5XnN6DDf704LkD7lCq2WUnjSD5ULnmcA7efFPM3Tk/E
OTqzFEpMW0Ik8JniGIbKa3c0uTRGs1reCo8yNlriocvYnHxddWWq7Os7E1URe/O2bVnrU+c9ShhK
mXZN4jeCefOiZTtIBf6NylmaEBp5BfB1t3JZLk1wuvhtPokRWoB3tQcOhYdKZ7yM/7Y7DvemIXKy
R3+MdqUc9YbjbXadRP65zbouwA5FGQpbGxFxMb8QbyHr5oEGxeeRSkjH+JIkQ3HI91ekxoheTDLB
2NrgSuQcCwJBCfWoDRwi2Z+9f7/1Ev8DPBd0ky+mBjgpXHvzAGTLvO9B7FURwTjeenqqc7O7nVfd
Oab0MfJ86J0cdYS+PTHSPPjoKESjjMw3AkL6YPIxJQuuLJq6LbtjxuQkh3cLyOc2iv92wAdpmY5y
Z2uRE+ec2Cnvx2pgrfBfMH/Jum8ZPWa9rXCi6lHtoX0y+4zgQMVjP22PiBCLbH2CBbg0R4pzbv/u
YUZTeXQADo+BSfPFNgOxhZ+e8RAdLTqoB18fIhnhgVp133/Rg19IwkziVfG6O5rgru5/GJUfLuYR
jPvgr4ii6TrhlTBh3JD10+z34TNz5ehZmkHodAurajLuLgm9JmUrTn0JJcmm7kRI2TDzQuIXKR8J
sjAdNH8skQrJCLPRLLfkVfLHEJ+rF+RKdPq3ngF4J3RpII+kB9mAqMVnmSsxCMSr6ymS5BpMOyDu
mmczBYnWKtcjNPgWevHhHDJYvEAdWebmNo234wVbr7I7UA5RoNmdYgb/ZFBXrRCFvvCnZivovvLh
d80UzbIHBfkaBgWjlNCiuLTMPo5KnDKTqZkLnlc696G2+fQQHTNeXubrYheEX3RrBwveP0/XqnLq
8X+Q0+t5Ooa7k8bE/qgyMmfQNkFlgtYTaK3OOnxVJA7weSj/BmJilRHI90Vmic7jTu2004j8NWfs
esRRLhFBGMIZOsmtcdeeUVpy1hohOsVCRpE2vVTUoMJw8ki8gWdW5JW+NHKrZ/lI0i1GQCoRgD81
GpsKOEjczUDvNCV10g3AXyNW8RYZaWYCtEoOstmFpPXp8L1VJdN1sV0xgtClGxOZ32fk0xkDUcnb
Xur3JjsNQ3jNpIwiemUq8+p0HUzczg/5uo4A6pCRoEFkvpRTKKeyb4ox7Z1da0h2EsMfcP5+j17X
9u9DrewhiKL1WldAKx83YFoRDsg9RnW42Pf9YmXEzeYCD0/eUxpx1zn2pwgSW8AaJHN+sl0geMPS
vaH1fIjW/m3WkVmEjVVQm1RAqCLDAAKyrYzugx4ivLsWyiKff0yxNzusrcO1d4yo6SdLcxTPdJr/
aI9v1qneLkR45xub9c90YM4JYOZYwlU4/6XbtE+4isz5XWg/kzVS8h/hxkzA38QWbaoAjY5DdrJ+
jLHD9k2FMG79leNQKqQTXeBIqDfVqVOYxct7oWIUeFJnX2gYFnAcvFzKdIhw7o2fUekazwReR5eJ
t/RnfKZIuEohRnX+WAPHt+FyaxEdl8V6ymjH/ZfNZEVL6gQqv3GRCydSo+HcDq5g03AXFosf0IY3
Ej/sZKrntS76Dg3CTadOhGkelWdyVSY+leRx8pxptTk46PbyfyXk8vna2FPndtKx1lDrg+BMQv7i
yF1dQ3R2DgzGCgxyzadEMQ+r26D8OmLWNC2jWgA2hF7aTFEyGVVSAgCa6PxL06SuYsRGe+yzFjcM
97qcpofOXQYS+idGaBP50zadnSxjdvCsdacqHJETGC/ttdXxZgmi35W6c1H2EP8ml8z3DmGaZT1B
gUTuWlHft8C6jL2f5TqBxjV+FAL0el5DUmQ4OyMoHcX3FGygxqPWZryhJhllYD0o1Y93cgzh24b5
Ph35ynvDUYGWnalFxVMqN5J0p8hYyqT7FJ4aYN7IWQct/xgOKYrkFozrUeAbC4Fv5vxiD6uSyi21
cIH2ZsOmHvE2u1jLzPwBp4vjEBxv6Cc6+bHYg6BKa/fpqY2If4IzeII3LrPWK3wCnOXgG0wJHo0N
1rd2sn9vD6KDr5xzDFgU0UkCAbkQRJHe+6WGvIbRa9ViEOzkWiOGLS7jCXtp3098l2sY5BNbKUtM
5RMDmPZ2ic+XBfyC/dhmDoNN+/4TTChwRJSglbstGMAI1n6wjkKnxe/KjDvvgV1izyHHTj4I/6iZ
KW3v1JwqqDZenuxBrgDHgadFocBjBxG1o0cdC+Q1lDY2TiKLuxdoDxeu5nZF5xhFqS9EwNizfwEA
fnIewwPTIrMBSGsPFjxC0l+bC4CgDJwkzdA8tJCewSnSG6IttTieaSu5UFJldBZZUsFMKIauuTZO
xHcruFxxusVgBHLURLOVYOaOO/hFZ6fiNrUcm/RgCqVcWbSJYehcIz7UF3xQwyBMlDM+9TGQuP+k
J0uyMhHjm4j76nFxEI1+YpkyrQnccRf9CDW42pofWLPD66DPHEjha6sswB5KXM2sorsEUy8uluLP
4gNenNV/8ypJ4uy1h7Onlp4CtX6RrV0/lBeWi6Dv6DHSB42FC8mcy5dmjjOWr6cHtLaghQjI79mj
HuUuSWW8v8cwfn/6x1eg5KQF4iM20SwK74DR2nefHQ7fMsonukzvqKxkWUxyyir+aJBiK1Sv7gKP
0h9+RpQ9uxAYtye6WkFO2ciLNyYySUAjIupjyJk2EeBbIrskW18MhLdZjQ0FI7/N/4XhuHOh55lc
DR0IhVWT+v0BAklOeOij5G+JvP0DgUMIXxj4tvdzGFfYOMBqJfiq9OO+/9QHLVL15vHdXeiMGM6Y
dm7ipPbeNEMPR7twRE97+bCSxq4VePYmare6uM8F276vjihruEoi3z1hk7V5o+lQa1RPV5HY/b1G
zM7s7X3dypKqGGTJsRF8W+iTMK86S4sDx7QPYb6vjAIuM/icnmUYrVlQiwAqW8ULyAqQup0MxQpa
tegEDd7DOnv4eQQPqmEWtmIq1J41hfIfqN7g4xuyZGtMR7qN15ysrWd2bzRN5H/R2E1GEND+PKRJ
MEhntXvL1FHSJ3NCR6MkMhlnLeYccVtfz1UHslrZHPKvr7JEXnH2cXgTo5o/APuOTjiOesJyGGOm
ywY6I5M0joCec62ug7cR+JvY0Z8wBunLwuOj5f2fvar3W/4HYvzE3bayMADTT+g5tv1E5fgBglye
1ZQtF2gszM8h1/NT7ADPL46ZQ+33ni6BUFzYz7u/RD9qZfrC0IepbVphsaCsju6VHx+DRCN+HhCJ
Ap7VpaS+Podmcf7Iv0MbKOyMkL+FrOrgYjpdeAFsqVqcmij03l4d4/QveJgm9+l1vlx0BpUZNtod
CMQqQIgQM53sVbKxzehp8ban6kLKDebRoduEtlH/13MQaPeWZIMJF3WBAMzstEiH15+ihJovgAUQ
LHwUGHX5xNDZl3NqAg2v4QGQy8xsTcKr8vyvdmPBXkmFw37kMXUy9oW74/0F41N/JJcx3710D2Aw
UR4UyAhSqRCCUgHP6ryj4nFK1KkBanz9ZtyIjWSQdXwfJXYDtuV32PXQItDcTpecu158RrlpqObQ
n4nuOhbh5vf0mSSyN/85adwNfOM8ZruDUaL+i5NhnZuW3ho9cfW4rlW/S2ddklgYpGt6HX2xIutu
y9ryeQzQll75SbFVzaonBJkHvST6ibG04TbI0WhZyysKTPXqj4jKJ28P4KBunaTaXCK9FNIaZ3bm
m2oCHuWWaoIlmr+Vn6Vvu2AUrOFWHiOaVieo+Isrh+yNWh7Nwmx30zItX2bC3QTykFNvWgHOoMdz
cLBuj2QrTj32uxEom+7EYtvlh3HI8Bic/1GdYxGH7z9ZxxBn+p/Xd5zg4xRlumBFD8uOJuRDlNe9
D2W8KhnttcOBIzJ0RfXtMfk4Alym7MocfpSCVl6RPPUw1z/6YU2sfiWVsY8RmzFgAlqj+39BVNCv
KCswfXNroy4YP8V+J+81kW9P6x2tnfgv/vKnQhd/PdE2km6Cp8Lk2yxHUVBI/62tpHOiYpouZFCM
qm3wwsg1kebzHYym0oFFFC3ZbfvmD3m/GWkFkntv8yOeBu+wYNBr7ch0z7yc+cNa0yiVNoPlYheO
1La5dksbq1zZMPrHuMgxUK7+IPiSYOYjnTAi4CX6LWXXZMjlVr6RwBLeVqTC7bWs1G6G5IA4o6Wi
lu9QTJIAVMNd7/YedxlC9Wf1aP786jC2oGwIm+7Q0CwkZC2exMcO9RqResp3PKR15bSubFc/SxIl
GTMfNKjlbeObnLjdg59yVu792wi3YV1fpD4IjbP9qQTZ8reQ7PCfiwxMvxP4UQL8t50M3pZ9NOXg
F7cnV6KipCq7uHlOk0PdRNIUKQ6loHGknCmL8Xljy1eBjsXQn8uQYzw2jDvrPqcC0xC+jjuhxZmx
WLVcl/u7qTLTI8fc+JG/cMA2+qq+N+Kj4lMqDbyBhlg4K2pffg8BfcbCTK59rc+TK9sRcn6toqvA
OXcjTS6P5NNU/vUVMeWtt3bM5EJfz57OUmZBHNRTpcMyu3X0EzgVgPfgnokpNqRiAphdKPr25vh+
5HYqjJMRVz7kGOpHNjC6RJ8vQYCpZm7g3VLYMCPro3ltvEIZJ2PekJQnb5kMO/cwntwd7CIK+K7Y
HnmzekYfY+1SmHxAPJBLrtfP/r2a4ZEffD00gBiPNFbYHzE+BLdI/kbJ123gm/nKQabH5gUvSUla
h+TfUqQ49bvPUeS7GMRKkMSoonFESvp2lMuwOxaDUv2dwD9kP+cfScB8+yUnb1nM2zKbhZ7cx8RP
CfiNtFPWT+Jw8ZsXBmLQYCZI/W+mmQ2AMyNxnAZvsEzrSlLvjVr9PbboltTJ3fJ0r4YQCmBAByhK
+boO7rGktSHAp0/wH9o52vq+w4lxNFZ2bhVRrgwMe5gcFhFkFPBPm6UWfNTgKZEbRKflTZfn5KmJ
L0IiPCVbc/rXVfSOPpq/u7Fio/KBmkEuqVFRIgltFtofy6GKMBXpN0NCOSP9cbt7lPZLeM/A/4wp
1YcgemIgKdQYyIZL15nJhk7TAndLzxEktDfKW9EtpPP9pPw9mZ+OWrC8k1G9JtOO3cQFVxMDEfLr
eLATK31F9glKXEJv4at3tL962HLVsQBOwcCraUCtPnJtQsbVzVjUEC1mjDfYT39n7KV1ckU0XTt1
og9wG+vFiOU0OsOl2rkAZ7mHAXDu6VNx/OmwAdgJsy4ce4I6s4K5gfKpVIliKR7C4kXzDy/8Napl
Kleauaq+AN9dhZkCl7I0BIIaMnmTvvThvOHgfXToSaef4j8BqkSJXX7y3SFvcIHSdDtxPHFDotsD
TWRvhrotiYoyog6bahF+qUK2q93689QW+l9kXUl0QD0rThij6TG9c2WTAzA7nO9OlH5DlJ+J+rhl
fkZwAvjCmSWicKSb5G9vCip2e/CSfFWRvZhd4IVuyP/5NaQdIQo2OblvVZ8ze8vdgEansfZWhJbF
PCo0AbkdMRI4FrNWyCHgLPVDt/0AKQSXdjyEgk/OnLRYuYGN6LWfLOSEqlPw33O/2eObnc/2c/AZ
+o33k/k2ggTKh+pXF7EMgV3ndJX7+MyOorw+hoVbJ8Qx8UsZpRSFO9TQ9CXZDBeEUOL76H1dEpNi
kIMf5cZLwLBIBOmJR7M5SpbIVQDYQfwJ6rMHTLCWoGvqAQdT/Nu/nqeVw+/jxEYLqz0Sp92rXEmJ
BPn1Z4cemRHpkF0lMGNFL3g3R2PS51V9IYpEmsH6p6AN8k5slg29I/qjeFQRBIJylPPfKVZVBe+D
bUI/TiyZihoXVq3O5+H+kxl8tda1gmKZEsKmbHT0LZvIrRPHMR21/vkjYhQqRmvF5dmFXbCTFFD3
mUpkvwXWR6FUMbFODAcUljwJImaJvmSAac0VOa1sXJOgJjU0708xRDSFNjrHFYRWwZy2wsdrT735
HEgNW9Pd5qNtYCrzjrZHwhimkZCpFh8g4VI7kbl9FnPfCnabNcaHqjvdulPD+gfgXei8P/B7Igc5
igWP055hvvV1hwgx8M9LavuLbo3iq59AFjNVT4e/zA+XoNtLQ5dkjF3wtIDQA05Pa5VLGjkcUUXH
vT1/tE8N/N/X9/jp0heYp3RXZMc7nxkZcyXzXVUOfeQt463AjU5xSjTrsNT6/1yWt29veftqqV8E
I9Kz5ssLxBpk5hMZaTgzljFmVgB0vDXKltGnq0cnWkqzI1UScCcO6x9PGowMbB6EXWGTmNckcVF3
6dygrmDsCQ0k6mZvxLwuPhTnTx/Dx8ZqtYwpb7ml9HRz3Z6mhM5dzbfonSMc9CT5WGO80+q+AQ8g
QaY/NGY9McsKl56spgdzgRzRthZsWpa+9ALHUOP4a5YGiZqRasF6BziRnrFWXAHm8/12XlsCu1b+
hHFA87SiKXnAh71bDDr+V0lxe22Fn9UFKkWzSgHEmazQDq6jXYw5B3dhLdC43XukbhrdW4cHI6A9
UC1WHKdoeRRGmUUdOSpJzz1FaSytFecccZ+RHdbdmVTDBzvyeUq1gHd7KKQJFD8IMAlUBZ2bV1qM
VnKeK2LekRjQxSnG7f78/HpKd14oVrJuGdR8Hs5cInGsOLdzO27HuajHIRImdsQ8B6liMf3+YScu
hUo150zuHEfdONjZJZ1obJFsStB3B+2ldzMQangCkg9iFxXtHwjBE5uCb7OUaRXf0GX0lD6o7p0d
c1shZlWvG98wP07QwcCqNcze050NdQCRbC4F4GRKxNddL62TPVMxl4nxj4R85v20nxsCB040ZVle
wjqKiKanesnMw8JByvHBw0lFCpfJqW3y51lw+R0iALv6nY8opafDQ4SBUvLdvofBW4QbFUHKHyF0
d7VH1RrXC6I2qjXvsLTgpLin7RQ6sHxWAwWmNsPSBMVT2KTk7zhPAeCfDP0GWzDHQhji/hXLo/PL
N6q1NwtLSjFYStjYxCkJvgWuQVzWT2sDYJKK2XihPA9YgmooQR+OacCtMEo7EzMLRbSFJnb/wYIo
qTi/ptm13vaBhXKAGXnEQPbWrVNyasnwjMNUcG80TFJNMj0pnWlyKuASWNdAwDQnSYZ38FFSZ27i
N7wc9A4Q5y4ck56UMCpY01oqgHy+CJeUKDnlYWnDG12HBcgCp2HKtS4/FNJeRTX0N74EhZ+Itt6F
Ml+Ne5oAPIMorDQooBELsBAA3ZdccQBgbuaDW5z427x6+SDF8YUzZo2chk6XOivoQi0R5hdAiGF+
prKiR7Hl1zLH24/nsoi0JWKrNWqWtUG5ebQyjWMgVIP2iqIjbVpD8P0Jfee2rgJdwNnc1Dzsw/qh
/CF+ujHrR97HaKEbLI+rA875Yv1wQW9KZ5+7PxsPk86c0/Fu0Kkv0tKM5UrW1k3IZY1ytAnryE5/
Y4ntkhV91KHN/DRlIoRQpi6dxMeURCupxfts7m32NbWY/tuX2WY0umxg75IstIGsHthYhXPKM9js
zPvYr0gI7PTTO4iZgHSBzxr0XHoNt54UJmodeZ6R0vFUZx5dpSK2e1+nyxh5c/qCwtRUSChcK7KB
cIs1klfF+hZoBX/LzN2R380WG+LJ1a1nR8ru91TkRaJAU5luWolUdMuRgZ8jeyhIwuNUD7qJ1Wpy
YiyZxnZ0/Ykwa+2Gz+GWDYFhXvomfbUDFp451uG0yYpJN5tek5yMOq11mKASP0HxWX26KeYbgThi
RC/ERueMBZeC4utizx4C9YAdr43Hj+N8ACxrx7cfnUjn2Vx0k0q1YWCek3YNhB62UWqSZFGNhNwB
eWO9rGfnAU0WcdzxFhmm3YDsq2jNvhT9TeNhUqGYsbKR3hwBWju3fyB0kG8xHSLWuOpQZseYLPny
7gwZ/4YvVgXIoV3Zqca+qItqM6dxNENhPjCxusHUbsGpWiGUr0sTsyiutV0PhvNezls3U3QypQXB
j2Ctw7DMPYcdxa1aRDrjDzKXZR6NfQMctpZ8WMW+mWQXqcyYke6n5hVhVb8nfKlz9qxeDhsltLyg
uAqRrxUrn784wU17WnpmYxr3sn/gJsIQSXHuvHjBu2J5uVY9pkWPFRjWrKMi8siPGwVWPTPErAHg
E2VkZm6JiYM8ochb/5t3OYKzisvV6pY5hD4IoQmH3IGJoKxVAFJX3uklRKXY+aNcGj5wqPHbW2Vp
7mKkwsv9pfdQH4PEyL/JAL1R+tDLlgiwxyHkWodbOHtAtwVJBG5In3muNK66uVt5fLoC/iIx4DEO
8vn2nYtJ/3Zd1jhny55MjOuA5P3CMoH20pPJI9wcjN/rzedEMzTfSwcg3E/Fha8UB8G7HDjDI9lo
4eixWMiu+sq8Q/gTD6O+n/Ap7xd71C8DZlTrLWxV29EYisOAYjuHsdVcW8FMhKUzDQD8QVS3jCKH
1493UwVjh9czRAEZCutX4repfeQ5KNgHr4900PzAyP68+nnaxiAAxpxt4j5T/I1icIYOhcRuE4f1
hn5Nv7zfKyS1ckyvAPmfQWasnZ/3OiCFwhd0SQ/HPDhsE8rwLOuHdbC5tP3Kv+nrvLbELnWVYCGy
fUZoi/nzL1/1t5qzxcl2vROXyyTF5hBflNfxmWePbHoNMiQYDAPwMpfCx2ZO9UQIYoW3b2l6Cit+
VeZ1MobYbkPEbYF1uM4hmcvIvPMoydHO9GjBlFuIE3Rp5yMjiKWHW5auqp3Whe/V+D+RjB7iELAM
dKMI32GjZjcKEbfxbv3Gho1TF7OBw6hwdt9erVG2JI/zzQbGxnRP5YRh700Yz7gQGP7l8wmdL5U6
u5n3l/+IOH7yo5lTcXnoGG9JF/5wASMpiDegyOXPIJRgGB0n3xkr3OSzYtXzk2DyQQazaN9MTLlz
+0ARJWhVhvJSKCki3rpQAnfZqrwLYNVOIV3nkjuVfQn432J/pRtkfWVyQqWLOjfEovUVibw7IJEZ
fcPww8VkBqDDdEKwEoAwasrhk095y7LIaLkTEdsfGHgEoW7N2UZPyrCxRRNkB2UFtp5ujKRxY/+2
0KSleBYl78inAYABFpuCxRljUy/lckxqDL2km3Oz1UkQXT/G2aFcX6ZXUZxe8rU1W5BabMBVSLdx
aOMj2dC8b37EakBNIo1HFMGpynzOslfVz1eNTq0V293deRmMiqUsrCuSGVbawdZMTTxbwoP8LCYV
mPtOzHhTjQTTZenVt1L0JEtCOZssazd0FHrZObhxRbmvqMrpBNIZZ1YBXgxkmyUO2RoIs9qkj4CU
Z0nBBD95bwQbZm1lup/tPoVeU0ouaVvaFRrijOAX81XkcF6IrviJkCnCRm2MIbCWnlngj0kqDXCO
mXFEGRGyOXARJMMTnhtCfN78mScye3iZ7PYNdFpMkrl4j85MKUiKBjqoCNPeSD9dl8IKZvhoMO7Y
nLddVKqiAUlkMP+iHSAv50PAnGz0lSx+vpsBqe+ZNFsckuFPjhKYAvRwxmu40ApZy54/F6o2r7oT
Y4eRMBdFp5s13bI4s1oyoi00ljvCr3Athl1kGJU9dSHcO3gzaZI9HVC7IyjTazXEbl7q2JHuRhNt
IigozD9O/A7WXSe4DCnh7WD4qFT3IccklIlmOb9sMnlJKmzyyGkOfUW3ael81OkT2VoT4bQfbjRt
pxEtUfYeQzyaVv9cIbewFV5ek+tZeqD0RMIboOPwj5GoLvGtQ+I4cjl1p+6HhRzVvYwzDTaYvigm
BwngDcq0E63mY9Qly1hIEZlg/afwhWYODfcDCsOdAGngjzR1B9SRST4QSMV4y8LPjZXfNuERmE2r
YLFVWQMXmKkOVEPw1WAxTYpi7Sv6yhhx9uwHiyDtWPjYc9Rkf95NUgFHd2JlYR1b9Uqs4FvULcH9
ADboSUfdskt3onvBLHMnL0SIcPR6EcdwIbbTEKZc/RPplIz5jRwjXq955PPXGSWIboqG315dk9xD
/4tnBUt3rbwacGiCT93OJApu5HaFpI8XXcp2gYDlXq2O6QyRr1T4lkt8xTBYHZgHfYwYUskCgm+X
8nnNTnihVLALifrDn7pPwMZVcVvm83Y+N9Ucea3CMV0Uf98a8ogkYmQBO0WSFIDwPVGnptjRLezg
O1Z+DIchgBNiGqdFtSbd29YLM7ixm9UJiK3RHZ7/SYO5StS7Vk+zSo1tESWnyKLzAZcx/M0Fnf+U
m8BPq0SZFFinEHisC5mN9ggosxJWCW6VE4G0DfWK0HsEczisFKJPOaBtu5jqhAaaDE0Peuq1RKAg
oEvBeWfwjaIYNXBKfMZNGMA0yvcsVTYoPLzLpsydP3XCraCpq9yejJc3jfxzTlTEv+Yp29eX7cS5
cbH8WQ6aGvj+k6apo5FXGsDt9zBCi0nqzEfcoLO2BB4QhyzXjn2cSy4ROaFds3Ve6mnPLOQ16YSD
0FE32OAvX4MT7Mn2zj8fBiNyEi9Dg5KvC/uvDfnqkCAI0xAhNjvucshwRVPkqPnnWt233kzVO7pQ
E+BRv3I9seLUwkgPV0DBL+4ukjqe1AtEHLAB4Ms8lwMYdQHk2TEw8s0TJYQbTFdyd1v40Tgv2jkF
R9Pz5wj/Vr8HV6ZefmDrKYkYwegOrShKE7SEaxDDrKqJjCOXfCd3/x5jBTamlEqfZJG+EOYjS8ML
a38MZ2/nxvdk+83VsjtG0TliCTNvARPUOnM5sUWypcQC1lrQgY3vtURcRmRXAoZBbPepzh7oZ1Q+
AM6DGQN9VHdZobHbEIPtx+IHSpj+cvCD1yBeyiqyPnEVF8GAqRWuUy6IgX2KvuNxe6H7o9weUwhb
pI0uHDx4bEiecE0b7nYsYD5VrzyuMdExhXGBpNOY9BBDKD2bm2mo7+Ht6+6jFlAX5oIiKZDaht9z
gPCQLoV+MsCDgS7mPzmQvFetkPDgbQ7eeununCG08ZIKzSaAD1ICSN0CqMAfnIM9Fl976f6IYIcC
zcBuObVYGmZW52Mnj/iXMTFIrL9Iy9I+HxLrnA7759hOeWuQfJDv4R2jrwX50nYa83wyAP5UL3i1
limGQFx+co8fWlwF1SK8/6ke1d9ybzEHE3Vg1wEGfWndlCYirM7hBuSrR/dG/8K2k6adwW8c1oSw
FfBu0IgFn1d6miWr5izBubPIr3p4X1FlfhNB4OGJi2bxhqlplq/5lF6u5S4EzztdVOFjg+qPdaLG
n0eBTmphHMFQegz3QpO3P+LNQhuxxAhhxdF18cIfxkL+1/84XaDqwBXgkEbvsY9nmzRjATU2E4u6
mjk44SMueBLCkXGzXR+o39eG5nAH0UySfvTAoxF28e1kXsp0llPXUtb2X4igCKjmQYjF55YAm+G5
Jh8VdmSsB407mD9AumUs+vpk4aOzpcPOSEu8XHTttSI015cGBHMGl+eU8eMSCvWnpbUI1bnG5cm7
uygriMoLjc8ORs3EMXGZ4+8b1hUze16Y18mdCTjcStb9jSgkNAUWJhCYmUNZD5KlzSANlWJccoBu
oRY4xZV7XqDwqdMQr8OtaGOZl5gPPEptrQQ+F3543wnPTUGnGsVHYworyFZAun18JACB960yYbgK
JmV4UGcYr1vw8xdfMfPmid+JwAImdQCshA7JBT0IRWIl1y6qjFyx+xGJkNSHV28zpkt8bkb6e7xh
6x6fNRYEzceqGl9NUz2Ft/zS46Sm1Dk245TN+NUR1c8Ckucj6M2VCBSW/0ng/BTepcGza6tM6PNt
THRIs4cIBuK3BgnBF459FaAXLfJPn6PJf498VeQRr4A0Z/2Ui3Cimvj4Cp/etiEa24gTNqAdZNOU
rnI4uyshcWhwhZPJ5Gss1rKE9lckjVwfxXTIxcWOVT7hl5DlsLNYUFfZbvUh5sGhSZk0t965qxR+
UbPTnL6q5EFDMhqbUrSpp2uesbSu/6sa1fd2LWsFIOQHmIhYZ0+xJpxcB3DnB0rP7wzSgZMW+m0m
7ogem5k8W2ZbmVgaI+93F2NFyrSO1gIkHOmb8MUHl88JvpppbQtHviwLfPSuwwxWO7cAHUmBf/lS
4QoeBgH2pJIezMgBWyMomC2Rhq7LO4nD7jFx5AAI1ZgJPjm/uZ6Mc43owLV0DrQAyxGKkBLvZN2Y
TcvAtemEN6tM4kHutPGkvX6VO5btN8jES1W16e5DOLfGHZfHpazNJhIF6kdgiYS2R8fEuZ+39KN7
z15uiPAzQZRUmIq75q3ezVafw59vG+oeCGLHdxDr654f7skqB8jRC6D3/rjCcuuBBPV5ZU0XewtW
niWdN/BhZTwltKzqgCtSz+O02kBDO5rLQ8EuO6hcC84O1hCFHAsa2xU+drhtZFkCPUb2xYssp+KH
4YfoyC45fJ8gAgIUbkk5gNBAvzO3TairrJW6PvRFeekcOLKjjmeJnmJFuVLoFSH202M7nnyk5rS4
mR7a1ml8FoQ2sDq6zRjmqAWGrUjvJcvVaOArBnvEG+JT8UnYU5SboisUq4/DS8acGfZr22s+YfKv
zXFPwlqMF4sZkTyEYB+kKU+z0k1sa5XuwJGu/JNBENIDilAENCQggZkpAhlibvL9hqfkWToqfHMO
srLESYKjQ2PHaQMNiSJRxQRkgjcuI/01b4qh8byC3aVEhn2b1obFdbiyYbQDW7OQnH6m6HMrw6Cg
YIYZ/YfKC11gjr+SWh37OFv9zqfGO/aM8yMikXWRjZSr8Hrp8tRBB6V2tLdrlzVDo9E34dShdmdp
ve8xM2QdkqkBy/E7YwT2g8gdCLzumoNELr8orRXYFMyMIacmhn9P49/kxwq9SKsH4ijdSj/79pMh
xM6PzKIkjWzPW/VECvUyIb1U9joBWk/5zpuFO5tyzQO0zoL1Lmcrlb9zai/eT4uI22rf7OfYYHZD
eorm05jZghM7qHIRBds3RiHR16S+BA0+7bVVS14/kYHzWU6KHBxUkXpmKfbMBEf6vZ/g+1iI2fHA
DfZkWVE5FaivugLHKAnsX6JHB6O2LQlroW7gTUo+KdU0Ent84ruiZV9rjbhUjcOgD2I/TL5gIriu
OpH8r14zuPv9i2Ysdq0aWK+EtjkD3A4Um81MnOo91PE9hT0BygewIjxU0GauCwNoS5E3GTBU1N0A
h0mJLaxEe4dhvFuxyVFnCqWCeREqcOM6dg9M12s/YhSO21EMnobFEbNwG2mur3lwGqCoMNnDq0x8
a1NXLnymkM+xqsaMMpk5wlL5VCJy0cWCRNUxFpfeXBKxFSw1y0yxgl28/M3UtabxYyU9Gx2KiV/q
VbaNxFfWWtJsoGoLqrt51BP5ITI9tX2VHZq6V8nhkxBwuwf6YzyfpiJui5Mv8sWj7X+LxgT+61Z2
qlQyfyl8pQ4xtO2inflQB9T841KnFHplE8Ihx3y2UnWbZQP0r9ZImDw6iXvnrfp6rFC4G+2jAfXc
1qau+Yh70O1orbZ0QCPnASdF7FIvg2eRn6CmpgHp8p4hmI0mJg1pGEUc/eKEEBxafkAFo/YcJu46
iO2fkIAgfvWqjbdT9GxptOFEUUChjs+ym6StunId0WFbc3wsZ8EGXg6Yoo77TfoiExywHiBVhFBQ
f3v+sI1iMUm4T7DAYvD5FCq9fdkE1FT9ulqk0CgFpu542sKJ1NlrLxraCesF/TvEd9aPGNL/s5aL
wLuM0IDdYQXfmF1k1ZifFxVXc28xLSAubUEtViU9L1AS7jANaIVqPhmdZh140fTOTcuy/98cAbcX
hMEamd2p9gmSFIEJqNPdD3J/uiqIHlLAHThvueU8XJkrx09ovam1dJGKyEv2OcQs7E/MHcctjm+i
7Vikabhjhp8un5Te51h5OVqij3tlDEwJXTeqPyIMUVJ/Vo19o//Vcy22jkektaEaNSpl/bc931z4
1w0vBcYIlsXJwc4g1WwXcYrpVfPp/n9Bfm9Q+vizt3hgMsAr6O9+iVXmqtH6mAMakqcnPpWDZjQU
+mCMtp+T6RTQWGIsi1/tZAX0QV4cg7R5DN+H4NwvWyEi77FoB63cc4UbQ7GYVvuoBLs4fDnQo7tF
7plLFmOWaXiUY6rLcAb4THy6u1uRAY5yZNUvFYrWj2HGBE/E7FJRWB+NFraXNTDzDFT71eh+f4rF
wcmiDihEwdvQIotfZMO8NLZ91lBob+K+L+5pOnPtMk7hJkB2EJFz9Esf9UPv+KBN0cVGsjKUVE9z
3cvV+hlOVBOKtBRzAntFQvlPUjUxi0c3Ja64Eo/MbI3C7VARNCyezjQHNRWAKbDKOJQ63xuklP5M
cWzpSGjFLZ+DpvwoQHbpAOooxxj2PFvmZtPJeZ3FmxQ0vdGJSuN5VD4f0dymPXy0uJcOHG+x5Pdf
b9wH+r/S+lkqTlzGtsZpTxwJFgTbSp/aJKaIuQ/r3S1WlIy2+CFLnSS5bhfNp3gcwCzDkPjsBOwq
0eBFO8UZhkPYw3Gx2estQKxbY2/dVs5yMHyoPtaDmOor0PlHf09MVyt9hk0tsJC0r9NjGe157mVA
FmmE8AZRJUyJVOjekFrHJSCx/yKxIWOOvODPziV2xHcOqXlixmwuuh4WciqUbaDFImL3MCuf1dAa
klNmE8y41Tx7gqVVTNrSKQcvM2gos4WxFyuyy+o/Br+MqAHRjkjB8LdpFpbrOwpCVug9DONK7S+s
1+wy/VLleiFRliywwxy+UHeeFkQ+dvRbrbSnF6Z01OmelmcjzIkvvTJth+LgMM5quapmCmVSzwpk
ztZEfwDK6ZydVhXxosSrrwW5CZ4YmO6f11KKirsGTqupgsLwk+o6oSyakKiOZEvPA2+wl62EZb7c
tFYr6uoVRlWQYxylHUsVHOKRcNetLQ9d4/hWA3zHPVcc4Cqu/0d0InVd/Y1dj5OHt5PLCw6FrMeF
VXi8glM0GwyK94QqW1F45OQ+JKfc0ex1Uq8Y+AecauOCMbB+FobJaZZR924dDyUs58fuBfauAuWt
bdtCml5W8/yqmE7xHVnahvrcYsxnXvz70IzZYAJnlg7Et8UaSq+q1EXzq3BKue6RdL+gdW4+S1TM
IQ2a9BkockZxdLjlCdz6gDqyx92zF/YJXYFy/x48sMzzqfoEkGtI062HV/p7cBrdhqzrKWkP28cn
Q+sED40o4M9Y+wl/X6O7aP45y8/LLCaY86g63NEbuSVO0ri/WwgIXkEFPCjXb1dpkHtClOa7r8TW
CfL4xNOetfh/kimq/rzB7sxtG9wVrECCZYcwdesZZW/Aw7fIJjLgZKoDoG+P+0zHE85Lkv9R/Br0
tT5IYiHIwP8+KVm4ek09XXsKEaMxmYl5ziQy+AudNUUMhWkH8TrTKvk9GPDy0QPFg5c724+al3Sj
r/uDUwEpUiPXj+CGyIVGXrlly8Q5j+Vicju2FQpwXgzLTrY+1KlJi16P0rdXb4bkphLJdblAWdOY
TLuoicc+btfUEWUsovktfPKv8kA26PmPorgNXzuY3TjacEBa4Dy4QXIV5DraCNCjeGTjE0pL4cXM
QZtMLHhZfXUosPi0FVikqddu5ZB6zXj7ddEYs6mlHpeB2NzOG9J+mSYCzbBAKYTyjyBSJajrk1LX
ma6EwGMuJWgDnPOxbx8d8sy/5KQDgjm4wcoBl1iC86Dthk3WZfTwC06KWPQSl4YGXaH+wpLkBXeA
/NdjBqrx8/X99i81aaUcIuWw6dOji8vZGtK0fDy6hmV/HXFYr3PcDciGh+6UolhvQzCekr4dhxof
gKwXrhw22cw++Dz5uLofF9siwMXaiW87blHOBzWRDyXC6ZvpnATd0jgG/xQ2gSoga2IJWTf9gGq+
0b0X+JenKN7x9RheE+1iUl0PaqZ/aQcqx7x5PZhJI9nO4YuLxqy9iSrRcGEdqM+HHUEJbUMABx9a
jwFUzcPocs2OwTPDs7mFPl1Xg21ZD/Vzg9rlx2ERnndy7aouKpn+dQrN40KGOUVnhw7AzuVuaomd
AIYz4gtvGH2mcETUWJaVLnzwt2XGcVjxO6vyYiC0F0ArkpVhO2YbnU9H/6144ueF8OLk8x7jzIpU
hR7llaFbPA8TzsDbm9T9JPSqWJe6SVmJ871QY13q4iAe2EO1kKyEmJXW9udcYxBULwvyeksTL/ye
FSEQzLRBikIHqNNi2O3uPt+sL3WHeAtSkqgbsUG6CQJeYLwScWvpbDspFYmtvcC8p6AdEFvJTbqp
SjPrUxCtfSmuhaJ+jjcgaMymsOkklE9mLMBE5GLNvz/fdDb1mlTayeAP956OIy33tYT3m1TU25NQ
sXcrTBlt6oR713kjr7KE+lDKbRBetbUyHE159x26a1o+UAqKx/8hlkeCWRa2OgKT+/v6Ih4VKBm4
ATw1L0bYMkfwHq+RFqzr1LNdQ9tI5efdHz+4Ow1IICEyn/0At8Xv6AhUD5Nhnxn/bFRK+Dif3VH+
zeB3IwEpKCYLb5OWAkwC0kRFmf5064eLP7OW7clmWSOcpM43vWMnOHQy+mA3oU2PRrZl+jCoTtfZ
iaVFhuA5CswZ4KtzF92PaQ9hBY6i0T+ahhap/DQbwgm33sJTr2VDvDPLrRirKwgxLCVfUE8tukVq
A/Q+MFaDiStgDHm6eNjUxwU7mAqt0m+RYqLquZ6DUn+c/cnxnfmmyx0tc8zKvn4XEPAWbxUW7zzg
ssq9e9oVseGL4OMIcw3q6lG4sGAbueZnT9kstGw+m2AQa3YFtDoWKQhstkVTmOrp7jysmKIrIAHM
cVo0WMETtMiU4plxl73QKc1PbXZytyu+lnQA0TtFkxpJvyJ+A6xB6/X2QYKPdg5y/ItYM7f5gHmf
k5glwm8/2KutH/96lbD2evzsOKY3Mdz/LtlP3Z3uEXWnKNMNeforf3CvSWSVFJX16rFJElGmyBdj
6Dt8FmWn8XFuCwWF+iub0t33ZB/BTbPy32rxgeEt2+Ycy0stwCi7onkrW1ynRexbKj2rbC7cK+bn
y05g5VXmxA4SKggBgnAr6/6T2eaTw8awJUTZJsxOfVi/6C+aOPd4VeSMX6IKQU1JssvUpPNLI/he
m5IHwUxlW8Tis4P4/itV7y0Dbm4X4kGotAmStVY2d1yPwjhbm8EZ2AwcLeP/LftKYWYrtXOOtE19
9ULUlTANAYOEpevKNG9+UK7lyumh9RAgatxotGMQnbPif7n02OSb2i3xG/a1RrBoef/+fSp4XfZC
YJQk2GKSGgWEKCh2X3g7YfKwtnCRRGrnayGrDkIVH+0c+SezUhTfW+FwIUPJ3BXFHBZC7w8rn8rC
9gGXKFgYZsJWg9WPbHccXWF09pwM60WagyzNggYWsoI05Ngpql6ziRtYEmDVmLJC2I9TyvLCuCSr
g7JZaMhW+Vx4SaS7PVMBH0XaXX7Ts0+7WHD16WHPaC+SFqcM0VSLPwZznN1gkK644+8PvhlsfSDb
RE/pMQLy19UxBlEkhnb5s6XpfiCh/nwCmk4RQUskxm2FrmjVX1uEW6c3tiAGLvGtGMAcxs8IvMep
efKptQtolR1sy8JOH+OG7KrzRlTc3LDEYDfG1nAQM3d4COz/vsvfGNWWmEcuikjP/nDcgO9hHcOq
kI0GZR3Pkl024AiueB2Tef3P5B8wyNt5xRuVSCAtVIzey20u2EgWHDTKRsZhanrq5BAZzGHoPJy2
Nk8/IRbPrMumX8VeNXvo1ebRkCvq/47nKwAxaI2HpZwQF58qG6/X/AJrP27OhYK6J4ZnciK3W9jW
Z+LihCC9afNP7n28yeJRz3XgS7tpPo8zHryzlg+SNqKp4LSgiwZA2f0KGPmigmWMTmwFCn7Yd806
4AdFIPhJunRkyw5OiPfPB9WP7MQqOIuG3N26KcX69KWjxeV4nIkpsFH2gPMkmZKIWru3EsN12FsT
xWNlTTZKrLTrtdZhyCkf3V1Jc4lG7Pqhy3vnvo2kCsbdX7qFK6ba+tFUDAWSRaNG03kPPQd0y2kB
at7b5jAiUUUF5COzy99FFEfu13rJwmXjU7ZT7eAR3naZSynEkLpJ21Thrjj/m70SNGrDJqTk6p82
Ch78E9kkTcB5qF56/lKyYfAJTwDUnSS+oC+8RLNAi67qpJLENMAUGbxRluLWnsXfD/OvZiJDN7A9
PD9jXuEuSJXIzqxhF0tpayCse+4640LbZcdE9iugaKfWIVjM6Lf4x1ne+c3qSuy699Un/KAVpEaL
GCq+363OZ/FT8Z+bwRZCCWrXkSzM1dIcxDAhfQr/Clqm/CQjkl9lFEXVGqvjplj366cs5cCG+BuJ
Zvnet4gq8rFxLEoDFLzZ5pZAS8vV0MyR8Ei9K86UNmw7oTBNqLHFWMq5iDqA+suoN6syW9jJ5G4N
Fcc78oofD15w4dOjBG3b+BETK62++OD2Ux733iocihu/eyLoete9B/234bnj4v8/QScdzXMr34Il
pTciY1elYYdCNKB2qB5viETK6v52xWEbKF+Ph7yC6+5wKx4PjdrM6/I6RtZ8tIYw8kFkMTwi2e6w
syKAnHSGt11cxgOG1Rj3TLjBzh5BdrfHmeDR2HKajCtwMwbNAB8UPqphZP6D2s81sbjFqbjza8LT
9SwXk2oEYypwW4i4Z2ikEaNiw4SlU6Ygom0qf3qJJmOd7WslQEf9fvuUjRPH6vXZLBka/7N3qCf/
vdLEF5cSFus4as0iXo1z7p5d8QZOPL9wX2kClBDvt9oRcMRBi02i4AmPc/oXY0gM2yezVUTinwCj
K6x6hxp/OTLb1XDjuvndtBwwscbkQ1ScOg8MZuMaRKkHji6RJK8KxNuzBNnDnysxgZQTgk3t6yaV
WeQ1Vbk28sKW+LniqVMGqzTJPdfXMAkm0mIhX57PqUA/FUfxsU190wK4XAqMtRLmpomNlDoWQnUk
ECOULyFAmy4R07IzCbF43DBn6HLeaFh2PRVnI7WXTSmnG0zoRCRmqwpQsVvVGi6Xiqf+ZBikmBa6
g+T1B1Gv5dwBhCsOq/IyO+L1sfAZCBvu3hm/T0zl0njztETmmdqJpinf1wTlnoUEnT0UUwq7FRt5
V/R18p0PIcnYqIrGknk87coHKaST8t+Jo/Kj5VmziSDyPbn190mJO9lyGNSluxZWKXzZMM8QzSH8
SFyKLXORow+g05Y+plLJgsoGrBFrccdqDEhBV8vD020nM6ZgZ3snDucqjeO4S0E/vSOWLzZn4NVP
D9wR/qzUwo08e+oqcjvJ1of+Qzf7QuSpd18wVw5VJU7wdUM/W7U3XX9f7FwQA9yeKqW1FHQPNA12
q+6g/a5RE1RaONlKunxW8yNaXPI6+CnGcO4DTSwO0E/u2uZXBg4MRkkLJA/HxhPy30bMNcWFe/yc
MalqSEAAOhNtCbPsNdZRVUzKAhfy5YsPL4a6X8HL/XpBVAlkYdZga9To0MDhvbCxccg1SMrEf6mp
tuZlHgk6BG5c9qwSVDUgFT05PJLnbyOoJkX0uD1dB3toupCLAdTq2KfVOKfOogsJPPlRIsurfWqA
nf7zrERB/Kd/PJg86P60FkJphdbBUcO8CLkTU4JPqYJAE+excvSUlZzcpCok4V+4EXtPu08bqgAZ
5ryz/nOmwSa3ZmyEGetYZrLP8FP760w0sx16H8rF3se09rBtL+ny97stYbSnnyrreS56TNbdhhdm
Rs0xnTy5XBHPoHom4DrvL62XsD6VzmzEwDEv4lphw3mXSjSV10nveSKwTCZDiIFf7OyAFzYiCvaw
xDjjI1n0NgVqqIxT5ouAR3WHfooEl7HxwDyAZWN8Tt4agCDFeCgsDFU0RUf4x2HwnfhAKflLsJ5t
oi+DQdmV0E43lGmAQZjC6QGxCR/DNSAu3+GCqQQKKrwgyd772SYV7GKrpz644y1MFo6st0brW3hz
MGiI6UTg37YYazbsq5b5KFWRD4q62k+MBW9nNzTMfRkfuUyi8qzjFZGFGLfWVSR5/6nL2Nrj0fzq
UB6g7syiKMWvoPmqq7JOZGWOkJQOY6vxd6z1DJD52kkWeW1IAFPONVwX34MkpIbvMjTPOx51T2Mw
fea9+sgW9dRlSrbBGHFn6wV4KfzxZ50Bzc+/+yLtYX6fglvPioQLLqcyrIakw1b6LG/0Xju3Q4r+
6OqLH60yzPcQFw3qZ3sqUfTLfHdCJyzBzLp5SIuH3CRlH+Oc+ZXVrKa5nTmxhJrJ3aLuMSDhOWvG
P6oYgG7MbNUBA8Yq1wi0UURG+Iut0vsp2qdwjhltMJWMuvFBne+3h97DjFF42c40/tJgIopPS0zq
CemVr/HSUar9V4jj+u3hV4hFDQZfty0tastzkETStun1DVmQhu7hnc15d8PQnrqNpAZSd1rU2dyv
fHeXuwtjPs62vPsUgjBSc+Es+xTOPPilXrt5vVJKQOKayaw/Msc/5X9XURaWphT2AIqsK5+O4ZST
yjVWodnerTctYOZ0Ha+otRZ6uWGmtv9n7ZgcOLdF64fR9mot3yH3LZ5rkQt2yKyfi2Tw/uITnnoO
ZzhRvuYEMwm4vP4DXqUCNdLh5JAhBEZNgFf2/t2wft7psUdWa5PFy85JdXP8L3Bh8KqpXul07MzQ
csDmVWmF2XyeVh5khqFI/Tn8QaBTO3YxufAgEjh5s2u+w9Dme2oVqN06dRwN5iGBX0+NNrHjw4yg
5YhbS3y+MijXBCoHjoAdZ98dkoq7ETSAYS5/TywWQ6CWnd8+riXPcUUtByJ81QDfLkHQuqXCmpJa
nsHvlc/dfIwa87hc6jML3lU+awOhopTircXSDgjJ3XFgeNn9HO0q1CRO8pXlzJSr6uoBZCqlxz/I
2ZdZ/y4WAigutPm0cNxdIar8SBEj6tWGc6q3DbdThVPMGKg0cAlrz3esAy6H8uyvYy7zADREke3f
mg5/3OLI49P+lV7CCZB5J6AP0BEJqTcSlyyZ06aSmX4mBHe2U4DIajVVQRgKPJ2YCa5JqRAVSRn0
cAzy8qu6K+oVwlTmiVaSenlSwCicOPSOyaLM8vuSXvKdp0gyc+5x3WszLGTfbYQiulJha3D7JUe3
TP7MEVtPTtWuqwstwugbxvCq20+NGaDXU7APxoMi+KTQ16FkNU+uq7Thz9IO96n87mY8ZLcHhz+d
gkYj98mHsE32Il9kD6U0QS5W9VE2jfCDjLNIPDmdQb+SSp0snojFOfAl++8cpVZ0290P6L7I4gcb
bhh/wH4Vy7i5jReWbcN0gbSlKDXilKrqAli/hnsAM5LChIfW6mtUgWvj+YQpNT7voo8OLR8uWrB5
mN+/GFGLEqI4l0+CdqDEbszGs0pyP+iyJ4wTzWm66Lmgm/YnVtUzQ/+vkr7LvZ9udGKj/8fCeLmU
5+YbEZKrsUsIoYOp1GGQasPCWDEjc4U/BEVo3xjT8eMb7KdCg2yiWWMHrULEx/G9osAefXnp+omc
LGe58zMWyLAgApqjwVgSAuQ3/8zvQlzhqpcseHmY4PdbSeEHqWXIRnq2Hkihk/RemSTOSZQt70zx
C0ocjr6TPAmfcdA19Du3YF/JR03/XT+xjOwcZLqet5IDvyiZs8l0s+TFSaj2UmdkTG8JemS3LnGM
iFZkqZUqbuMaru2Wn45C69a6b/iXiKdJttahFDtfhTBAiNhwaIXwWqv8lkL+0SkeYpv3Qz4+oduJ
9LQfTKZXWhOGhx6LYgqCOahW63p9Ij9mgnETeqkQcp7gdD6FBeVPiZYpkP46Ba47wDSbV4DAGIwC
LG1S4QU7qmdU/Pjnd0YMhKwAOw63hQ6kfXFMH1eJTFU19V4jw1TtjjGGhemqaHKDikn1KKQcO3nR
V0xQ/bXJZvWnEAevnP5xXlhdRXKmacSZoVs59HyGkqGsp0J0JXwQlcIjUAfcc3gCZvJJb7U8Qu39
/f4cnMynzgS1R1LGndi5u2NZsiEpmMJ8uDVgDESiL8m4Tsj1vp8gDwBijueqoJb+dc7ut5bEc02p
2xw/yK8z0kUe6yD/NQIvUD/s6+f1Kz6gDiVnocqliQ/oDFz/EIH0HYgLSqRyQtcAT+qHQlz2dvSB
eG0TmaZxG589waymqDnrnkWBDF7u/hpxxj1hP8tEhr0Xv6oYa54gGzv7O4YI0jO6mq+zr7s3hOoC
SD4AfEoYa/Mq9SD9Ujo/FBMljr6PvWAkz4rIHG/C41lSS5T2LEeDLNKXobFbuZbZQeruhpwtsHNk
db2C2omgoDl4FpCWfjZ2Df3iVn6tJKGEwn8+eUfEr159gyqpqpTKHS/Qxge3nxt/xL3+o+OKuMjx
eFY7ZoyUpXDjSUAh6DpUn/vVMVRp32PPBSeHTnoFXNDCXVQwSW9BYx+Afxvqf+Y7LK3+RqRoPEmD
zs4ET0sUtj2ztO9FxY0Q7FXLFWHi7To3LhM+EZdieZ5LsuVkYq/R5Dw9J9/RhzZz5agTeJsSlhw9
9MtqZ5XsFmLgT8sfEaBO0eg58VVG1tisxDJyMz/iq5FYyQvHnUWVmYyo9r8APtLyGb4xhEbzDDT8
x4BCOcwA+MSHLahMRJVyn7fBklWR52/GSHgzLRAV+ZB7cqWkA2MvcbD0Q1ACQ0VaLokiwpRPaO70
dtKyfmwHL5SFOTMGPYJ7uj25qclOZvwr5oDHbvl2j6nC+dkhi/fgOLMDANrj1AFoUqe/qRwuTIgK
QTJvcA/vVeeE/GqZW6LEL6QRVzQqGI98Rb+jL2tFswTjQoBsRZVOqNmStPm2W3me6O8XVqltB5Gj
EtEHlAjI4/JWyYuRqopHmDgcEYbiFfMQ5ILh+lcMC47hrCiPOluVlNc1zcVUV1ciCxRC7CA8fmOz
0zeWkNVHBGGyriKBx+1QSzUw4ia+ypzd1XMdLUHscfvDKyO+hNkC4+UsQI6Fk1osdXnWmsvYSM0O
e12zy65bMECj82hCgcRIgbpRDv8jXvJZroI2kjMrZoLqJwqhb8aHXMrkfY5DCtQ/ZKjk+rrBO7j9
3np345Qwjt58ikO1oiVkzPcc6/sSMu24qNABQ+9GM6vatb6prHSko9TDl5r7rMsJqKAt2mtXtSmx
/ebwlj5gGGsuuVxCM6q8Ilk4+ilLSprcKkj8FRp5XkIOPm2PR9+7iw+6nm/yW8Cn+zzBoxMXUwrP
LH9RI/dSYXNbufEEViO6NlWQ5yk/wY6fHkgtIQ2GOSBBB0pofmpqjftOlzcNyR6NpYhY5WKzOlEc
Wy4aDMH2fuCUV/QP0YZ/WVd6KCy9/H+F+1MYVI50YBs9VDWMAm21WINzTiHN3ihhBYavWJvbRMSI
OT3EsNYOE6lfGUX+nPqW6sGf3KzkHAY5xOFsE0UmufWG/WcSOoovqLAeMTI5E0oenuRTPyOO/+dW
LZdisoJy7T6B1DZmh3qcKLkgp4PXAA2IuQR9GM6e0s3oY/U7/eBIq4D11qsKUh3E/a1fjNqZCu01
WMGmeFD1WyBkEMEFsJu3Bct51wvdcJWG9aPps668Czs++yNbm9+EkY9mmcZx90+vLZIbHvMHMofW
OQbbDOmHCHEkM489uTV28Dw4sUSw97ESMMGkDJnyN142BE92+UVzoKkHbULFN+3vSd7D4isiiN/v
vuyPtsZ4wbotSBzLiOclKZ+yPvZzEXX2VBMTxp1P7mSogXn5sLvaVJi0CYlXvpXb3/95+435eEou
cbA1EUMdH24TnLTh0qKSyKnGcetf08Uamk+kx4QnI27wGHJP2MbaYIwKp4CvZB/kcUUtHJpyvlxB
BSOSjCKGWsZ/vW3OPSkkl/bO4zirVX99ALvF2QRaYg3ezqpAEz24T9gv7O4IP2189Wq2OJUVWy9c
HUjw5rxmodEB1qcCJasChilD9Hus9tghdNBCIQnQ2k2u8X2lBzT48VbU03k8Q++rGw9DHa1s8fht
YfeeTA3KSyRe1lwICf6YOKz/uEhMSrKP7NuUtAqXxmxplgp16nKzhhYsu33uEvd7muSdOj8u2MfI
A0G4JlPPY2WUiu7Y/tkGDeoHppMfm1QD6H1zc7u7iqQRtnz2nymPcXX1lWWwWr7a8KTBlA86lhpD
FtiBsnD3GSK1S3tFSOQwiQgQ2VK4i66vDOj6ZmZ+ZuF1wRvyFfKISciCj8I7Xuetf1Xdc3kQNETz
cODNQ5OQPd+RXYJDLHo1UZBrOIBHtDddopXmA++JJkkJg2buyMPaDPVx3L9REo5wI0smaJg7s5bl
8kVsZctcJHLFj+Rz2q+LWemt21yHk4P1KBV7OgQmFxtPpfYr313J0eJaUOSY/QDbAA7qoBol36Jb
TFko9YHEidienaItSjtqMjTORz+Py67PFhV+NlE3Q3fjekPb3OzQacebnghfoBkmTPU0vF6TqMcS
KRL5W2t0Ehh2zYrzaLGkf0MFg/UTtxsHOo1T9z8Pwq4FY9phgzMiUZj/g2OOEZBKgBDssy6/unoQ
ZwCEsLX79IwUdZx/wuG9QFMPDaZWcljzocVIWD3MemZsJuJ/5dqf0EuAP+1778ZqPcZgbb+iFNXa
uiY+89A8jZJyaiOgv3UjZcn3LlW/vk3YzTFQH5py8AMcMifdBebzpXN53uuy8jZojia4UlTpQy9D
dOCRFbrqfVviXjSoZtPTE9fBBJfMB6muhqgZ+Jtsf9kcuC2bj6BAmCQIKW9GAOtK8ZhSdZmY5uTf
fZvlUAOzlLpEhryvsTsUmOjOb0dlFs2DWOi9Mg9w9H1dii8kEs9QTBuV1NJ6kQDUEiMECCc+NKLB
oi30d3UW6kam/+8pnXO62L6KK508WIdBkw4kUtMg0Ndo8U/gFczN5u4Xc7VsgbI/KNz2NBGOJhuv
1hbkrt2Ym+y3xx66X0QkqLPAQZ+Obnz79OOCdWJg+fm8ZQXBz/lhCFhC4CusxXTOUn8H6o+qEBm/
VenawkMWiSW3FfEwWBQJoyIgZGpDLZOQcQLMUXqev6wx+QtA76JD62WRaFpwHN51GARvwnckOc5o
EfzWvc6ZprFfixvDiSoaUREUHyxL2XtHUCZY2l2stn8B8SHWhUsDskqywCfRpZCGhutcxoEapyru
igcI8cR4Rs11VvS2dCAd3/0vCbm/vyQtJ9DgGZFW5k1BkEn+ElEmflnkJJLHMfeFj/EyTvp6rR7+
qQfOP5N/3iJJ5olj7DtjVK4mnVkTRaFUHfkWVF9YzQgduN+hfgKPdDZUOm1WYkKG88O4VI7Zigli
CO5Yo4s/szcJhJpVoPIr9JHqw+jJjlYiPClMg+aUhmy4j2Ar/KS34Cmu52anfasZP9AMifqTdiip
kGRyM68zbj/M2iilP2GFW7v3KJKRk02Mfagfl0N1FKfvIpWhqXeGyvAJN5S6nDhtT52ZojXt9tT2
seIoutJtdMdJrCVUejx83aUhtITFhPcm8chGgNfsAvT/uE2D8GPan58Z58R9UZmTny266Qv3eq6w
VJAOBeFcneN1taXRGHR5eE9gZuhHY3/+R9paRD+gychorTMpqC+AwF0PksRp+YMAUmuezzStl7DX
zviErOYJu8Sk2ti46S3F6YlqFvGkxGfiTm99O13YLomoAcFC0fN6kXOES4fn5kP1erEwrNStJ2y6
V+oJp1HOgZTrjQ8deV2RzYlJs0quhwS/OmOD4ViUILhGm6DtQqxhD58g0OOn87B1A9/VTUTPwXgu
mBRngHWLBiD1aRCv7wSwbu0SWaFM1Z5kfleWBQNSUEbl/TwdSEv6dB9hnzKBhyKnUlsJJHJ72tfg
uZ5IQD0JxGUcAUC40Vzb9ReQeoHLjeyXZJTIBZaJBGIjGp+0bZExI02THh1YSTgROQ1/8SuAA3/u
u2vURLk6MYpGV8cDoQbA7eXK5UVing8x/wGigSqBih5Ipi+E7/O2SRWltD3kbu+PLJM9nJBxVcRp
LMJNeV9UXUFs2Bfwi0a1DbPzywMF4XhIuKCQhQKo1KVqIib3p5oN0HjBT9ivEfVA0lmXmBxaljO2
JdJ69XN9tGp8KwFJOQZ02Z3UdsoNspVb0XKV5FLN6FBz5my3TadwMeugEI7yJNNlc8XK5s2A+1NJ
+kUBvHnKXNpwK9mhdbUJkUCvJq07jq6+R/ksLVbq1NRLCv1xtSSWmbqVpCu6pYcmoqdG+M3N+kxl
d6exYewKwVYL6UuzO/txJLsai7WxdZgwnj1f2V/lkml96nwfwcpIlTZQ32eeDPDnzKAwdhhHe86K
xqp6tQ/zFTZsBQnMj9Z2r8eV2l+WZLMyhHHXLD6BOstZxvGMgBjf5uZ/Ecs36v+aOmQeIyIt1be0
JHNRy1d7H2nIlUPuB2KPzxFi/uSlGYsTFeVOxQdwqGA44ij/8Ia7sHPPfpUqb2NH1saX7FI9BK13
DOc1eImq6AG4JyB25/T2cx73Gl1OB1/mj65xCpFmxoXKsEdGEj332nCPbKZS/4OtAQBgbbGC4ZeT
tLg8zDchuAlS4KVc38P7cAzxe65hfSm3eTPQ9HZ3chllCLAJ/HB8dNLymy0mLkyfot+fTGC/1Uip
uG/MZNZFkU1wlvdwxFCLBKv61VPEQPPC3gbIyo4qh3UD7LfwlImAl1CK8F7DxZdFu2l2MjLJd//n
2WFzs3VAXv4NjEmN3oNLE3uom1AyvryDEMoTg09K76tJ1HQ3H0PPrXpvmeLTrRuGHBkUqdzLSxew
N2qrl1d8xzVa2FsFr2JOhbwe2nkQYrkf0jnintkTryesy68UKrKzSD5aLrJI0I7Vroc5Hgshrhv9
w9cNLy0BnkTKzKuX43PzCtliZecOYxk+a7zx27tZoUfNdM5MyBZLPyxBtPazRmTtYgTccPZoMPf9
r6luAIH2kDqRPylZ18+MBTGnsuS1G7UA/aoXpkK0XNGkkIrzsd6OKf2xeQ+4hTMf33V0YOQVv980
4j0nBmmx8DuWU+PNW4x1swNNwkJt4yJUvxQegaKLiCi8HswBdF1lTEIabsWrV2chGHIjXEzcCE8b
H+DpvBHaIB9pfcQNoAZaO8xh+V9FYyS9AuHMVQQQY8KJnu6wCkbtCZe7Q7W/0tsp0bDly158Du/A
6BNW61k6oHVyL5W/ZVs+nzWEMV8/UEvRWXO44+hiXm8Rg5+/SzJdBpFUOGg9pV5ax+hkGHZF/LLa
iHlUgzeVhei7cLIQYYkDCxDThFKRbc66bUwAYkj7XAH3QdRmkFEfiCKHmI/eJ46FTsg9nS8rxew5
HI6KrARCIZ5HJ0hko0w9qnd8zfqEB4bWfrSOv5E0s+3EeImOSeymFjxN9ZliA5BJ2ifm6F07q5Ba
PSIZTff7v5umgjQE3J0d7Mk7YdQaNOPZoHZPfQbdDE//f8wkUt7kqtXutz0EFx9fq9Nx/uKx4du+
YhFesduL9HAkIxr8Wpu+p6OiDyuI8sJZQFXxHbWPnZ0eYGqwOlOGNpG7JVhaYNfImHKld5PsufGT
Nm6yIoNp1u4lxPCqhzmHHM4UBCW7/kJsE+ycZlzzyT8PNfNbCcNhDVGlU/kRLBmePA04eIKzftgw
/TbVijfqPc3uaYThAcoMt4uO1bT5S0Pb8YNpv9L/dtmN5pcvRmmNF5RFMmgZqHkZUsBdMqeCdYdG
h6PKmOAGB4Di+nQsy48KWdtR7Evhiq2LPQkgxo7vsW99z5Eawe4YuHRAdwcHsv5ai9bv7sAvyMiG
RgYA7nIGHs8YrSRSLCwpcJdNfVoYd/FYqYudpPHQUW2M/DfQsPROLcReIAOW3XVfh9Np5LbdRd8F
FEvWuMlU+0IZJuz/SeOngknopLOJOuZS9njDXVlYM+cpqbxvIFSj0dcfmzsvvZ2tn4G2gXL52edE
kIUg+FU1GwYlArEc1aDV8SQzjBMiaiEuT6RRUpulOWqtBkNfz3RqO1IM+EfIs5YodU35WCwhCqSR
mMc+ktr729XU6nU0PgDFh7DeI2rtGw8ZHayXR2VC/zyyzidMsrhnP1tS0Hbp9J/wXvbA1ILVefw6
UhhX3AvmYX89lR3fhXIuVqWCk+yYe4ZlO3yTzmkX7ftsnBxn89NGwBzpEdLy9jaxxo8wzRSCUpuA
dHGA66x1Mq0pTZx75ydNcs0Z84MQA2WMPK9xUB4hF3TsR7UYPvRDAa1UsLgdE0K0+ULVCT2JXcM0
TS92Euq4z29ueXwuseJXjDJr7TWnLSzoIkQYIZps5lPK1U7mXzSdY18yrKaZS1pCE0qQqGpTJncv
dsUKcNoc6voQYMe6pAUzulurRUkxRdmUMe7Qerzcpmx2D7f+71QEk2C+AWX6qmFLTwEifXpvTN8D
iWOkwH+rku/FSYJHAp704L0E00v7I05I9XvG1CaJsr0YkX50F9OEYSZYlL7yWf97YHU5MoUF/rT9
HDqVT4/jyd/6oLU8UFibweazVfqqQrvMYWtw4EmM981RwBSMbd3/ueRHqzW7mMJi/pbNNd6AdYU4
PnAcz+6exkJjmku6sNSgQJvQxjsuzu2ziIL3qsG5LiaK7vEsALccJZHX/1nstsZWue/sNCE2q/Q/
fz/X7pXyxwAFIaCWJ4P9tCv8V1FJgS5B87pe6uDCQwElRTbxjG2I5gHHqllR9UqRi7t8kX+G17f+
0TFIzhsPH6rRpplpQIz00cGxCCQMFpxQGXjYhFcx6qF71TW3mQ7RTtlQxwekvbdDgt2WqZYTL6wm
vN/QrBEy30PQuu1ZaOvTsrrtT55C5kBQ1ZVqFPACWUx+toL7ucQdUN7gmRzI43GAWoic4jyCbwKO
13lMLwdMoZwUcAE7pT5U6y8YWBLLOASLCtsp+znbb+5lwbH3SDUfM80Drgc5cshdde1IBTGLuoY/
K+rczc9oTy1pehXokTMoS/oPojIeG7T7+a+9uSDV4c2iLV8zuM3C725V+bn8H3VSARIs5KHH6Pzn
wbSiz5GEc3tMQl89OvMEjYr6Q3BDtnaX5RVRRC1WWmjsPrlCiQ0gJeCvFA6XFyJSTRZGEANKQCZE
Fjo/mqICHL794qgVcCL0UqMCNgDvDSF2Dp2UIm4wSrWiPpEb18EQH95yDq2u0eb+pg4JMXCAwr7m
ProWjcsCMxNCW+0YRORYJh2Otspllre3l0OGZRbO+ht2vL+6QUXJ6vmTtdsdRizqq9sY8JsUDBDB
PDf84jqhXoHOlIBsOcDp5uQZJwTnuyZWr0F4WrCeuhwtFQl02DxtceHTtIKOAWFmb1uZiL/IZBFe
+f8u0/G3eaQi/o80Zmi7yBX2Bi5/N/D2q6JXUNIkxMKMNZSiZqlgXSUvryzwOv3EjrrmRrotlOUT
2oSCG+kKmEMTzfljVQNKdX2BRwZGVNWcljVwFjbknHfALEcaCl4X9xZSrTpHBgBh01504raYGH+2
7Ex3AnXIbLaMK06h9SIlDaAZjHSg+o6x25YdZOX2+oHjmneg3Y1qvuqnV2345VLH2AmHl7X1thg9
b4Mx1om8x2jhUFZ5/MsITkXTJ4hvFC2z5cEVCcmZqOr2wpZnWFqlHURNSqWn84OZBIuqs9e4Y5HM
5Y52VvXyb3TuGJXlK2ozVAVQwQCpq4dBnRApucgtKkF3xnZllKcMJ7aDadPS+RIRzQKu3njcPADj
3E4iIsB+7iwu6CAGdWDIMZe8fsz8LfZ+0OQIve+F2XuQ65/qJubrtFZd2coPpOWAV+bVMWPSqHVh
VKuzR6DfSoP8YmMNWiWsNHqfKaIgM8iRrFZcaRFcJEduc9wltv308x5hvVVN4u7RYOM4p2KiNPGT
lymZ9Zi3H4shAn/NHuIblXU3eqVULqM2zdLYLSZZJfCzOmxmay10QWG9nuJTE9x5ZkxDs6kxmNzk
uPFHIk8YdESMHDvBxusoK73s24Bqggk+BtCJHeHoMhQZRMMI0lhdGY0Xj0vvtw0fVkojahODUTLZ
538kP/bWH+n/asieuvX50ehasOGzRUtXHcWfc0Oghexkp1gmUYdV4tvjvnMUsRTXvJhlQpCt7Ris
yAov1JYVRdbWPG9mtgFIWU7B9NKG6o+VI8RIr/6QX1GZyPmwZ2L7ke9BK6HQvgfTK4v4rc3uvlfQ
WpPWN/LvMqIdAlYEYFYXQxfxPd3GU6RDTF5YolmJqmYUNgz4kWlykZ1sMcAlxLTKdDLTlHFpx9hY
18c92uFi4TGzjCakVl0VJ1NJO9FUCmQoe3veO0F/r6ph0WP7Ko6vtADlHDs8wbirPEka3tTtTuFX
y7MpQ/Js1DieNK+GTciP0Vq4rAk0k9x8fYz+Jwps35gkE5zx/D/Sloh+1w6CKdkvCJsGP2UPWKfw
ipSOpCtgpdGPxG6nQMtl7liajvqHSjVaxGIcqDnnn8gxh9Tr7QZ1wgF7FTMqNXhlWNMi2cSHVbWZ
Y7wBNckRODqBh3sPqov3m/JQjNLYWf6xEdkm8FK24GwM3jPg7XRPMusEuUjpyVSpRp6OY3GEwhdC
Z3S90nm68uJzERZxSSqrhSQpNAhXwVV4OU66xEorWNE39H+yqhymAZHotrMv9WFQCih4nH9q4ns6
Zt3um/ZEKUVZ5KxlegoScfQ6dESai/mBNi4rXRkDTFH1lYJ16/aJcbso8m8xV8k+//BossYzT3Aw
VoyE5qj2woFiv9JjDLTZYXKeJNtX7ZTZltGuhD9YrIpqQTzvszeBSOR2ZAoikb97nt00dmLss048
eT2+j8bz4bHvlSe0uyASOkq7+NIH+cuBfEPtbjfziOJF9MPJxwQ6GQhhLSeVEVfu9cHHBmv5YNaV
oqumbV5L07Oe2iOY8tm1CZXnA6Jynx9Tgj1ljLyfpmoOg8zH+yZa/N47d0/Xdv2tKtuVTcP4yxQz
/OkbGkFPEG64kpo/IiNKifVBiDqdYS2YPpuqW/T/ajgmakSYiyROyaD4Cu3UogvRq1cFeYCnCIQw
MVqZWFQcW1J4M6OlCDrSIiqcUlRVl1LD+i5lfXA1t7oVPlWS0eJN5AL46R4bPuQ6B9NrPXfUMY8v
JNjegkXZQ22dXUxUh3HkZhY55QgCFKp11Uqzjz0Z3NC2i87TuAxiXLL5LvJCSrp7ihEmTLucRgsQ
59mJVMGhCOneMSbK5sS+mAdG3pEwf/UIpnSXvLQGoSg6jXanNYE5tRll+EGCNoKuaCApruDweqYw
HBs4xkkLn/5nfMzIhidmbaMjeLybkipUhsC/5m0+ehuiuccDs895VVHYhSi3fkI2TahCW/DeEN8g
unakHDR4I4NLlb2KCSFyRqSvCRugyBB14PvKmb+e7a4ssgH2/hgjnWDC4Kswlb3JrCxU6bxwyvME
TcCis/RqYu3wZhskeayUnM1utvwzV6HKgpMR5btmoj/ntB+5l0scBCNTi69C8+eZLldfMFOzLop2
NUT5Wq9gS+Mwjgsbf8LgxRRsmioHNVn7n1Nu7R9BdnNcBlNr+a2nBCydeQ/QCCCot1R2gqtaff0J
F582x6Vo9bw5KMx3TvStoYxS4RhCCzegls0SedmchGaNQelIACuWd4Ijzfnsovpv/ZI5x3i9bYGE
eVpz5b1qps8+N8Eq5U9t87I+ZWbpzLhxTGwWW2FZYuGfRWHzyBfV+McmzAYqw9cuZtCmWA6WrGeL
Ihiv9WuqZNv4pl2aHxjGtFPZxQo4y5UB3PCnndrrdrTee5+/aztyHQeoPm8ueTZC2Sr7adDas9mA
qb0Y7bfxFqC3KXWbdlo2jnd9Edghk/OzG/sch2yXrmIzuyRtPdw3VwmxrNuFcRsQDcemRPxkHWtu
5WYHqDcTDxaxNxJXQFJN83HxvXqBI8HDanc+QLNyrwYbUCTNN6yMdH8X/N8aRAvXAzC/kIodW/lZ
1V8+Bg3En4hdoHpnYjV/NOG6oF+eNFxxu95Et9BAh3mTw3tWlpC/7lmOAnCNTw4f13RUzXFLidHT
BIdnvHrddXQpvDFzQfd2V96g/qi2qy0Z+0+ESFGrijlRMXhMTQ2Ot1Rs0zBMUbAGWgMBuJ42EaIk
CdQO8WNQZ3pY46CCRHDYyewhLBYbTwt820dQeIKcYXdI2CKSTbBC5aInHhhos5hTKBV8/2FaiXeC
b9yws0s8p1mFbG1HEfQde3cqRFY//9Ht8oH6q4K2CujmqsV+ugXG5oQE+/JYwx3auWm8EXdsacik
oVoSGwf2FLlgfPLzs/1wed+080Oc5zKtGxgzNOeEFeboNORiK/40S6M/SKTffZ5NZi0z/NIdHegu
ON+nRWUjuPJwYSxXbl1lx1e3c06wURIVj4a32yDhrXOFIp6DoV4wQshzpqsDCXH4wtAt9NkkTUXc
e7zoQKAztNaHUAplqG1d7KyejGtWqNEqxPc3xgjmZsnl56qRI6o5Bd13Er/SFQmsMQaA6LhlOCuq
PhsS7qeW2X4L4EeyjutUC46PiGqeXa70colQUlRs50VeEJNukoa/QFS95zbBVxC5LA8EgBFKM0+G
oERlq6Cwf4GhYdSw9lBYtxtodAGIP1wJPHh8sP2M868tDn+XUsRM7FYcB/y8CW0Gf7anT4ZSHAZz
V1jduT5tMn1358Ralye/zU9EIsJ9tkvOXOuuyj24FHWnhsXrsDt6EAo62gqr+2rD5RLfYBF9pBda
ZUVeZVwKI/+nZhyMlWwcDwdB8YfMJ6l4kUWmX32eba37ly6kzFioS9kFKGniNkKl0soq1P9NRu/S
Lthix+bu1MZesI0dRwFe0r8QxWbvB3fWFGF8kZhQO/iNkN0rjBxRFTFNJFp+eT4PaOqTZp/ZqY9f
cPuC6jZDYBjiwEn337Mnr13zvDs+fFNEPAqakv9iNLcCHFrzyn2Ht7EoT1RMq0+wPXVwfFJPpVVR
EwO93Xgbv25MmvT/nn1Y3mMkU4tFx5OnVcJOZJD+gP7yTIh85etlkJyIoBPdsmgFvqm9U2AaU3yA
Eb0hEYjIo9iZhPkQIuFXT8CFCMTXLrXByLloCrvdSCGA9odST40Qq/QYlpYCyiZviaXYkkbkYkK/
5WOFN/cj2DUpzmzHlkpiGbk6y2QgSuuNllWlEeWFIL/Mt76HTfuQo63Ix6YJYWRpB4Y/4A+CzREM
NfVe3+x8dk/AFrdSRDrPq9zuLV2wc5S8X9KeDImiJza0dhfBZ1bLohkKjz9XXNvye0kvGvC5H9sN
zIx4jK3fKGTXApIw0e0p3dv1ERcG4afKIIr+5vYk1stxJy1UTwdhWo2iQ0QRy5x/kQmdKv+I8Bq7
Hbsw6pkumEk/rPhtuduOFPCbBN3TKrPRKKeQc8ZR/xrdrvdRzL+KdJ0Wvo5djIRn8oUzIq0EtFbS
b0v3jnuo5KDCmwVJKigBNMGbsPur+HqNG8+Gg3wdwZy0w1KfUttd98iTDRNIAonBGOqb3U8RJe5E
qAxueDfutv/LmiyTA9v0gF24I04kz5ChSdVNnyG1ewmp4NRTGBpKDWNKjfVXhkHZ/j+OugVUzK2y
8PxQGh8YiOLXPJfqViK+uzpalUtGjsZl79CKMBva1Slwwt4Iq6AV/5n6xTGw+TQujMHOFw9BPMbI
uhHeUzFptrgSfb/fBu9mAz32cKN4vrbPeppBjpxWaL9CrBPNjtZyu+pehWFgxmv7OipqUb/PGgLy
po++azONAcVQpVeH0ajiYAjfxpayZqkGHUIfzoQB+GuwqW65sRCXvWHNjBicdBxaEMXUHi3LXIgh
Z2WxTEaxMcnCOqMJff3k//rhoExzPDx207PyLfRaKiBm9Nv895U0hRe9W+PFEe5BWeVHgTmWv+tF
HmRm2I+T9hpKlDu757ikOA1FtwvTmIXpEUGySJg0ze+LaLF2gxnx5gIQuFGQAi+hUiAAg3+b0qWo
h6Dv65dn+pr6Ne90OlXR7JuIzrPxRfdBsEU9BfKi/70LjjWx4tCi5lswwIgfJtjpC7ggfzIbtIH2
vvo8MFAn/2mSWbmpyf6R+2dV6P9hyZ+vzBqpmZt4KBpnH5vEIbDG/pdPr5mUu5Zha6eLIbF1/d8C
JhqRhp0dIgMc6Uv8EQIbDMXeVLJ+N0Zz54NEAiG1+ZuI4NqG5eDUmpYQ7Qnnt/EZnQ9kHcDiDfiP
/vNOsIDCcR4xmT3W0ygGTMlzVt42b3ErwwBJArEzw8FVJCLVVcX+zKtH+voTRd7ZAxuek1hpKg8A
8+XPX2LqQ23iMEKkXNFZpSNqmEvWE9tDqATiYw5EhgKl2036kmnbNT2Kwfsulp3AFjIH/dyBhXCW
//e7gxWVioBczxwUy9NkvywUMZsrjKozlKSfmVldkMgcALuEVf2xkbvIxa0m8Gc9ByNwjZz5+mWE
uwhrVFqD7MQffYUcFX9Dn+w1jLbr9TL/iZVXleuLRAsxadUOS/ibFde7Evb4y/KwPyRVdpTo2kQd
Tfm8YPBXSSN3xjmDQ1fSVHGr+JemxIwAtaaoalBdkZv3Sr7Muwane7PIM10C8pFx8OOABY0J7zhb
l7G9tRptfzMhamkxkkh6O2lDMBaTZt6BpJ13EhvGd4g6+8Z+Ee3hlqevHD/qz7db5xG958VN8J5s
jAGAKO0eEVHdaFtXhXHU0teWEThtqAlXlEAU/X0cIDwuQdCMDc+uyzqMBDfo5Og9FTsvUrPXMb+u
WvmkYsdjhUwMxCiDd6q637YReEh9Hc9Xn0b8v4KZbpgEVq627vgnvzHMRR15Sz2HwLfxdoCB582v
bjKnU3V/qgxrwpeinuhKGkhKe+VTRkyqu9SZU3PUvdpqGQ+u4XS7cCMSeR7r8+srBZqYVD1rQaa1
WjJLwt4JVLRL1zJ3egyu0Q9xnflcITyUaySkmZ68ve8F7tUOnk1mXD+03T0ZgR5dlwkwJBmqYnMB
FHKQDF0QkDpHk5ucKhj4iJCzf4blsMetVNR0Ha519PIYHLnnWOzFvMTUw5PLF5EWF9PRCgYI3Vui
3IfTfZEMkLtPU3kY+RJiTgwwH7c1GHPXTAKfciGJoXHh45Lyx31+qx38017MwAU5fjLRT/V1e3+7
IMepN46myrb4Q7tG+bBMPbqGmPDtRV0ukCeR5Frkp7kc9Z7jlO7gP5V1Ai0TXhPr1l1CN8zrxdLR
ZlUQXdnLJC1FdZHkdJSUETJu4YugglQtcxXD7vjpjM95wa/hNIsCRtXWQSsn4dav6Lu+qu66qS0a
4tOLipAMTbvKrSpa0xtS2GuecwRZt3gBzFK1r870Ydv91MnQfDo7MqrZh9ffwgqk9gGylw/M+q77
jO8W+aZ4wfmwh6Ij269gHxFrfN8/qo2zTDRHA8mioG+DvvKgS8mn5ObVtPhpjOlVIzCbn6TvXweV
UeJiJTl0VJdJWgUr8KFhinhxKbZPhSzP68wIO9Gzi3oBmEZyQ2vh1Jx8cjMnEqoNFYlwzEoFmNnp
4kpI+CTqLg33iDk6OM0+eFndurObmxQXc8m9EpvZb+CtFldVqmIRFRXhrJCeDlMWw3xnXTs42DWe
8dtbvUynLJivudaha78ASt3Y/sOBk6V6zSkTSowcNStVAfvo8zA1Puk7poqmaAree/skeCbSNV4B
07S90gCLcJYuNcYvEAWnAt4IDn1KiHD+XFqflBdi6cEBeA5PaIGGOV0dsv7pRlBhnm0h50HIlez4
LJuN1UAiW/n+BoZ6M92P1RgQMc8pdJiV5dzc4moUjt5xh1kfkFtpZ52Lc2ujq522Q533HmuJniZj
MSIWzScB6ThrcBIuLq+oTA9Ez/0ppqESjTKrDZuZI+tRLM72+tV8Gi4AdJtmCP7KfkWk02KIr25p
dbfClAWTJldu8jXZvjNGE5jOiHAJ3v8gEFTyjFmmBLAgWUnjQmVZTXkp+wnejMgLm0APNd8/Rinl
GnLOJBseRktmORepd+4RkfdFwt97pT6a2n3QzOIEPopcAVDFrDFVDKZEopEtc7O6Rz67Gi14XoKy
HooGaxUUSOj3Stw+f+0//I1R39ULlrd4Ny5qt14venIeVhIxPmnGN3m0JmBS/xlTQG6IWpoHrY9r
iyFHQVFJJ43G6SqPQDkfNAMyYQOGVi91zxOExdaTX4d7krxfb3bqfsVe9oD6fypl3xptJiFITZlo
vusLTDLbTTL8W66IkxO4n5o58hngJd3FWBT8RnFnKh2LZ8mjHnAIIIVh91reLmgsuVos0LQDVD/X
oJ28UdgtodUVo9+z2agqdPmA3N23wPYt842X0fbvvvBMIPlNYmYqXnIpP6kafsk97FzFmDBqEUr1
Pz0WVy0dd7a5lX4x4y2FbmKLykl9kymncIBqnjg1TH0fv6Zer5E9uQESVC4sGruNDEVCh5fsTL86
suyRmvrI2QDFaTgqG7TPVUQQRzcr/n7SirzEaTc2GL4L3YHuzV+H0CJlMEw/kzTffou9DRDaD1Hs
2Tkk6SLlBH+sUy0tQrrsStCA/w+V7ioYTn+IlDdBGl/gVn+xrF6DNi6AcVyjOEItiq2VhtIiTQ/X
fSVihgrG+jPpSEgJ7YLUGOKgLdWa32VwG1EoqHEpWuFnrFb/dMD4mQ0srBbl7KzcW4u+1kVsGPo4
1u5jKFSZPczv9k9f7HivbZC+dX7aaYXYe3imiZgWhBb7Ex9GgBUf2KXN/esmYVKKObSi7l5K+fhB
gSACQ/BGwprCtxcG+SDV2JBTJbZiveERKjGnn+1YkJTI9XbZ0zgscIAPqWdQS3vKCg85m2LO/1ID
ZRrmq2Czh+07Tyz5evylSg5QkBVttPFyyWUemIyaLAMA6CU250OW5UC73H11CuxosdptWcuuycY+
9u+WrGfRYKESj3G4+ERxs/pNbFTKTMk4j5FAN+2qkFDEJwqE/WxumH/qba/lQ1VUTtZOpLUDIBL2
93cOhHEHbaymSc0KPWhAQJ0wPLpM5aIbrmZL6wiPAEvJc/wsGORT/It/EvMBY9EIEow4X70fZU9T
GnnreebCWk9zQmO/vFtqk6cDBfA4/mRiqxGNkcHnvCbyh0KDHxim0iR8l2o34FjrPBGVbSEO1EGY
P5S8VUusGCagFNkG0s+PyRNvwjTyeRbCKm7KuOLW6b/RGoM0DO/odO0cH1f4WNUQQTk6ryMGVzjy
m5kABLL82t++XoR+xSkhqsWzDGzeyB6WX1W01STViNjecS7zJu1q8MU3t4JkNRtwnaPCA2pF2tEp
NDjStE3oPeFaamjp6E6UiumbHFQO4s/3gnd/zvoCKKc5UVaH4MHmZ6khGPK0cbJ5U4xXXndmtUO+
wQ5JIOQDslnM7D0uHGja0TAinEF1WFDyrv5tCQAovc2NITrDYL81+1N45dq4eAiX+r+8z+AIJu1U
fw3zOf0OgUGK1OP/RVxSfOHJiKrPh9vzvosFLNZ9V5uyF3f+4TpSZ3tdJhSFqLNKX4I77TszjEQw
JHP72hA6AYinqclY/lM11Z8AL15tqiLE0ZgSjP6vGFcKaky8vYonRaFL0krgHkx4+dA+nBiyqiVf
a4aetF9Ko+X6w1dJbKYbEc0PObhQPz5n6ZVNFRqN0Mp/q+E/noLgdE09D3Zxxq7W1r1CGsARx27A
mGlUZfMIyzSYpV4Ow9+1XTy1K70ADgS1kb0wLotYYLlU261kKZBKaHpqPK+018RYkFJGBcSC5+uX
T2GhhHWEWZEp/xKn6oPsTpq6Sa9C8GIdP8OBOx/CVjS+oceRV0chPoZWOU1/jL0n0VOVVxkjLzbQ
vjQdK+A86+XhbbXh0cQCO00QO1QWkhbRiAbTDiHYYwK52F2JIA9nDbOafLDnWdGiFXBeLGxESW7s
qgvS6B27VPJ+TFCEGVJeFUkHAbV4hssGFXOPz8fiZWFTqDJJ0QjnVvkzLDm9natD3WuP1YDml6ah
6DBHCOsMxiNYtjVvt4693Uvq9s86s7nvnf8rKtMveTQOFKqi2vgIXXSTwkrLPdxpjjIYzyapoJxw
E+kOVwKEf7VVHc1jUWna7YXWilg5GQWucwenRsW+E95UDTwYuTzysPux4y57KFHiCts3Jcw0NpVI
r47C9khui9uGz9pVU3Qm/zMG3mQf9oQop/J6fgVdNOc3TuQUnMtldEqCdN9JXBYt/7wFvoRmJB3l
1sqcxhwfU1i92zcaWuYxK88VTJ31s/nDYc2euC3mPWWodsuvg4hOfvvRiQTqVe8w5m2ci3v9wFpR
tHwJeUHRt6K8NlVP5I+qQWYeiIveo/b1K7FSBpirjW2Q+b3NkpeEoRHs9/rhmtNQcyQP8Fj4qvDC
4vLeZ98pSQUVI82N53WlO5L9dcRwKwuVrfSSDheIbbaJ9k7FAZQVHXFzfsTDO8zTrLsPv8YebRWe
NGlvxZ4beEtUohkr/IG0G5dh7xCyIvNo9+ez+iRjTG+VfAJY3PEna7LqpsVhj+rt6ueYc8xj1cm8
ryam0GOLDAOx9L71/q8hkhG7VVK//5V7r0d/wIzIVfBhoGHNh9eUClMq9+76yR8vZc3ZntRimJsS
6o9J2YbjleiPLzpmfjAois/KxQTHFRsuF9HmTC47TzBFAWgl0VFt+NIT2l+sxJ7ax9ZsValcvsLh
rFx6QgJjDPh1idEoJ2TXeaDqxB7bH3sRL3bpi6m0mi0iqq1cufxcSPPXz4wVnD/T1/HOfdHG788D
ahjcAlcJ5jMOFzm4Cbqt890Q6Rl1UyszAyhORQR+d52JNvXKhP8y/J5gLnx8XE/hUhiIP9Y3xPn8
jo7FhVgBniUOwVRjg1o0b26d6nhsut4vJNS+CB2F3W5T9sj3VbauP062xMOXlr7iZrQdqGKLMEMH
IH4OrX7tY0yOy/D0N9lCX6b2wIhVN19STMGsbwIG/dY1kd9V1EbVQAJvefqqI0y8tLv63FWcnJbV
AisfwRRNtYH6MPVLmcCS9F+fw1GVJ5Jw2jaKDY263sCqrO1vFND0HX8jhdPIWCzdvt48IqfBhYKr
pUkjLhVMG6NBfNMmefyZ7viuo1UiQppJTradAiRwb0KK+hd1YoCyx92IIzq0k0xCAJUgOs5cBOyE
pehGMVdZeDmS+UxvA7OrKSyD6UpLb49bXvZa9IN77OIH7J/nmWThdmDrI0+iib2RsODSZpySJcqw
sK6ftIykvuRdHzAKd3o1mE+xWx3p5/vU1DtxChbeTg205Ym7gs1NyxV8xr26kvcazTn2WPzcm90u
Ji+lSQabyOsZCaXsAQPtEGlIUuN3bmZ6unwZRcBvcUUfJ+CEIe5OvbJzPrWnJRQlyaAeSPkqJxMP
jh6JfmRVNSO/2CnkUw1lyncUj+nhiWiePi/ST/6zTXV5yVoISi4Wis5Tsgdvh+fjI+HnMW4fCOy9
sFLL6hoOsbRc0XXrepkZ8vG9HuP1+qyhRR5OE62DoevhDyXqkfP42lem7vQVxiWgqD4hWbeY0cjv
iS/mFi80kYJUesdfCJCwlKy9KNiw68TY+m8fCXI3H2ttQymQYUtx/5cA+gvqvjg/5o7SNGQ6/wje
MQd39yGjc2hy8wBXRBucaGisvPTrnUAyqg92kKyVCzSyWHWeSvHCdmqIPFdhCHJX2R2P22pxojVT
H+CVNl++ZkKMdqLaQvRR1B8v/zVCr47GUPQ7UL0Yha9gbnJXIjiSCgqWPa8LBRcoBmzy822bBhq1
idu/EsIS8T9ZNoMYjfOn4Y3MotK95CjuWBtWAN+wZZmHsd3j25MOtKajZOVs0W3tJmNep7l3opNs
uwZ0Dxff0ZkJIC/Rs6u2KCoC+tXkVNeaJ8Zl8yQEaqgChfQdFrzdKoDVczw04QX2XZ0++6XSHvKd
+F+TIgskkklZ4o6S5QqOjS8rfPVYaMnfRiFyEZqtkPzg3oEiwQjL7TbJ8BxX5f8DYTklzpHKcpm7
XCm4h39ceesTJZWZ36c5S064bKwClwCQmtyr4WOPieU/OKxAtIOReeBDA+VaQZE4D5z6jg2S301x
DdIzYlRcCnaY2Qj/VPixSMfgOsmhF+9ddmKsmi1JQR+0qOg+Kud6OY+zUswBUuAXhddNgS9P2cxU
eq8Be44Cszbgf25irPdReAeWm5EN+k9LY5aKeX39El7T7Q/X8zBeqblG1QQNMkyvneTBhz75Ld6S
pinpXdDp39q0Vps5ENAye9mjf1QWHF9Br2qaeqvK0lyOnozpHPOt49Hi22mHgsvJGM4jP19l9WBE
QTLaNM1yI0nKzYsCpXMQXNPB+As9lowpDw3vGjMjlJDmHKFW6eLuaMfEZgttWP4MfhFMKT00jvMf
2F7KxPcLsylLnpBwdLlIjdYle3WDOdpxalRO6tzjh6RW4VRY2FIyiE/1VDeSQj2nX+WAIEaYwp9X
D2W1/DnPEjcX0gj4VQ08UqCLXBHiYg6pmsbeLntdwNlwsxxbg2sQ+/+F4W19hLSXa4UnRvtuW65q
QP0C4Hyu7RmEshRjU24ccw2IEpz6ceXuxtmiQqKdsWcVJKl8E2bzb8H1R65pz9nCtBAi98jY980b
aWq0II/OgUn5LcpcvkMtLMD/FXyuELgj10nV5RuYMQ9L2AnKGT2p3qvUxm6UuURlc38zQkj5N6ca
wsh1QFBXdiidEP5sJDdP782/3ZPtRXminWP5Xisi5U+aOLdoZnv4KDgU9DMnY0aAKL3aKe/oivHn
IvtNV/YAihw3yphH5Xec92iiNbstB/asd4rpaUubzphIPA9+ArYVDlpLwb2umSgUvjvqRhqFvNeY
oGuUYFYlFFH1J0RtWat8CRhHh61oSms5EIhxn05oqEHaJNEsOFepD2zR8N+P7dQDk/utWWdjnjBK
2+hKdC44xYgeZ2MULdcIWsazvV7ie8bWQCv+YYaKTNZPxuOJGLv+xCBRxPzQJyfIOOSxhRfefxWd
/W8luTu13QPjrFzjTEMOWcsJRPbgVYiKkUtLYb4UJRT75V4Qec5m2OoNA8UNPS2dA296CmVGyPxY
YuBP/vT5EF/oPNPftoAK+7N8IukWo4gW6JNQ5VqNLLzXGVAoItpm3L2wy1WLJAYLSLpy3tFsG4Ii
WE9NT32Aepth1YnvCxVHd9dHcM6mLX7X5oFRHcnNalSq4y4DqBol5bHLu8xnv6hAhWhKTTAfEc8/
71SIjLDuY4FjHd2bF4cWnHEWGvCKi9y1kn9MrqKQZotRQXtXI79ItG/O6zjo15R25+HFn6KMgS9N
IZW3X+N65fEB7ya2c3o+gBHZknzmiTazvtyOfCJb3GVuJm+TLNvFQ7qRgMydFUTr3IamdPkJoMaS
CJRXTPACyOqURGCyqaf6d0hkjzQ/zuoz7mp70RPP460fTUnIjI0zbAOnNh3L0up0FrrewGqmB+aj
L+0xYAeZdFNVpa9jGxVrnyYyE5ymdBbnNRRskkxxiC5jovvkfS0Xk+V+GfZLcqtYoXIt/uxhy39f
psebQfGI5TwwWfN6GTPLZ601ispxFbC5QN4YnJaBYn+mxilM6KVjEOeCxxeWn7ngsXOZGd4un2xp
CwR/qG8hlOnPqVx5RiugK46BN4V9T2s96jF43Va/tSJ+IJW3QzZf8o1qdSsnLmvhX4jJtuQq42ne
eYqE1PN9adqn9V7T6tu2n1RuWvItKTYTSlUKzZamiGutYg9+dk7g8gyg2TOBb48cp0cuwrB7iYcA
SnB6/djuNTbwTe4D1BiniMMV2yTT14Y/ED1U5uhxeG2mxDwMW06B52cYtG5+TsZ+CEO5TtMQsGJC
Wxjorlhj2RornNWd4e46sRQBkzYTu54eLByMc1olPLkAyjtlHZBjZ5Z+LEzOjsrrLDoRl0ANYuHO
joxib6eAjjGm3dvzKwXQoxejTFO/F+3qvhOJjOKHS7nAAOHaIx5eNeTr8RFL/yzrkp4EFesk3+yh
Yi+riTGeobZ608ViAFq252/sBEDt52QL1CNaXABwOMyOXtB+3/0qADWOcjfjw8y9WR7do5tDuhpe
wwi8fwu4dCV1ec2RUOgkaR0nvmOXeDGd91br/1TbcswUJq3GITqm8bxw//A4SGEPc1/roghxSwtA
0ufYjdI6FEaBn7nEABig+TcKyM3cvc54SLXex58FUXs2vf57T/lvWckND8YPyFnluvhbHeIDgiD+
3TwjzWPn/ngIfZU8n/K2lP0VDz0h+pCcSx/RGq8jao4dM9s4FQMEWJ0rz2aDPepIAYiaCkPXZemy
Xwe9R/WT2Q6flOpOTMP97ljMsp0Q6n0U4krQijbPjmtkM4qFlMdYYavjSJb7POe4Bl9177T/lvlR
5lKokGT6wf6mbw8a9uXeJJj6Zpoo3oiJjqoz+gLU4ahgSCHiBfQ8yEP2+FvLGZ5Mt4svL/QYztg5
YhJQt/uXuNs7H16ay+jhX+yxyJLHcq4VAsVswMadnNrKzLNcWZFGixbfZriSn8E8SlCCRMhZ/Gkd
vF6uNpZkZDVjeCpJyvvHhdxDb5kaMUkChYZ6jXooAkzd5lCK/8a+kpLyo8V8vKd5dFYIFDhmBPWi
ed+IeKXBzoOPxZjHz+1hwyMFcTNErk2AP1iSkaT/kPq7X+FVCCXuA5MgRClCtt5arhCbYU0CsMDr
JGNxSO25ygvah0oCJXh0ksBa5QszXDtiHzlPKkZ6vVRFroJis5vyPi3B+ZE8BeE+7lNrMJHkltts
/JEzRwyoGQMnR/4RKG+Dyxk8r5wZMDK+v1z/nGxdyqT8sOMmyJtgZvtLsu2IfU++eMHYdKqZZwL5
KG4+cKOWqaYKXTr8oxpvFm9ppK9IyrHnN11ypY3cDvmmSu7HMwb/i3fZb8vgUvLnO7c+kpJPJl0W
aYPN/BFmt+1gSp84cY8DCC1LnfJMJ3CLSsNvfsTjZzW6S7IX3o6Dn0H/7etnlDGAQMjW2BJLYsxh
gIW9RGDHlduk77e9S2yjogfdgwYL1Fsd8bMZVhYHmctrGR2cffbpS5WagVPGvBtI1PohHZ7GF8ev
x0yAQ00ATtROdvPUygXmY2LUNkzInpAQ2xWQWvSnBTIgOjyTtEUWUBRWtEUsLtEdM58aXonQOhvw
ghAcz1Y9H1QBXUtRoBbdNnAbUixy1gmaUiCxu4cwIg7kBtZl1aZrxsTs4A8xehvBWjKQetbKtyw8
MTBAHM8bn0dk4WyApP4fwsr63f2cyNn9MGj+fXDvX25GQBybArs+A4TT47TWmcC5tlhJfNa1kqfw
qjd0rYdzfZ6hy8qiAE08IZWNyHiMb6AXG8XATMn9OMVorym0/9N/ynSRVcmgRfrHhechbmjGx4TA
Fa1aH2k46S6glGSRS72efwf6p9VR9zh7V0oSdLenzHVPpMXD48K0nDhbN/zZMbZciketFn4kAtG4
z+Z0Dc/gm75eMdWotcv3CJXFgQQ1NG5gxdwX6EL98tljvD07ziqCFWAoq1WiN2E+/z3xLRlI1kk8
7kpi/uI1S12Ux/XornOnRbw75i3bGg54xErDohyXRHVfAZ60z8+NVKGUi/gA1xN4wnbAstqexvck
xXw43ZXTwbt1n11wh9/cZKQmNWbaBccoINMVLUa6Sb6BWHkauTHNXWhI4v1q/w3K/Luq63ZSltv6
dp46/pVJSHGDRiC0EaaEoCHUGo4M4aBt/VuQQ64HNDj9aHljmNWBb7ecIp4xkl9j0m14S5Ael5K6
kxNKHEzhPprwtAqwsNd5OcoljdQEuJZ5SGjqAV6mrnLYtqUnNQWZPHyvf2NBR/QA1H5+SllElvcB
3DNwti2mBSAqGPyUC+RzF1OEb9wPYawAKNi1wzq6vigNs5Lx9LVN/wYu5JAh8sXvBQ650OUBay+Z
8LUGvBUR+EogWuEbs1ZnsVXw8LhB8zMJF1i8mgAfVBavwz5PyKI7CnfXmNO8MhubZfhrzmj5jEcY
BGQaSu6TpXYyaKwEOINNSAUGwII2m2P/91cdfBQZlnMHDeljB5RrcHHUsnqzp7p4K7GXuqhAdhUY
KrSuRRzCpq9eWs/FfPh2fDp2zpB/TlyMuu/dtdqWKmAlggNz0172tgUub+q41j5QnwmJsdUwbSmd
+D1/8G7RngP4wm8oA6oI4yDhWuCQ+6wEm6IL69cnWa8tnQvCAIVS5sB3akhl5vPrXJx/bHZ/dvuT
2cLGmv6JvJcKYAJzkcTO+tORzmlZRFYumId8lxmBVG3FN4HlDw8sqixUgZ3hE7X+Z8n9BLawc5Zg
2RLx/yeDQl6VKrPnYu2s61bCqiHM8WhqYUVg57nQC7tnWQrmhd91RTdTzuRsgVGypslJ1rql3ERq
CVX93kRrMK9bm/fchacv2XV25bondjk6Ux48vcaJ8lm7fpE3TFfdAIe7Qy+Si2RY6/h0pFva5HjF
IV7La9f2sftwk42cp/DgOIyss92GL8pMZjN3U63V8JO5oxH4BbUcpMM8tE3hETr2KrVOsGbP/41O
q14g+hA9uIeKMU58QTbiV+COzI21oYlfddwl0xFaffVTwWG41q9j+jCiQIxTPC695hsN/sEK6ID/
FIJYthXZMj+b0Bs9mZB2i5I+jld6Jx1p8ZtoEVaEb3oUsZYizgBa4Uj7CuOiNG1OYjilVYACqsy4
iuhNumTcpmQC/U54/HxmVPmsd05NNKnxYTXjmwDpV/mlNOa0ymVHwLIrHw93Nq1q+dG4zX9sxkB6
D+hcTXHxuJP7e4sNLLTrZM9bo3gODofqdwr5kK5x+FLdVogDYFwcOqByaJl3NWdvS4ujbg5u85Xa
ko6pHNov5CJUYD2w15HKfridz2f4tpig6B2ANG02neBZ6AdnVoW7C6mI0lt8U4ig/wQ1LQVImwRD
OIBUr3W2Gpi3ycL36f6bxSUzkyKUlYHw6lYIjkx3C+VmmsndSPsNqmzw3hnZjmLUixUOfQOwCcJE
sTZg/9M16Uu8mV97ZUSrLkkd3PKy+dXYu8eMs1fXW7EJGDvrao1vbgw+8Z7VF/dfBVxmwF5C+0mz
9CUShYWi9tmWFkQmXtAb+aGiuncPovF8WL69uljkZNbIu6wsWm0tXiWkCj94cHKbaeaWH30yLS9u
Lt0IvYKDHLynTOgluEI+SZ4nVawnLuQj5cuFcuKXzIDFx7FAkKZXuQF/Wg8u7qaukmALrHMpLNTf
jAfyjzAQNwNKV7AgMT14tg/8GoC2dBW7H33Uw0nHNBk1ULrDmea8zm5+j4FX0Q1EJgKUic299YJK
FIa8Jm3KtZn1koIeUzjiRqFNuNe/ePEeldvLSo5A5Wj4kqr5TWzU/+8g3j4q0EwVBvddJBAFqx5k
ELSzrXwDy1eJwBa3GlOM7SnEpnnbk9cuHFrs5XYdso6VsLt8mejNyQ6KyPWTMfCmzh9rNNKPvYNN
R6z0pqwCHChbwfVVtDs7EKU+5gzxMohH7RU/5i9SEBoLP6M0RQ2vNX9g1c3/B0d+1ESOTyjQiWL6
079vE7OHNUb+JeglMDOKB/Ye0W/st7YZpTNCjGCI10O8QRfpnVcy64gHI76W5k8SbLedQ3rc/BXY
jzOzySCvDAUf8Drnrch+EWzh0AkZOicn0BuTzaNwlCSBy5HACvex6uP1HEdqCQmqJoSpx+rKO3mW
RBEpti1/KRGtNrUZ1PDo6ChFRuvFcweoVrqvZV+ls0zhyydseYi58seGw4hk4zEc1wrtR9h1yTuN
UxoR7jPYBWvO6nv0VhYfhZv0KdvEjnZSy0Ub00ng/hNHpOrra5KOM/00KTywhCK7VX+Q0cKIMJhC
2vN6KSzy/d42d0JWA9LzzJAGD4XrhhESN5ivdjh2KVL28xQSvAaKdGFVMZkOZHzErtblMv68hgUV
YJDa+k5uLvVg5rZuRi1ZKbZQ0kcNsg/X/UWbBE3eopyjJalRUqlOsSrNY/px7R0ebUqapqgP7+gH
ExqLFhXiisepzquxkRMB+jCeV+JwmJ0lZPci8QjPKK1HfLWiJzr7V3igFmcul/Nur9E5kkADUANk
IrvWl6i18oGWo6roMe/j42ubXq7edCYddhsaqeyUCd2PIoQlCCVFPXhk+xvpc4+g6R9u0KeEl2EF
qErQ6EE87YP0tR1oG1weUkHDsLOiBTsnXq0bWMExDjox/1vW3CDfpKlgAxyHlUWLA8sYXezebWxN
C9tVYWWODA6GeWDBebGOp8sHrUrdd9Gu4aRFXBvI33sGhhUOSWW3c7HSsoUltPYX4iWG42aJBgyY
wJ3WqCF8ma62qJ1B9hSLLhAIvCYDaSAINMytGRyGjt/zA1RCv2dhk7yGpfRi7nYccUxI4pW5Lazw
GMEZmlRS1h+qHel55Lf1E1WctrILYq2AUrPN1YAuW4Cl7DJsN103G9F7weWBTMXERggHVcbWphTA
VIADy/FA4i2U+Qiv81/d6mwvo507CPDOFunRFd7ziQntrY8j0DGXmlAIgZ4d3757cS2f/jC7jhIv
RiHMkv+JwxC23OymVcY7PVJVXtdCcLBFYaXcUWdD7bNIkLYx7EJPdpXj2UJj0ziDIKYIZi2noAFB
9WbyEPSfV5DQuXQ2cFgx/+V7x4zNKkyizmzCf0R0c9SNdxShHC4LRKq8Gu4IBJMqRV0K9IyMMHoy
zpUxKLgPdOI9D2mYDL9WJWhJM3Y5JqXgpv5vBck8bjAFRTF1rJ6ya/DjehSYFBena/mf1U8rspwH
UugSytOpVpuNXDlD8eTUOcNEWWUymUtlXRTdo1kyWLOawWQHgoskynL+IVNEYU0ydV3a/4XPick9
0H5BEbQfpQ3D4pnkmnB4SJu9KgFcTdbnVmXO0EfM/O6jTPd7jv4wUhmg7oS8MCPuYJCdgU1B727v
C2egB+qB5h0I1qXNUS1jMRTybDKt9EpOVKiMY2UZnvOOSppKwJcBbFh7cZQQyIpVgQ10Ji17pcK4
GCEaVnsrfltBCpfi19cGjOqFECXWbhHB1q8C14bb6ZJ4Q1tH4ghVY6IqJ0BBwlA7k3ONaa3UDSJT
jUEa8yaRQTv9g8H1hPj4oF/tZMsGlspBOfWGqU1AxY9qg7q3zMmrhXmEufk1UDvond6Uf8KRn/Ta
a8XOzLhzOkut8yeqFSPPiKcxqX9n+pi9JMmfIxMy57j4jEM2VEKkCXG3jZh0Dp85u/x3Kjpsh4Kb
4LziLq6l9oVmYLT9ygDSg7SufmjoolpObLUtY40LFUsZuzt5kqfu6d5MAb3lBDkVFtVRPVR62SWV
14xItvzaC/LywEi5g/JS7eFLuxrFBqjATAzK91qKALbM8U+09vUYNOybkgH4rS9vU1TB0zkPVev6
haNKcmgYmA5bNqGuhrczDNQ0WuoKzRRBsHiX9g1aWrSTbQh0/MPLZNSL2Jobpm8BnzQ33getqIKf
XanVhp1nP4UDjd7e+NiagOazpTv1vSbuxZaaQ+jwidKDPl0gc5qm/89sgfuAqF7f/R4QxjQ1Xvr3
Ng/yoCDWk/Azvgy41CxdVpHkBY6V7RZnVtzhgIrBWsoFsY0IAJKM3RhOqQADo+ASof34L10IyiRg
YI2LCMXA/nkTNxvrEiGa5brugH9GmjDW260YxKhDmN377GjpmkSeAMcsEo7WjhTjRDNg5JFlgmIi
XWGkL6z9D/7UNUMypDmxXcF4PTuF/RvgdBUrxXzXOQ/Oao8QeAUNgZw+wy0irZ+Kvs7o/kFEi8nH
7l9zu9jXBkxmwppIyLkzwgTgWU++XJ0WA2FRFD8XiA7AFlp1BCCMkfaeVCHhn70cWqa8gC2zJci2
SK7QHGBLQseye/KtGs44ex+zi8yrgm//8NGhAzsYxbIU9TKqLMIKlLOFKIJ+gMCBifqpLL0gvuLq
mTZQg13U1OUPFSH/nkw+yF68c+GD+I6+1elH13tzN3m2nX7cCqTYZA2qP3zKVTcO34SMPJafUadI
+8pax/7btuurMz0WRAYHAjVNEeAH2r/XVU1ybbUR3kkCXZwCGR4lHUzrO/D3Ckr2xvZq+ErhBkLl
dv85AZIFwO0CBZ79nxdlk/Ud70Th+nOOeIJMDiRbAKib7XxPM+ye5ZYAKvMs6YtEtHDLUaiKpRDa
BbCgqNGU5bLJSS0nLLydKydtN4qstXvhMDzPd/YxFCHpdx+RQnMMf3dKHrN8cOqVCoTlXKqATj/t
ZYP5uIOl3wcYbTSsw0II6k0zSOIfQooyXA8NRQcx4fAus/EEkwtQPSLvrv33r/KhuLmPJpAFonZ5
TeEAb3ZcdM910eGeXiKCg0u9Xy+BIxM5ZLA1H5euFhKg2oT0lqYWkC5ovw27SzxiGkpvdnnNbRMv
8sGDPHeW7DUc5fyt8UZG/ifyDRqo6DX8dcjzlx7BC7C8FY3p6k/IWP4ytF+4E6CZAJHGJGYbxYaP
JEDy0gEEvaj/otV9wQSwgESavEAEWPZ2j8DjQQ94iD11VvCNoFVHhdpP/OZ/skkoNEx3BTdY4Ln3
gKSf+iF0BmQ4xwsobJVTB1xAkm6q1oyjEP/YHdfIhXLT/SK04L3bvNjBIf1VPrKQJ6ArBb7PXlAt
hnvRvdtZqrl4VJ6GchbTIaa7f7FqE621pMtUPQqlEDWwnFk4yFaealVO3t3i5UnW3YsPN8GfgsvH
08uHhN64sEy79g1KhdamjIvtMU4MPrS6vT82gSXK0qVxLZf1vub6YOWPmxM2AHJVX7hW5ZGA9a5g
vtgHEb4z7YHGRPgadJ0g56dXM1R2OLbtqr/9gndkOD+kOGlDVWcaekKAxcwqzQ5Tazd4LNsUkF2K
xnqvyQKd17v90DjCtHoAF9ecqvUpQIo71fAF+EbLW+lOOhXz67FrzoyH9h8eUwX7GyJRkTNyf4C0
5EzyyRDGg9YiDn4eUdqT1vRp17uAz46Q9On2CNSj5KbO87oB2E4CD1y6HS+iv0XfYOvj2w31q8r1
Aj1+b8mRMOOBqh9wA0nMzdredAodn5mUBDUbO7NgjyVUTINZZzOeKurSbfXBk4t4LR3Fem1hmaMP
2gaYIeM8ghFELGoYl/dhu08jmAi61ct1/QhjLrgb0eaGOQvrixOk4jESXnTvvQgK6Csj144mCuu5
5iLiBiplJSE939r2tC56zm/NrubSKoV6Cx43e+QYrjvnPdOnYSksSguS72Vvs+p3KfHVsMMJ5E88
vM4vI/EvO7aSJgUDYI/QRK+qCAtInw5PHSzGTvTIVwaBqcGkgkqDr4i0STKizKQE+7esv6K8lNej
rKCVLbTCmYlNVtArAU+wNAMDO0FtOHYswXeEqyP13DReA02X+RrhNQnkYEGuz0ZF/Z/LKOwA0XmG
JTiJYTjBCTqwjl3b6gvv9Qqb2Gxgvq7+KamH2j4O2qjwEOaMOHeBsJB+cZqFSsjyJMKy7EGSXtCQ
1ERsf/qqKrra52Y9I6oYVKrnnaeRfQcqpGLM2il4YXODSS3l3DjsSLE3GwLIx/15TOTud5gRihKR
r+C6UKLgh1pN4v/BRnx7nqkLUxX1sHjp4D750hqRtZah04IwbP5LdZIjP11ubpcS3M2/hgyaHvIz
m4R4FDd0lpN6vWYVEyZu8gwvrvZLEvoa0Kwy5U+Or5lmmcdFCMIaEKYuIfAKHn8ZbHLhKXhMLoTm
CZ9HbBIf8zv11elZwZzDzpvrYXdgMWc4tnyn2565TX5Bz+4UTwol/ZeOK4yOdZmQPKNCMNCnJ05z
p+xL9sm0cs5t0rLEIwo8zOvlThzVesZzYx4FlfXuWU2hBEYHqWKG/EvxuDbcxv6CTLSl/dqU+teH
OWs1KR1QousgAE8u89Jz1ll0RBHEujOdjecZ/6DMKk0iK2jI4FkvXPqXdzuoMrdUK7Lbvo0Gq0Pw
7C+wlKjqu+Uc8BSD8URZQAPlK9zSI8v3rSvyj2mzl74ieqUxJIymGP9G4sSjHExMRSBX4fyf2QIp
Z940CqpGhvD4grCSMdU81RB5iHvMwkyb6Af89fKKND55nt2phP5EuFuk+lAYvoHvA0o0XvUMVhT1
mHMGq7LzszxBrWi/8Vs0avfbCbwlhCHu7Nsy2MrvFymieQdEt0rjp66HhppMqHQ1/9C52Ez1cTqk
HJwWMGi7OiLwcBDyoxkmt+WxBcp+iJ+5EEzYYmDzAbF11tRSCM12Ry+21D9RbSBzGEWUJOpuIScZ
lxRtKrs9OuSMIGdaSDsxaJtch+K0pxUXojvJAoJvt8r2nGzHyIWFWzuh/w5Rh7sAigMyLfBd7ZfV
AVV57uQ+3lm6E6IyHvTQYpuF+LLRMlN9XlkiXhh074nB05n0w67Cf3z5M5QDgXmyoC2APQPTKnIb
hePKp1fVWExHG1Twi0lY4IGm/10k6ZX/tMjKAWMYwlCeBLRFjWI+Vkxvv2nL5iiqy7bq7OpIOl3f
VI9I8rMIETdloBauBrJZI9umhOez98a7ZewquoDIlW4FjKG46+2brky0D/q/2SyunahgD50ZR9Qt
gyfr56acTySOrpe1VsydE81DZv0BaWq20P240xFvm0eIPz9dhHiVcf6jt9olIxWfsHTzb50CFdpE
+JgRy26lMFMO2zm1dRcOIs5cN3TBLNrLoZRRPbhA9n60tvcY/LCUZPA+eoifdI3Nax+u2ZO2/CV/
3rzeOSOnJ5kTZCsiWw6ugCsIyQ2HUb150J6sRoB15YR1fc0vFfHJoq4G0UOaHB9ARlDAfPEWQQ1o
DDeLhcH9SWGGOSbemPNl5e8j+uammpbXMLec95tpMTEHhVMwsS/E6sAEs7Xai458HKFWXEBVPNFi
YdExSIFqRP+purXB22W0I85s8MG+Vf+0pToyNil6R7c8Z6TK2nMd1pHytFpLfXX8Dz1OkyIwz/Bq
KOtjFp/3Chb4qkyl21fszPaIiz668nXrDopYUvg2Yz5m23lMBWQUpjrkuzsmHyKIt+2ukGRQ/4Us
jCirJGnOHcvtBUPQ70+wsVoTonfWHsstx/572TOlqkETF3jsEJbdoaeyUJrOCM6Xu8OdaffYQabM
Ow1T25ToyZsPussxryI6tUBHhIfNC8Jj34aw6AkGeOmDceGg/BGseOc5Wor+ShcMBQjCxOBxjYY7
e0cuq2aePoUCpNk5hIDvghlZW1hhTcUFyhQL5643q8ql6KKFVAGmfkS4NW8/9q4Ta9F0bU86n4v8
HSN6PG/aOKlwvk5YJ0IydyU06LeXlhbfpsAbQ4FNCjqynI3c1F8imTHDMwoB0GNXp401QYpx04Fs
4sR/KCIMlDDC8OAJ13ggOpuo5+f5GaSx7xqVBweU2I7zaqplEq/bQtFk/3R+fqzTY661Qf5hT7t5
sp6Zx1TNYlYXjAtsiaXEM6YKNHZapRESxkUN8DvOAXlBep01qJ9pJrAuZgJCv6Nh90B+LdmapzmK
luDjWfRejqI75czffcT8l2JsWPV9+ns6VDnozKYUsgeU0UDPRikznc8d1V0cIQtsIthuaLzHoPpY
W/beCb7wZUBNwRRfP4Aa8Tqz6y674aGkXk2x8LDDKR2eqR7WEdyTKVyQbeSai36ILGNoLvEfDPev
gOcSjHeZKWcEnkaOaO5GKuMym+Sb0wpRpwaM9Qd+6cuT7s2TxY5LfKr/jyjJROsIRUkt99Tsaksh
M798H2KaVRiyWrtWqv4nI1jYrXp9QezhO2UlkcScBI5UV0o9HqUQ1mAvG8x7TxGq3lsISCHo8CSr
NRDlZJLR9B/5SsaRY/dTAseSJQvy2FRamtGZX7GSulkCvBk8x4ZXhy+oWHYHN5pPKtc/XBvYy4Tu
O+NBkrlJnRJk9gdt8WQaTT++oYOzOdtCHpWOX0yS0WJVOI89NDzFXNte6NRMNdpJPdosS73LhF2L
G/wlPebEDiQR2pLsd+zrIEvW3Vuk4hE+tPckA4g0S7/X+Q8n5V3YZeN5h7BRQfr++N1k3S0RxYk+
iXv4Ji07FYGoeDG1JSZ2UdRg0pSzfB7qeejxGzMRduy8oYK3rgtjbBIHtcSrIcwdzkd4ID8ToXZf
G4dNCIkDi6K/netYapx9ghA48h+E5zeyRxufRl1z/GnqTS3aV8ANbu0VSswWPl7CaIRnC4ZrCzKn
GBnaDLcWCTvJkw1JS4+253atntflW1lgjTSj1lL02YHpv0CpGdZp78fGbuhzrwczWtqGlsDVPJjH
tWbcjFv8O/WLv6p7+Z6LnyHa9GgJfwrl9aMJu2Fbz9PiOxmnJqeycn4vpkPYD25Z8QUnRWeIe8fD
e5l14OHmSJHLSutryqbuRQDNuthLej1xQtowofVTaOeKmaG5jAGZ+5XDu7/slpr9+FMIoVUb5SbJ
bZKnalKrbpxOs6wPEuCaW6XlkQhQ6F/0bfS0DeLZmzqyFJzJBKch7tuoK8FgNq91EMPwdNa8Jz9S
FmcUp/NNDaEheCsQfU7GHJvs9aeBdtH4R09hzJNjubdh5+czCz0zKPcJYZDr7HOpCZePbx1eW5bn
zPqQUKAZz1Jrh6B7tOtagD4tSEFfdrnwIlf993cs1RqDONf1I5aAdeUUkTglCaszK6drUs593kbt
65QaJhrxy3sEPxUZIE0LNLy02M9TgZDc3PuiI3eAaHJkSrPnfbGv0erUfP6J0XSZYuqAIdyLuj6I
X0bvcL/qD9ahYesL+UBd+naJsh9Cv0HHhqk63EAKpKuQyQ8eJJDRQyorFAbVG2X+CyYUzHHeVIJc
g9Dw9v2b6dsq+d7ALYFZP3YgpT6szWVvbkZaP0xhhfydGGadMiR8Dxs81NYxFACxHPtQO6dRsna2
9qRFz8JThVMlJBJi/czxG9WChsg4f3nMKk2F23DbCObz7jSNM0snTYQJkCl2bGBxsiIadAGULmZ/
7DgX7SCQ7yqEingyK7N+N1F9Y7GaMbVckqMuVSKieINVVXRH8BgJKWmFAuedEBcxG7wJpNu13qAp
ozzOGdhJIVP6qzyTdjg/TflQdaFod8msEZrAtJxk4NCLtQaxmUTDekZGeN3ZXnZw+VQWRrMKt1UD
tdaIlMu3VZLRPaSr3T9UOiT1+mLpy/xoGPfJHXNeZM5N8Si3WdbYUozw/JlSNS08Q9e1/TLzqOqV
IrkQUYjYf7BRhn1iOtWID9Y2uODhM0eL2SxMFhohadMHqxczVWxznvHxJwvkLOoz1NZ2JoZPwvsU
P1vQfUZAm5006g+2ZetSBHazqLvo4KcQNVXdqu2fagj8Zx4a/J8fUcrW/X2v7lRKOVnQmQYu7EXq
d9GGqJUHagw3BfudIy9F+UtvuQOMrhFG5UfwNKzjRPOeV2/uw/2L4dk/r6U5ix5XXzwt7TAI8M4A
nHsz18JmOxVejNwLhSDkpSGrIgTq5d6HHK2WA6dAilXiyBI6aPcsHzT0yv6up0+woiri1G5uT8DH
lbVRNNiSYTQOMf/pNtHEs7rQegvgaOcZzwHjsP3rzHR2SjqQ8pf1ARt5qat5u0FE8oEcuNINeTYy
0N0dikvsnoETrg9sS4iPQI9P6DL04LSFLDlw++Hgxkem6gsbsdLLfAhUDCxj6XSDWx0epVYfwip9
EUmNwpz2MnhmgB77evTxQnSws3HooObwbotgLPHh29kP4CY/0vhtrmf47P2gli5yVxGk/TVxBTLk
ALyti9GQjeOTuuhgNVhZqxQqGBgoEw4zkr8/jHv+hA4gXklR5Okxcb3M2SvDOjm8GTBl4g4e6AtX
nJl0X5K8YS6Ak8N6ZKx2VGw33muYdFrlpa6gv/mi45nu68qubrmhLPIvktwb8vjNQnxaWwrDyGsf
5M7ivk0sB8cNA3BMhxR7DgI8B3D0mtqlFu+/um7CXQ39myrfiojjdfY2aLMRv8vnGJASTyFxwP8I
IzAUXPcWAh6Zzdk6L8DtKlH95a5iYf8WGHuq/5ZMu7FuJGg+hd0qBuQJEmm8yILmpiAJds16ps1H
4J0ic6mWVoREv4GtLikBOFkCeoLgodN1gSQHvK/gvtL5U0ZM3v7GM1Rnfnlg0XzHON3SmGiYIAD9
wOuJlUHvafCRKhXE6jZxJ60ifLtI5z4f/eFlVqz4QAJoEPRZUjgjny0U1FpJjW8oit5+BaVPVjnN
F8Dl5BxVonj4G+hf6bqx+bsfFb/zK+GeAPupZyLcyNiXepU6IYdQid0ikPhjmm2SmwTzuK/h3enR
cvXO7VGuzmSVsYV+NS3RtJ3Qlo3EFsZkTtDs5mNIdmLcXEwanv+fmAZEjX5gV1q2J6xX51bvRO/w
cahpc9QtitZBsP510W/3I3JLBFP3j7C72Ki1+VZ5vsOei+8FM6/04cGwjf/H+88yFYDTj3mJauSI
fzhWvLg6C1bpIAulvACxEkYVzup/LQXh4++QDzBaQCymCLVvnUEhvCtu9pab34xFqEQgyC4hIIBn
dE7Ue0jP5NYXzfJmumtmlDTa42wVBUcwLZ+lNGsKY4cA1b1nod1bStV4VzL/zg4Yd+LGeeM6H1Ks
sDDqbKvFtX71+AQx2E5a5zxVRnYzGqek6GOsYeP0KtFKklVY0EgVgDBpbTcatWqd94eYoimzxCcS
Hu9ghQD1p6Iwvcy2EWpXsBRbHvAieXVvO2X2KAkQow9awiJ/yxhGyNqnjY8Fjwt1enWdp+9TUtRD
adeO5qY3wTUBTaBaHptTBDVjSJwxaeQobtYrYPnQ2yrHKRUBPBjdhwUjlC/4glNxxpNOkuP7vfF+
zGPjJW8OydxObjZmpxW6FWSyMlbeRxegXZ8MAxQoPJzMoZFzlWuwDIGme5HHTia8TudIGK6sNUh0
IUC1yNyjwCJt08adDFi7IZIwUDtj7LOKyAPnKIoWSzx7DCymXCBHWLkj9ui0d+B75mmhgq4kpnZV
HEk4ChR7yCac8SX9ppXBfJR8Owx02FYojFdB7zSplpHpzXiWIgt/p2VmuWEeQpdqnlYcdrDg92wP
mgjkK+M4Pf3pbI98O7RwnaGe8Qi9v15LAcMRf4e9yVOiADr68V0zjtBkPwx9zqtIuUc/vvRCcHMk
wd+kdPXNEozAH6qVSKS4S489FBoT0gMpqBJEidHp8aHcecWN2wS08cfykGxhUkOSZZ6s/oP4/h/q
RyeTH+GHzAXy+dZs3Tv2m8n8n6EbARlQ0UHEsV9MY0a5pF+h+N0sPGzwEtH9znb59+iNKKTCB8qe
ik7ZzgwANstr1yjWuyAtLW52sOswa+d0Q0HNYFhGCePC6Rf1ZX+L0UQzf3Jki3xShvhrWJbpf/Q/
IPUXWUmeO0vViMzVe8Pk2RrFIPVuYbbu2qW3s3hBRMbKl8F50a+1WegDRADBiyX60D2+TV9/il5I
lfLAXJPHXDK5oGVXgIkzdBKXnkGTmoaZoX12y5nWKe8OYbPf49GpTlmVMSeJqZH/0B0sKgMEhFKX
Jx6R4w+VzgWEqm/2AR30T+a90XAK0gIUoaOVQhItNNVC84ZVW8w1iB/WKY2y+13GRD2dXma9VKi7
Wfn40Rf95Ecb47ZgSNLH8KQ0SlBEL4p959UHCDzFTrLVJIEZ5Oje1NNlz3iyTQnBUc0gR6f2zc+K
yGwSr5xCKnjDDh/UUa9f//uvhHu0R9QDd3zHrirM07csEuRsmQmUu07GS6PidU/5nC/dlSYk2k+l
5dEcp3V1EV9FDGwNApURadB/UKJljsB9mCh97ol+FXUl6Sgh0RZSzIvI7WUHmlR1JlstiA6uMwyz
vX8vC+FVtyeMPFDxhYlj67LFMbnDaBkDmRrp+w+jho+UMfVtYPMSCVV0DMWihyzFaQEYw/fnM3gd
v+PhLwcmF159I+kLmkbzDuRBFW/7VwvIxgfYbinZRSYnseuoWNe9r9SfVssGSP6ZBKBIRyKr4teh
psvOrxg0KXhEp/3fx7mK2xay6CsbO/VLBG08l9Cz9iUIUl7iB8QhBGlh4WvT893WwBUCX0eg+SkV
RIQqP9iRZVEdrIuHRkcOBtUuW/xZWbVrra0v2GkuQwOGQHQJgy6y9fXk+aZEFOKwIg/zm82Xq5Bc
luaqh1b1+mD2wpTelaWZGHZNzGy2BLsxGkRREyaLEHc2fu4h2F8KEkJV3p4mqOlCfBK0k7pnjhAJ
/TH/AuPyXYRaGNsd61wViLBkRCEHqX6jVkRQwWiVhuBBSoGJhedIRBIfvaNS3Z22qM7oQmW+euVR
R/bSiLDZj0ZiAMnTF5L4CsKA0F3vxifZn1WsuAsDvYrtuzaxJY4vBIImlCLTZ7zcmy5SNymHYItR
+IQ9YW6HTFpuu5wiGNOwxAJxTv0CCa04H65v/J3ya5zfmTEIOQl3rgmtHlnAO9/vzCRTYT3zhR63
yAQCrn1cY03Zge4v3sF5SNQS+Gl4deaZVOMUSuovZrYFvtG3eXVIanCWqsnxdL8SrMxTBepKL/vr
RrI6hagg8Ik+plURZhN5o82IFKL+HxvGu6znIfjCgjMlxV1S1RZ3gytFNnDxu+KIiQsS5J0Wnd9X
dJwDix+jUB65yXuymmUPgtQNCIJnGkH/7gItPPY3AiTGCsdGDFF4sGfijl11rcT3/LUf9FYW+kd6
QOpUTDKEiv8IPnZi/QH9vJgUIPdzHOuup6LeQekSVyIe1K/yjEpTtNBQY5MbVyGDHYMWTZtTnTFG
9/Y5YDZrFNZRXJMj2LOM4dtQWiDXKGd8qTOl/7YYyNc11dIclFZRSarAiNyWcjMpkIGcpZYknvjT
peFA0VbOSRsqk7ZN3kEeGB2Pn/gt+b77Cq7DjOJGNndHqALengFwyuVbRki4pxlGJZu3RGh0lA3/
Odyqh3oLxUmHqY6HbTrvXaVVvcGB1ZRymu7dQ0oH7e0tySTUh4iwmgw7NJMeaFxZAJULIJlkMJa6
ycXyr+4sND1i3TEjpsYEOd1x3nwoNYbL69/o3FIBB1bU0spIn7p1qIp2rtBL52BYo+ebN0ogWDrC
iDlv9Ez/+LwRJZoTEOQEDzgfaE0x+2GuV2RwuBOQAZDT+n09Rja9X7kAl8/ogz4e2P3Lf3lXUNzI
cEQOS1dP70ASthq/EF3b5NP4n1j0JyvgRPJJZhV1DTkIQk5A/3uB551d6OzNdPorPdHr159q8xld
Y3yvpcZJlKX8mQ5dfhHIAFRlWV7kvJ217XfxGC91hMUh8/ZacC39RDgVos5jJs4pLjk7FYE3zhhA
dxI9G4cHaK63Jv05PJVO27osPdfbZske0KCbAThLjVhfzFCMnjvuH4ln/dnzSRWmM7UAWzgQq0wJ
ea2uNcsdbgbKJQQ/ABz6o0ZQJZ6lQC51kzVrzmSxkiJ5bUskubdktE+2QDjr4CIRY2A/2EIAnV3A
MW1c65n7E4yECjfZhnUzzLT8x9JnEigTaetf9yT1ektCD6FW76XapIlTAuDuDsuEBNiROYP0s+gO
wGsPDqMuusOJbIYzvwtAGoci0I5S8KRsRCZIOp71JU65HjRYCR/nTlnR7eELAqQb9MOnh6p4RR3S
UQ+6UIIwyt2yzpAa0wfCeYfSx/JChJ2prl8OjFOVDg1CLA99zdoNdgRsJuCTJvqnCfufG+2Rwh+T
w0aM6EE9du3wQwkgqax/uOkDiDzogE1vdHvG3OaDec3pecTz0XVKrgydtUxZs+X8GxdOP4FI2Y37
6PQUHBFv5luKuYVCPZcyyA3jwR+VFcS88zxhRw5qENUipVnMSdM7NOMHkkWnpdzzG0gbBh0JI3Ok
+Mw9J8sGezAAe8mMKP4G1jOsZ3nE7I9/rO7sf1ZM0h0ucRg3THKqii564XnbSpCXo1zUQklMtJvO
ALo9luiw6ecwRf9RRhod9uvjf4nklt0eEzvSNYtczH7xmSW7aTZq8fNGSSQklj5Rmyu0ygMVeqnh
5UEj+mIsAIvqDcp8yRF65u7DYGykYeHMqU5eNhAtQEPNxGtlzYByTtR42c59nq784KOb1upVUltf
um8W0LWxtp3yuz2SfFf2uNRqMG96sraak1BqXg4IF/Vl1ZfHTt0AHgojInaldkK+zCevprR1sjD3
Yn5v+VN4JdUZ9rgVSnqonBy8Gp/80f7CYMkq6OSo5IYo+05InSkXQDhftLEGR2k144eId7f2+ixL
7zGUB/IWpWgDx28YMAFY+aivXoA4HTm/ilLzO2ktd3eSnR0ekb4WVKJbNqidqPqb3PZ4nuqiRfVH
WCNE/7yE9rwpWLhvryfXNReUi0oAnI6NDO1I/SSSKwgUYAfLRMOai3voPmpdz3sL+z08XZwJqGji
cjPN/Wkt894ogUwjXOuZLGeYLc0yB35yPDgJawgwtQgS+hSbcFyZTphDqsbN431sm8NBpGI/vQpw
LhE4e8jI0UzS6Z3TwgbEmuzAtCRBJLzUtgFpzLxa0tvGIUdxLVYjWyluRBW1nyYduh438zl0MW/P
3PxT5V0vA7PMBn11oGyEtkhitl3R9QbJ4NVoa2Ei3JrMZzyF+L2xk+dCkMsRd+7ygbUK2dN8/oYb
wFLB0Qitjf0VKxXGpYgAiFj/Vt3k7SIqSE9KWPfoK/qn8KLh6peHi0E5wuJ91qUZHus7jyzHq5H4
NE0/2B45IfJM5ir+t+Tcvrm9MQBFUqw9CpxDOP1JSrW+DhlK3TMq33q48HnECn6ssS3CyNO3dHEC
8TVqwiJOUZFo36XTr9PFcl7V+K9FW9tLy5qnb5fAenxyAc0LK4tttoWhmChbyvemIDj4NKr1LOaa
zTsjw5rQDqj74tpIasHkbSKPxGyt/44li2beKF8uZlR53l6waeoec7PLMkiUJq5T5yRH6+GHmz+e
SqWOaRdScJH5rrEwGohIhLVyVGjEu4voYr8pCAEzio8RAqefAZbQED0xVgSVafTNXq4iwduuSqji
/BaaM6/H655woMZAdcTv2QSI7gA33QNDHRR1vzncCYbJt8PCqHQ7+i7DUd9wNIE0cVz/TUMp11ih
ZwFclcj583oqXV0+78BglfuwaFUdwF5vZT/4myn7zj4ASn/slo3OlyCvbsVqH7VoWNv+c47Q0yQj
Nr1Tww41UT1CFj/QMWaw4B/6L6f0SrpgbyV1M2l4jc/mWF6GhVkOnjsGUw04tATBJzsoty0sxRsT
hK2bekpnKPv82TZiMPuEY1RnaY3RFKPpl8TKtkyIM2VGRuSLYZqS20VUjSRZMb/2RWF6rvkLnnqx
1LQQNHmUW0mJPOn+EFRPr9lAy9S627rA+poKwHee6bJhypM19lozulB8BVeaah6Tli1Sgt9or9NV
UCskhJpk67byhP3kQcx1dCPX7S5hVJfxuNboB5bbNe5KlAsD+mig095/w9s45vgKFPUM3qaiFkhT
8WFgpFRKo7BXSW00GJmUhTA1wrTySy3rKAIAov+fZL4rHfvy5j8u/yCZLuvm+mg23/3lG8i6wMg/
K/nQTKEHgZ9fwOhiNl1QHACY2yzjgnbZdp7pS6UrRNgs4NNLLn21Cb/WFsoRjY6iz59rIc8bS1Iy
DD885otwDiyXlbV9zx+QyUMP7/n/Cd2IEL4xjSPO6nuG4tvxlkmLoKbx3jxWmGepNP5pj95cMAGs
L/ym/FLHeyE5eSqfkoGe7Y0obGLdVRZf3AG+yuxBFpPjXvoIXvwsP7KnjVtke8V2F2bESslZsDdD
RrhYhrHmdw52TNYSTHAquumvTpdCz/y5/7BcApajoKRICx/LZaEOATqq7Ed5pX5acy8m8MPDdmmm
5MoSazWP6xem9aWIhRYnMPN02mL9lnpsihcbBOI1WcFK3klUHCatnPXBOOdkH+qqLyv94mtm69SC
aG3OehXcnlQ74E0yjvEFV3tsJYhXUgzf2uOEmry6KsGg1a50/B4PB5rFtCE5IcAlUjpjoD6aDZOB
tUC1W3Lv02hYpdmGzHukseTtGo8Pr/crAbf1N8fGrFZyTzOwpoDmL+klzRaqfKk72+QUTpXl2E2L
dc63LbI0lJyEY+ynZqkT7MBeX7OQp/HAk9Xw2SzgfIwwsloNp3wEKT5ZSjzLdcEvpQBAeqHKZGS6
7wptUPzL7Ks7h5J+lC1/NFqB3QPj+L9WXRrNvUeFw3Yy05Zn+UJKEzokbR1QPX8PK3Q0hbJGL9yr
Fxnzw1RpyczdVNYqTSRoRngy7/L28ermVsYGp2S4O9QiYr4ait9zJWSKwC/621aFD6IBt1NmZd74
TzhM0uEOokfaBoLAAAeuZAFUdbvJhxImrrasfWQfdxbXD4xKR7TE1KMM0opz06E+KeAqxUh+Xmb2
vxXtAAUPf1el9rbqfkBEkFCyxb2c/ZFoHZlQZzzObGZIB0/SNbHdE+0byYoR0kMxRwY15k3HyCl0
FVRn7UmtMmdpoRnrYIJlzxujypWBHpd8FCLnFvn/afTRdTPlj4xPJjaf2b24mWYy/letW+Hmfke5
OLOVJbv8CHGm3vRVJ81tdyoAGhYLqssjoEyFPrK5a4dWRLEfDg16TctUgAXVWhrnfHjogZq/T+CV
3qiV+0hzxZyEgXwSX2No7WiKBaOjDahBrjMlRlSiaKAuvUXQEYu1f2AltCgPyhGQDCrNdQHSmAyY
+F76IHKniZ2sWsHuxYVF1OC3trCGGGZbLlzg85jNz2PJe2RJlxm7NkdaG+JE5Dj1lnpIY4/0Gtkh
h3itHsj5WY/bkKhy7bsD7esn4qRsJD97vJv+sWMxwBMCfuWhbTmXhNSV4Mm4Iupi081WnP8NIY+8
X4/ZKg2TUVZy44sKaIhyEAXhg/rqh6wviFnTXTaWJ9ufUxtfKtXGbtv0VXeRs4MAl9p5sP7lK4j/
9Z+kUZpr4l9c5eXvgmWhgDYKLBtl0dod+8MAtpLyIHYn/IXwSZo4rtj4LBZY4+9IlHmPYFMem3xI
Ly9KAqgld240kBY+CwsmriGDdTUnvUc6rLha/q/itWTY5zXdgGd+sh0I8u3BFTLUiKFqv2tOidwI
RWnBkHx8VZYQyNgvYjNZ0TrVKFDwihLEoOQY3QiHm5Vi6HWzpHgaVTpx9VcOQHvbO58HM7vREfil
KpJLo5Ql7YiY/OuHgSStVkb8E4RezGdEU/eb96fXXqRoxDcISlZEYCpA86M33a7MPJEjIY0+NZno
Adlr8cGkaiOwR+aO2kvqdmaAbJrAMoJHVzgz6qrbPhcSJ0bjQyn+ln1zl7hU7hr7VXs9jMK9B7Q/
AwNxtFz7VSBGhApdNbJbE9GSJpj2cct0p+yQLmy0hAkV5RZZVwj6EfcJ/G1mA4eB9+DViS/Abf9x
gdyy+w2dOZElY6pQK19wJwomCni6RIEAwLSa580qZWZ3k8mdytdZLN8GH/2iiaDZStVS/tmXFSUZ
jEZYit8cMUX1/eQCCQfQZzkWp2YiP6vlpWMfLECUGxQZF+zMbnf9jY1K7O0odZ0fMq2MPETIeFHK
UpUpbKglJ4BfeUGPwzeyU6/+EDyceRIOandSaPaDKKyMUbRjBqPZyReYFVP+Ab0WurZ9V3wlViRi
8z1JEFXesAOR2tNAQgoUNZ1H1m0uTN2jVSaNkCRkF9iKhayCuIbTtUPbfjjzqu4uTcMoBUEEQYdk
PGStUosHPfLZ5I1p7DdGcwc9tgT0cWD07qD3DrMppi4fEJsioO5YWaxP5eg0qJx0iEFvrPc1kGC0
6c9Z7NYhDFhcurmCb8TeVLxI0yPb2xhz8EN/+XLZX0X+7I8UkdkdT0hoaOPEzjc0pApalRXKIN4j
MmU2mFRGBRuiMdkeNcfJLpZsvANzc0YTixLVcGcaeZvYk+s2KhiNB+5Fu9qeZ5gPpRetwwQ30pAW
TvdKD0nzG5LfSmUvDXvkrdzkrizc3Xuxqquy/2BDR2DDgzsPAinMsSt+o6dQzBVJEa2+IhXbTX2+
+aoC6ftjcG8Sl+62xQB+xwg0EQqZhNW9GuH87vsUORT702madq8tUkdtjfUSKFX54nIbxlVRrbod
GTEL4rmnbBItWG7ouXMRr3Ec5PqHizqPEqBgjUoHJQ4bEty0AgbUH6vPqrVRhqfsQst1CZ3yjOdN
19gH87RVbcmmAjWW1y6B5E8QvB6QPJ6jdzppuXtLjdJ81z6YvXj7CQ52uWwneYyToUme2sS/1cxb
5RqciJmAruKVoHCiSoJXBnJ4nWVVvQsu07PuX5oRW1BEwQRC/oQqqWbcGvOXAxL98yCLUqOuIWNf
5UbyAhtQeJriaGTURZz85UdBavTeceBAYjwJjsCrx7oBzy8+JG5iYxY5BWJ2WEcH33HkUGBz0Mxq
xBrDAztHCaopFTmheUbkNg3WLtZIgGYsqRy5kdcq8rBU/sIDa/MhT8/9HJLFwPG3stM+G3CuxV/A
rDRKFUcM+mSdwCcQuJmoOWZ3qiwb9WsPAsc7BrMeRo4Q6SeRhEV5ymp7XZaD76vygydfjGFb97MW
faEMl8+1Ld1Fm/QX4u9MZ4ynSOlWS77C8G2fLqi3597FmH7I7A2q0bI5+U06xa02CMP9V4g7r3XQ
uth2dyf9/bihpPDgV6I+JOegI0+4/Vnkra6T++A//CPmkvSe2N7tg38mOr9PsJB5KPptf0qR+qnH
NmpdrMIAd0MBioUF82R8M3PnA/chwKvralejnoNErIrsFH/Zj/ow4l9WNVSsqvWeTE6ZSnjmaNuD
EhaAlJLRXr6SW/+z0wo2J6vcEgoCT3EsLZIFHNrFtVqEBPp0ibPAAbSd0kpBebtkINd7JpDGYtty
/8ftFJuQJwFN9QMOVNNhs7CGLXnFboPZ9PZ6ZfJhewq6rHXh02KzVSXOWmnMsDmLCqDxyw7tTRCP
U3wXx6E4XVv3k7z3ql/GhKylUPuhjcZkca3wOvxTygSqjZAjcq+tUbsyhEjwWRtkHeJtAGq1pITo
Bb526t875vJmpreLCfnDnRwUuob2AZ6bSGdCD4No3OldODtUVkniM/cyHlwSPv1EhlL11pMWhQa1
jnVnFzvM9bjXxojcC+76yzaalWl89EhgyBtJyDHiTv8ZTrKZfoakQ36o7dJpBELMRQOxrxf2iEqw
L+0WU2+QSOpn7ruTO2Mn3J9wkwjq+PMkxbWvrIXqd+M8JRyg4lRR4VXbQv/01mE36ZbJsFpDKZkC
r3dE7YarocIBbq4zIunMn9kVXosb735oBCs52tzJcs/6UqDaZZ9VGufIaAAPyYwx5rd3VbnX9LB+
0CKsGPp8xQSH0XkFcbg/frfNDuPdhoOqysd/78w9zqrpQqSrFUKrZSUgkRYF8P8qXedVlUZeYo1N
IQuykcTirh754GvUJsGUorwbBTk54KVGoVRUKp7JDRdTZb88FYRXuW6LaACGTbPFdYMi/mc+Wuns
OUGeaZFnnYTs+j6VRVjH/jfYxhcDDOw+vDf6sRlMrxP1dAMOx8Q64490PoD3pk7YZ0voYdEAbiG4
GKgQyNt4E0LgnOQ/P4ilN4MC8K0c/yDU4ZxzAPbijlPlWzpMVMpd1ln3QoP285BjYgsVWOrbu0ZX
rsOnVTKA8exarpzetL/yMy5IosVruLTqEdq9Od6qluRvTEOza4O1wZnprUtWEU9ZNckkZ3B4L0xJ
53r7vZ/w0yTDAc4kq/pmaKSyeW4Mux/5GA0XxKDhl9vcuR+4LmDTQAIV9pJUE9nKRzf4LfA+Q9RR
M1LjB4/p5L53w553cSZbm2EX5q8EATF8NF9yAFIg6ErdY0tH1lp4FGV4OU3Xhl7uLZjgYSqVT+NW
XJqc1b/bhIq7HLoQi4grdeyDWoXgM/rC7Hi6VUCP/Lj+DJg4tre/efkuLjN82V7yeMUqj5oJgvMr
QHZ9UnQAzrqxASZsJOdzX60M35kGUP24KQDP6PjYfbxWInyZdyCgJH+34nz2ig86MJeyfPdfefYZ
heNpoAXZa00Kqj/srZoL5qGMaUZXzFPoudt3AHRhBtwQRdUn52FVwK3dg10DVe1DDTOhcCbRlQwg
0DnX9hYLo2+bf3iyfZfPAik3pJRKIG18gvC395kWbT/Ts1LNczGHrZw/0KXsn4UBU8dJeCNVE7T7
jnGjCKCThwavG+101npIXjKDH8pyXUkCU2585NED8epwDSmryzdyOlnVTCV29S+9f+RlAgk9RL9e
hf6z8o7IJMfTt74UunEdt3u8ING9UCxeerKbRyh7k7NFrur0t8zf5Nn1TBcG97BDP8iuyrXxFqid
I5IO67D9z/NSGwyrLIf8YtbNDB2UvLXax2tw8wcqL9kNQntdkACTFQ6waNRHd5TsyKfJUakD0+Fa
QcGyz3MEc1uUw/cC5ae+2CkSggtUnIxycD4Ox+1J3iAV8ryIAfdkcBNdgSxGotWc2qTb2Y9jtrds
WBDnAreg2ImPYhBJu0vYFtA/zIdhTIILA3I++kkH1Q+Zz4qAqJeL4tx7We0KZcOO4pqS2lagFLvg
cDbhi7+9Z/G1YgDWwHU9NgYkExmaM1+KR/dQg8MG92E/d75S45PoqTQaeLwEJGdEyZ3M558RUBcX
NvHs8735X5dtTSoSgpLD1QF0aDSCIIngguECMYYjQGoU6V/VqjA5CKOmATCgY1lQj7EBcVjLHvz5
+4+26mOEGEQYYSQ93en4AiEK9AgOOVOWUNnGAwp+DMjp/woUPh/5wrc/XVZrqB6tZ5//Ncnr63Wf
7UG+ThuakRrIMFXF9lZbEKJEtb9xbC79Tez4373wV2A3lWSMxoohaL7pqgOeRypUJMEG9ln9yB8E
1lt1KfrbW4aHw9OKKJmgAXYedm/MGjRY7RbfwHNjIsbZGP87rP0wkXqQkqRY9o8lI8O7TYZboM4h
7RWgVfK/ZRg8VPIi3UwWxwBEPY5eTlWoS3yvH+ykdAIEwMZieoM8p0cuPEFsN9eTx3PvloZfTFNJ
a9ZkWHP4y5zaptAdCtyy2LtX13xN+6YMIKfyp/XwyfDKzocnWab1jTOgMn+FqFYLefYWxRAKvTio
TabMQ6RyI3XbZeZE7tUFrgLdHbY1f712SiqHcQmDhS4if1mvPAsCkAQJE7CGDjhKj1KnJ4Q/qyER
REevkB/0TrP9UEeP359qgnKPOCo6yF0MhS9Kw+ClLMtHtCFRnLLHnqUs5UXj5C5bBGwZ7ny+x+oh
J0szSegtHQoXA0wFHpz7cROiKlo0BIyCGODoLsn+a8y4GOOzHD6PBzyhvZxZH0VoEsX3ViaqtGjk
9y66ZvnjjUt8utwXWEgDkQi8hVAzylxJEieoifMUHHDVbuG97A81Fg33bdaZgof7uWP/Lj07snYN
iA5BClLjOGrgQOnOcS4L3uPYylUG7agwfkiYm9E5Nk5zJGnaYC0bNP2/FKirj1XdNWurci4Mdfk3
uJeNY/ie27fmCDRkM9nb79RTKcAkM7Yaipa15vcSyhsk0LgLkEozloHonXl2+eJu+HlB5yvcJhmx
fC+v+2Gty7ziSbRD7oehvQmxEDYjVILfpHgGBF/q7QKVINPzzqes/ULOlPmZ4uyquPhNDrzRHGHi
qmBwe4XOkBSuraxn1jYxe1xG+/vKzw4Do0mC4inC/m1Op3V7YnqOtvQma4UddnUmYUyqLox2Efkm
aU7DPesu6/0iUrNHaIQqqy5xgr6iVKQ2ZCcWFHSN+Q/93bl2k5ZXVZYMPrl3ZasDku21NWyypH/X
BCZRTz4cYcJ6rEaUR1Ru+7hlufgq2UuP/M06GTz/boA+n3O+nIvUmqg1o2qNbSAoI+EpP9R4jJrC
ZUkrxB0zZIHcluh0Sfl+b24jQBX77SoBcqHcrXS7k/y4h5Kku7DjSz0oYAxNWTQVkVXNFEQZbvJf
gDOMVJc9wZrTqX8f1ax4qUlqAiMjcCx4NjyHMLIpEubykknHqyhWKt1P08rBkgaF2eRRfR+8bzzR
f9BhZWeFHP3BiHwapHGXdElziaYFyoevT062gqZHS5NI2QJQOHFcWMnj8T93UlLV0tuaAXw1jwss
TInCYglSS6i8MMrtl+ItBGg5ikzivTA23cb1EtY7gA10s8IKIMejf9oj5H95DVT6/w/gicec6aaj
ynRvoEroDzb0ngVr9MgZBmL8z9qAms5JlGyzNMX7azyWW3v0noW229L68PgNF8+wDbq5MRWOg89X
HO3BRBYisTfVk9Qnewm/CR6mOzHVj6Un45o8U4cI4mZmmAIkkm7N9zueGxJeaDpq/rYWgdKJs3XC
jOBbViYDPb7bMZen9coViw/Ba9DS6TctyySXwVL+BcAeUZag5alwZMnlpq31ocKYW+dLz4wrTxMo
Sy5Nm5ob71069ZfZoepxLav82wMwA+GEf68mfFCR3n0q47a0aK6QBsai/ZtPMnQNovSoNQmGOK3B
soO2cvW9qFYsz94vygrsjZuya0BH9Rrfk3zkPkuDZU13Kyq09UbwlU5p3s4FZb5W5hbo+bH0mPT2
Payxm+d9zMJailX4n3MedjWnGq/kTFrdPrrREw4Hlr7N/GvHLovP5Cmh8YuBEyCcLlju75Eansav
EL5+LyxUfUoV1IuFhFrhqLRZ1rzippKBYRkwyCuF/spl9yqFCTxa2niGM8P/BLcDAmAoo2ry5LMm
MJEonS+hrYO3IN9758Beu720y4iDOUDcERy82cv1/y5gdbGOsQ+fPQaJHDi+nxp8KAP0e4l2/U1c
3KLjGHClxnJs43LPD+VaDUrd1IrZrcGtSqC3yZ+lhr/UpK7m+NoyAnopymjscdFQrHqy7KB94ADp
jmfvqvxkH8FFgPDxBR7LPUvNTXnl6ea9G3oDGBqB7IVbHrbfoKFDAQvEgHqqcy+HbZImwAahibG0
iPAw3o+cxhMID/EQPv7qOexq0F7cJvJGDEOJZBaN6hsLjXIbXzSd7TrjIrT0kUc57T0joMdbgpDF
09Fdff+oR52+drz6I02NpHjZ3nUkhaSxIPsQAMiYrE7zplHvaLJ/5eIEQstFca+Uu1eCniiCirD4
Wu5ifyPnngSiIjquaMpO8ywjNb2vzendDn4o+9nv+oin9OqdNmQ1wMhBRp/5v6Ur/N66RAt1s9ua
F/JKkOGG1ok3rAZSHDcWWfcaahSoYEz/IIVBy+lAMgtk+Ah6ga1wzAl9K3Z3BMdmvhe5U7+XMcQb
GdHIspHSCrIO4H1GV6akjOf24pUgqwPXDngp25O4/q/ZS5pZoNcIwwaymDdzb8wkxm4Zs243/ta5
S0Mxzqsd6cAZcowzmOne3aDYc4nEL+CkWCu+kU0MgdAxiWWceL02EpMViWiEurhy2nzpqMyaIvY+
eiROJldiLNp7GYXVvsZvCyZuXEfyeXLfu4hwuOE/TwDyi66DRN+ZO7AsZ1jbWJUal2aJkNFrUb7Z
wbNrRp02cpHOpeJX6o1h2RHcQmcnQthgHVAl7aaUyKpEYlwX9ui6ZAGfaPGQsIWxPSGnqfdFYpPq
taM1Ix559NZXSYvDgotfFuWYSXJKDiLunRdqEGs2Syem+Rxo9gcKNhe8CfPcIBHMYhJXphqrPu5x
FUmaIKCFKQbeAht/j4CszjymySBGYOyzybpRSSpPKukCdYCrEflbsmhbcdBo6NMRLf2Hjgen61EG
ZXdlO6MjV2VYoIHjADAEw42W/UpfdTl7cQ+sItzBdatblpTb9Z+WX3bTWTnLYvrBlxUsHJDAoOZW
VNi9ve1k82TxZZpEcD/L5tiZmdT7Enfds/2Qb1nuKwTOkWisIz4IFoNjOZvDjFq2pnBIfjx1k6ke
ilQ8GkrRnMVzQB6AJNHwmeUfa7QeQvG4KzNPn7NUqsbFmX/TEY7WMeBOpBOXMp3mQr6FzgYCtxru
rxrklzmKLeHCbxAdLiab3LzAHJzqYI5VNPvL75bUs9KDScXOFz2vo+7QMxMlShKiMv07FGaOGreJ
F59IpyRqNR93M3d/sNGmDNYc2vAOPZ0LmRhfEeY77jfbRr1ajlV53zaAnlf5rkJdKnMISro1Ekiw
oI83P1gzc78MWu0IfYzafcPb4VeYRS4pNu34N70tv2N5l7YPAbY3kSyNtXgrHmYGPG8hpEeHAXZ+
CLkVWyZEwRrzDwRRT0nL8xtsynl/+WxTOp2ipH/Rymwb5SojzPHd0TMoWk7PmkP5sL/FA1xhGZJ7
mhj4+dXlF91eDbst2EvnAOZ5t9ciMr/aQD3vT4GqpRYbHvsOVz2vEtPTB1dTizAfnBvNkcvbxC21
BwgGKzBSDqkto+ZibfuIroq/DQ2HJqimB2nFxF54RpwaFrJZ8bOooj2PT1ac8ApLXhmQIAm3UflF
QYK38h+/GYoDJ4h3yzyx+vEwj9RKERKzAIeGea00oknPxNb57B5Hxg5OhNZniu4KmNp5eU7IhZ1L
izGo8xRx50VsHz+7PO6llc/9lSmVuLmx1K0mrmT1qDU4wI+OMRV/APvhewEjXfy1bDdG1mpAhefl
FMBy9wsAGiK7QdtEdbiJAvM3pDNmE3mDziIvcK3xjjOasjaIV54Kdlkxrv5+fSgdC2HM4CsyyNTW
7DZ41jWjPyH9MlX+Qia3kZ/xUzUeQESrU7Rtvz61N6Baas3CYZvi8fETeav4VOamJ6B/ZhHx3Ntm
yIpFLS1GHRiisP7Bhdx5RV/UaI7zaVXxNX+4XrWuO/AkuG4N4feH9dU7TAbcqKqjh2mL51Gh2agy
kef/KDNjUHU6KJ3XuMrlX+NyCeNnyAmZu2Iu9oWBZXwq8P6ZjWs9zfcfaLDuuKS7T6DZ1tTSGyAl
ITavLdWAtAD9vLp7HnvYJ3xLTKtdw4lamNK1AbFoJv+eMwx/pASLtRfFO/DtfbwZogeGvzXyZ7Bk
NXAYgtvZe7qcoQCqiNZWgPgjESwKd5Bqr8R8US7ogB9SARbG2Q6wBF8yyv3hSP5Icm34CYUfn0wc
70ehFz+J3ldNlR2NKvdRw5l6PxKlX7aj2pFJPOJb55KqpMug+VXoXiLmlaFpsCDn/sUJjucWWIzB
gCKNBL2XS2uMkNpP9vqeqsR42ZkER28RLEv4B2+xY5fjakRbQtica1kVfsNuwckvUQIW/8LQm0gj
QsjSS5/+TZeDgRtLptqvBCuqSC+hepKnucfPDKU1YxIIq5D5MI0xcFDJRs0P1mk/0DqiJrJdjETE
tg9CoMHj9k63T3yWXp9m6zvWb7hFzfPydAHzDC24+PwWkOWjJFWqEoHaIc76qxGps11/L9YCRMy7
od6It80jH2I9adf4Xi6+/unGwSoepxlg6nB1IbQz+pmP+3vxF4yMu3WORkMzDlizUtbLWkdt6sOc
pRMLprDb76h+QSw++jsgfwA8TsqSCRwFRH9zHUyKlAk0SGvGewb03os6QvQHSLiK+DlX9yko7smQ
b7JRFgZ1+s1b12wdjGXxilrCySMjKhQ8iycdfcTEQJQI30T2vCxKR/g5Y9xmyjpCNMgXbqHLJteF
m+rA6VgdVhb3bT4rLvuW/4ROCJZShpEaq29LasqHRFWi0he0+G4vmLpkrI1/K2itgcB8ugCpcXzq
1aFs7tqkfSI9gvH+mv1GlN7XOTFyrAwkZn4/upoFPX3psThgKn0ELRpvVo8qYnzt68vJ7wGVe4t2
bKW20sC4FOcEYvgXoxwYvhG48lxE+a70ot1WZkc1E/CYH5kMVuyUU/mXJsXZDdSbR+yWjcJHWebo
uReAHQxxFpzrNnXDKaAz9omq+OZC/eg7h4NwFSUVZeb+Q3dqoK+ke/HgPlzemSX0rT9aoonU6QpP
V7G9FYtgjkEnx3HMwKwB5ZIvkzLUjfXyjJMNKyH7nHHbQW+XLtdM7TqyBi3pPgIDD0ZDE4CICjki
E1lw2/v+nj+MiLni+R3EzVaaAomQes7v7dcaYBZ+AczgBAOVyJGzBy2ICoO5O0sA4o4bha8TDNAg
xTgF75RncIj5NtKHAaXMWExACQ0JaPRZ1HKjw5r6SWYRDd6PuQI5r7m46Cbtg9WabR7N0DY6qacO
FRJsNab+SS+xJha9yUoxX+TE0HY5NYGFcfZ3KpUe8h+PLoyjiDgMO4Z+wWvSGS6mRuUGyyxfVeH/
X2UG4TjkHjwz330tAsNnGgeV8lNvxmK/vDtIi779wegrStNXbVQ9yqrJFggpszXdG8eRnFmwJzff
xYbmy/yo//R5BY/qKaXuDMiF10a7D0MOIH3p9A48ZIXBQVTsugyRCrDoe6SF/an53Nsf3kBfx1mf
gVDioxGIqFk2IwEwXB/0fYC0IibH/rFGlqNOQIqhTK3tEycgoF9Kq3tvmmM1d5tYSmL/c14MDFaR
i6TbFtBQ1V1eS7vkZYi2BcT2VD454c1F7IzX4wNrYchFDBRrRV4oRnH6oJUDhCz5h9IKe6rC5nvU
Stt1nSBa9E2BBBhqQMmlXFbiUMcGS/MmOa6lDqmxZxbCaE6KL/iTKCFSzEQskV0skOdGAA9Vc5Xb
2f8Fbr56lxxr1Y+H8LqgLaq4Ku4ndesf0JBTtsBm1BC77Od2yrVHt7DDpToUQKFMtiXnAfUkdMi0
GaAU+IaOLeNw04ptAWu1d8cPY0f4WsluYg3iKwtzd/eqxwhqw3DkTJQYAV84n482ijukjqLIi0XX
10R5fc06rQZQ57viesN4hQkIS8JJfItaw0DxjwOOeiuUsYWjD1Ymux2+jE5D3+q6ZoB+/yjGFVtd
EmPsoGNWlYOUWBPVYBOaBuDJqCkPwnbSFAwAUfAFGY1gRq+KLKyTizexdhyvXlRpWm5Z7z4pmvTN
fz5tYNjS4MJPb1dAsc275egmAmsMl8Jcb2CccxGZV9i8DvKY/T++CjP5ftAadgUiCVwn9L5P7C/n
zM9ADriAIzGMS1Q9wfihZ2YrFuMN1fAh0L6Al4lXH4UcxCtN03w8GdmLxn9oB5J8HI3pTM4SfVCC
KQZVuOsY0iQjZ39YhZAKJPeRpp2xD9V5Wok02NcexbFbE6iocBrGe7Luz05i6W19T/IvBdGafzy1
tBsLA/dnpAoCquvDklh7p5iEVYgpMHgyiRwSNL9JnL/2YAzo5qu8Bt9J/2nFuOhmGND66BD569XT
nih9EelBIEy+ndyzgPC8a/Y0g9j1PomKTEzjPKSEwGdPIxdO1XWGTtPp1QJ8w4NvSW4gbpTf8MGM
PMXgcFFBFEVfTKbflaZcBp1uNl7eIW+gucoJLwVbeuMdsQog99AJBm25V50qxHtP72eoGZhm6EEY
af/jxyo/jAjrP6/ofXYXRhCPEOfrZDiEe/sf5UQUJ/eMoIfvmm/fa4b2gMYGVMP+lYpCpiHFOSfv
maSeiTp8ZPY7PfwBoeLJuA91qcE3rbnRQ8qqdPb6DqZFLkNFjYHJ/bvyA8dK/7sxqqyl+Q1t/g/D
Hxxll5UPkR19rYDHMUobJ/suUOlpAqIAhbqNlVSnY6VKVt4NCxQzG4wNVjsYaQN5dQBRUZEH9/D3
fJfld0Dtj2aavQAfeCCLnQNW0q6CGwFS4feweoHDmlJWnaXnFLZWr40945t67EYyKNmUl6dY5pjR
Rl5EWF+YuuucUE0tfCbabNPpzqdG3EbQiIZCkzDkg8I+/xg0mdZxVta9/vpKQhROuZTu+U+58mBf
UjnZqwcu0Q1FzZJgg3dK5K9Ywph6sKMmxxnboc6j681+Y1hScR3zb0Rk84Mdzak6gVlGGCsqR+ry
1QHsrC+uBNXWgNsV6POOKSpFFqGKDNrrGlnprZF/baN4AOHXxdXvn5PLXs7t9qCeLwlYG+7gwY9z
frrk88FBRUuV9xNDQUWJ0ntEJmr8mcpjQ+5eSzrYmiQhuLExID0aJrFTvgmIl00zT7HwbYjTGUSC
ZWMzxvywGxZ2G1Ksl700Jn9zZDw87YeTWORA3UI0uXg6Z6zH5wn73Cj7WaOa5k+tEJ98Tv1oNHGW
aZiSD/f/U/c9RZpekr1ShwcQ0FE1zzap/ivcUMiekjpxf1KaBC4DxpbDRV2FL9F8vPdc2qZu7/m1
ct8sUxmtJsbtRicJOklUIKvbiM6NlvcA9b0Hchlc8qfeDRIGXMSbNBZDo1xSg9uBr9wD5Ks0sauj
+fuECNeeIbnFZu9jir+ZD44GNJ00x6l+b8S6CovDt0W5ZuR0XtUb/KfPEmiPYSlitmi77W60AyOI
qfxrbhN+HPDFaKDKvczrIPHiP2uzFqNlkdBnPjhpStQnlAuZqR3f2QIthrRObp9sshmDYxhJe+1h
aQEB8VfTq40PBGWFSQvTgKv54F7Tm2rR/0GsPe8icq680j31GWOwmaWtHCD+ND7cbFQR3TkotMjV
2gtwDf/MnracJXVKFBFuX/kP6O09sEjKlYdSaQUCumH9mF/mBb3L4evYbTDTW/VAImdtXWfBAF5m
xsGZm77N7ki3kKB/9Z4TZ0EsOzkpOp2rAWNRzndGtjkGDEVAzeEd9X+uakA0uEv3sn0tABPhdfas
RP80iT1WP9JX5GatK47elgi6bJW9mT1DKyyZ2/WZychXxuveJZbladHiWxUhmWHkbUZzDxqvLRI5
TTescSsEOASJv3XQE0XptS3YbBmXGj2x9AADKU5J5ESBZL5jX1yEXkX9o5NCnxabXO3TTARLzLCU
mlbCF8KomBPzNlolnK3EtLlS6XnQGrqEkaPsQbiTUmeoSvGYHhVwmTSFo2wX/MgaeeUcszkwcG4t
A3fRASfWtyc8Zwfy7WZNvirzvALpYuER43vo0wY5AxH0lJfaCGkU7s2Wfju/weF+J2x0z4/NcgAM
J/WkodzWF39gbMzFCvxDwUMIT9aHmX9DuxaqrkIkpk6+KGuKEgitZQck+b5HDgte+Ilfa1b4tcGI
Ow6ULDaGtnbMJfx0Yq7YKZFQfcMLxvd8nOsQPIMGA1HasfwrtWATo4rSZiKLUuW/Dl/kVzgWxPLw
HIlzMn/q9Za4EOLV7Y1QLLvqLmu0tPusRIsH1pAU9lXiQbeaultHaBAnaVpXmK7IpNp8WuxBYTjM
alC+YtgTTdbEEQmWECOTDjsSAz/PF4CaC/67umOruIlX8zQFsAOb01q6Zy6njPwW2VCgH3ipmO3j
PSHLXfg0tI1FaqA7IYQMMU5eaKpso/TiFVXNll4Ab1TI0aaalTL6O3yaFezmqYR1S7Y4wvNprRPb
9vrvtic4bleygXnRbKflsxgcBMTGnDMc92bmOQXVsLEPP7MXOyqSYH7NyPIEPm13XXtCcG0oNvvt
lev2GPN1qibOnDkY1fG0NCWXlW5uX8/Bs9GLMeXFoGvzwVXCaEuB7saWonkogzR9IExi0Uw9uk1n
k2UYi01l2dmOJ6ypwAeLjT8sKdkx15bFMISszLa/f5AZktssXgQ2Mbip6+f537bYdmnKUovNHitn
a+Ic0DPPVfZU3nO+d4tMP6PeFHCo9t+wFuub3vnhuif/+z3dPL5YhbLqKTWhjVmUCFsXgxWOLMWA
8dpluJwyis9egHIZKlQmyWwtfMRAeB+0jeY4WaknChzEZWXdABe3R07JBtzmNInsz/wmBx+Thj7f
w4wMeTXre1uIOLcfKzFA6GYkBzrhIMfylullalQqbfw4aj6J46/MSX2L8fQ6/PrxzVZMUgsBTgWw
OW7upGPTL3CdJ+ZctKvOcHdcIlLAXv6S7ZahgZqu3ZjSyCu9B1nGZR89GxLDoUDjiXFSA4d1s3Q3
D0Pctk4eiZsIKENoo38B9qESINbAcppREdCTzt64n6dA8l8Q0obGiOZ1LYhLkTwkQ7gHnIF0cW+Y
Xak26/sVpUXQXnVNu8OzFoJw6ATEzkphWPdZlAfKvc3ezYUKwGkDRfKlhWSIsHYWWzNSu3KPVNxV
15hpJJ3+Y1jXIwQlNovFGgZJqtCq2AnPkFSEElxu8A8fOCwYC8Ga2oD2six9taI1sONXPh6SUeBp
K36V41ZwnLCv8w6rGU33We53fxMFxNDBokIJhpy4JyL8/Di5FbP7VU7JsehnBj6D8k7nHfVfulqI
UfLeMLhpURVa1PQ6ItLXf7DIE1biZL4TZ5CYfCqRIitCf/FX69gpfnKqWcMXoaeE2ftygbxOF0eP
NKVVO0zJ3xidcfMfcXJ1vMEsyPPmS4anV4iKVmJu0HtSuK1guZ7lpt0StrXioFHTWngTgeYb6pwg
FlFWYwl6mnOVHAnbg1T96BUXJvyULTIO0ivw2RaRdv+UQnNFgshNVZqk+yAqH63nt2ddV7glCSrR
Xlku4+tjXkY5hkFSiJ0PtsapGq94nlfmaDvILojlLI0AjCYxMuf//0qjvCVY2wwfmGW16gBvhQ8I
tLcu5d8NtOTErTwtrKPrsRJdmnCW48t4KLw21Yx52X+GoG3nIzbWyqcDx/f60TAtIcPQfUAvfxCN
s5EWFPjSPWR6dRQ9A02pBUsgHQ9fCYvos4hJXqU+DnHbnCv8/wstqzYmt3LkFwT7ck8/meoi6HCM
FiH+jHfCnjC9cInpbzBsO4CKOFjkXfxycBiX8OAJDRK4+9RHSsk4OaoMyOukX+p8QOL2q9yXTPhL
7p8rh/AXv4BbJbIdaJdh8QkSWHqVoui2Z3yYU+8P+FeBf4TnBeaCPX0S2RA23A4G3yKGucrbtQpG
4EhfbYqQZxmUcy1FG4eyKdrbIMT9NRitaEa4eJVK7bR5luiT/s+TKAK+41fRgRUamty5cWDmdPrR
Wemi7jPCwxy+6UiQaVhAlk9CGhoKwLNow8YFP+OdiPPKh2kPdo4/SNCnj6y1eFVQLXQPH/Oyl6bb
oSv/XsOsmF41ZDoQBeMQs3nxJ/h/yQ7NJdMZXfzG1lzBkS31LyN4zpF30J0/S+e9hu/kAQEh0dfs
30Yv6z4jRuaAOQ6DykhqF6yN3XaIYRJz72/CuV+OqnULagrIHsnZqCXHOu6uEfBwsz81vyHj8p3O
jQZ00UHScp1hDGkD3q9iznz1HYzvzksN4pRdfFKnvwxRkoiI3ueezHh6RP5Lih89c9uWQXhwMr+2
yD2t+MseHiPpojP62aRd6EPp//jEOlUMEOxv6uJPYJxhb/j4nD0Lq5sMGy7QCCL7V322Rw7fv0TX
O8Vp3iZboBK+wn64i+5YMFg0/hbDRej1oS4EVd9pOkrZCeQEaXYaIfljSDuutN6eQXAPWvaHa3HO
Oi6N38NSE4Vju1ctElTPCJThAXgsKQFr0jRQksjyJn5f3sdGlVFArq/9eeqqHxYHOuivuNz7R8Ku
yiu25inLtcluv4YPbEcgSbkDiqFe6/2UgXvuYBX0/Jyw8BDSvQndOUoVJhPNZQtmyHoiE7naF/LA
yAMO2wGVDg/6t2b08p+xbbYN+Kdxe/rTwJjeGci5eE/H6LjLFhKhPK2O445zimnlJd8D+Wksw30h
LzyQrzdos73tRkXexp/zmJt+XgYdMwuvXdNh3Tx/FZWfeAEXlpw+BnAaoMa7kTdTQasXEsmLUAXU
JiNfOpZs5omtjUZNGEyw00KAfij0NZvpA92BzX53x3dXMJjzz9Mq5Yq6jkpVjXiT2JD3CeImykEb
ttKaQKTtH6HEg670ToUxD+IZfpuL6fiAwGhD25weT95kd8RtBCuUGQRg8G26Yv8JDdbP0QTk/9wK
2NDMEWvdp+OIy3Ls+AoUW4PIe5jK1eAVeKTkmrve2URLcnFIV7LbwhcEDstuaOm8zhh/V2kKIQu4
Z576/oHzlTh6m2S1csJCnnmhOjZwt7F97BEtU51TLu39fuIkidAsI8GSwBpMR9QaRx+cmu+3f+Lb
9ul9YDUeuyNXDLpWqzUvirsclfKIEcSf9l8FX93QOu1YgBU8p3WXqmYl9BM1SWnHcUA1oenBPnG7
PvUIwNvIGPEpKXZhCHnrb1v8D0dqyV/5CBFKMnn8nYaqi8W3T3jvOqhoclHGb6ImtEfTAs3T68se
husuTjFjU7ZtLSwkZ24owlfd5KJiLt9tWl6Os7D41e+JfxOxkaWg+RHkXAJB3P8U82ZJtNKFtT3h
O61rV3cZ+AZGPwxb6vJeZYEAQ2H4MQga36Zh1tACK+RKGXlZyyyrV9BJSOIZOHdnA8pZ2O2tBRno
+ilNctvx90E7/vxHqEGbXKEDXUOdrlf7wTlCsQLxIemFdTo7m6QqyzuI2C17yp3+GchnR1WxJI6g
FiDiM9BHq2fCxjqV89ZP8x7TcgkSGj86BjCPQTDSrjhQbonnYMfiST87lA8rnF2tnsHvqfoU1re8
dkS19ThPCBOWgCNbfL5ZvM1/Sye6XGDbCYOHJMU/RWhpG/KJX/vlDZ6qHsuK6oiP4a4Ycv/amtoy
wmK99YvOzdPWbP2H3GOUhuhPoklPQIiZkon29Q49NOkBYR1O+bvC0Dg79RnJtBrD84MpRmds7BGX
O9/HJSaDOgj9t/Jq3jRQ/A+vNLhK/dw7M67GLujvLUc/ZJWWwA3fr7uHVjYVY+cC1EFv/+500+/V
37jGP/EjN8wvD7gXj7LSvrGAdeWKZhi94DWYBpGW3QJWE0H602DNAxttaIU/9neeZSnyEcI5SrI+
2puOaKMBLgODLj+pL+KBbvwFxJEDAlL07QTctdcIfjpjcqYemZfIqUNBOHkLdNlR0GPZJxBbIrbU
JgK7O0gSTOoDlHGzJ+/r8MeOhXts/2g1HgzAmCVyz77zQ1TrrF18e5q8q4xe+LzLCdHINOHazB8K
nyznL/QpcbOMycdHh4zmNNzWmNF3GzcgDBQVaweL0ouacJ9ctTPvUal0NSHypHDfcQmtLcb7ZDHr
Xanj+HuCDAyVY2u+KiOGhcNNjE587SDZ0es2nM1wZpchMC3RY8hcIsf/UeCy0wTgGEfnGrz9VW51
TrGpl8DUdlbeshHrxGKyP0qQjBliIcK8rZDgjPPHbEEOrhX8t6fI7B1ZOYTCz2BIjw5/I5LS/Q32
t628UCnSwElYcMKdUQjNkEU5yFtBVrWrUK4suqVkAtNzf+7ZVRYRn+WjElmBDHj2Yn7QFD2abIQd
WE0dGE4iQKjPcTzU4FaLNwcotkZclWKBN/PlmM5YJI/+Krfq8rJvrnaG5epN3NxC4BMrG7QuqdXL
E0RS91VTXQVnT2emdaZMUtyzNjpXGNrkNZbz9caKB3ecehlgny33O2n/bvY5UWY+EkCsUuD+c45k
WP8pAmqEUAIXWLkYdgSgE2Yf7jaW2/7mWhFVd01htWT30cTIOj1qocVUWWQk36o5gQuiK+iEpSE5
S5IgVVG9fuRZko+F2vvydasxcrhHQZSGlVTtXPiw+68D//3iENwJLHmXxWxMHM8Eny8wZMltslF3
dZYJN6oRClMGABGrttUYZv3xBjXl6JjyInuwnU3y+Bptqai/PbZuqDGOVmnR5ZQJ6PYMXakEQq3j
nx/j/0go8yQyVcXbn8qMTuAWJEKFPKX07dY9bhvoNFlSBPQrS2HfbvH2FKBVy/4GBZtM18bm9zMI
JRNgsBf71pt8VwdxpIISpOHsqCZjaignEpm2RE4RsG13/BRPC8DROpLC2Mpjmpn5OWrt15efec1e
BXeHRt9Li4GWyMROfWTDX/bWAkjEVmClmf9ISuNts5H0GoGxpbcBM7h6z6RCFtWOFThacxc0F6a6
9xDXJwL6YakMnfkFPpbxPjiugcY5pabB0PPk+aQ9by2YZBdgK5FsA8mLfic1aXGstCvTkWE/Y11w
hXW7i9YQP45eHJWN7NaooahxEDg8jsfSWfdsPMzD9I7d30HTWviE77Cro5yabIlEZ1SuhNYjjcPN
NRZWCLvVNGys+iAFQx33aC1auUsXHht3A7tAw5bZSC1G9ojC9iJ8AadDeL90hJLIE1YKvzW0Y7eR
1mhoDoScerbvun/pmn6YymwfJdNtvLfuxXw6qQM6A2RtThKwKMnYgh8EaIZ37j0bhF9tFj0eCYq4
GfbcZi4Ila9dDcM0njI493cE/uOeM8Z/8E2Lg6417lxYInkzCQLqqPkgfVJAPY2LA4tzEq/BDfwI
+lxOztp6COC5+Er7u+/gpW4Y5TKXEeT4DyiDKO2RAaw8tyrZC/+WsvNAmiWAlz5yVHJetfk4MtRo
yEtqMV201L/dYIWYwqx/7ljICBy2GvulGz+1w9cVY0BkVjrhPO1nyTijGRTTVIvQaduD7glrSyrs
ZczHLEXNxgHj/l5xA8kFueABj4dltC1Pdq7+mb2Ykgy2qsqi2ygPF1p7GlT9bTrfbl6CmxEIQVFG
OYIQQzGqN0eq0gzTEDg3TtAGHnSGSe0eNTeswRicbhj3Ip40dctnjjX5SlFb6k9uCOgGhGRPp2ql
dkmHoIYV7DVHAwpwWnk5L4a7lc+9l9BqUZzcQFGlAtWj97M53pjTly4UhNip0NvH+zuWGmRDZYh0
Con0TlDUFzyWKVuNjy4LEphQFHEQ+mgyMG7NukCcAQnVeqxE5O7gaJyq/y1kKmBmDdjHltKXTJJo
dJL/yOCd/6FcZvajjBL9LA+TtXbSJAv1xP2WilP/+K2viKe6Xl/ALJc4GZ61jmmaenUnZa2muDd7
Xk58Rf+xK6EQcx1n8Zyj4xLEc48iXTE1rh+P9JW5b/4L7d8+toMBabUT8JsYMz44kxLMdKapy5XV
9m5jmq3QvGq5MUtB1oIPZqZhxcV5rstuLMhn/ABes8mlC0CsfpaXim7gNhf1//SRnrKrgkRbkv9q
HnnpIzrXf4TfCOHMROH2kfgT0Q77HRiHHNUPQbrs03hoWSEym+FScQH2tUG7Hl7vAWPzMP47/xbK
BRzLBOyRo6wB1ceMopEqYacNI4UV6oJp9wzyYNSrx0F12PS/f21Ob20QKnn6hmjDnLGXJmBAwayM
TrhCZLyPU16zKEU2PiJIh9NyMtPb9BI7XnzTbIjjwl34mrRCqDRYrXkMBRMfYFzjMo1bPNRDj6br
7OIbuKsYI0hgq3Kz7o33Kd5hXK+ZZrI6wGzH6Sz31ER+0T64MiAHlprStUfaAdXUViEHBP3ZeNt1
MlCKzh1EqTvo9oIR7XWOjTgY54J4eQESaoo2UtlA9soex/LdubCy5uGOmSPS2zZ9bdka383MMWoA
IsTW/FYpwVC+oNa5mBCUm0VqURxD6wKD/37oG383r+B+KJmSrXec5wjgZWxmqDDKVpAMyGcuBO4d
dLFwaZ8BfCZqp6xnuxbzYnwdMbiSdfwao3hTiYi3/YQUnUnxgXyNleoilFtbJ+v1Q1JeNnwhIwxV
q1MdDz7rMBZ9UUMazEnIK4FAHSs5qykWw51eyTwmFfR2YveC5j4KwPcGLfeCt63tqM8yTeWedYwd
4maJYYh9d8Ne5imjV0dVap9+OgDRYenpQeJwRzXLRPvyRazxTb9IIOoAjmTOQDmk/csV094FoTWv
kO+qTpBJVKxAEH6XInLOPocmTw1FXQPtrEz4KNZePtoc55qPNp6YVebFPPGRtJt/qTFssMfPedZj
wV0Gq/7qxg+38UOyXfnYm7t2RUmzjRu9Bb+xPjXhGrObHFOW5pycL7S+HX0N0upDBPuq5OHlsrsy
+xsn2yLKgsw3ynfWoaDkjzAkbtfQtsmaJUcYMmgAPoJkSPFbsrvg8O7gK81K5gkhSl6DOrA6gw/o
AAfHXS+CmhFt5+cllhIe4/jmeKHynxcEEjXB2wyQ6aWSeVpsY2dEHQTS0+Osto/u/UEWj6tg6jGH
o/8CX7WM9wUb4yppRrYlF8Bjx3CNke1nvH/3ETKmv1H+TPCUk+6JjqPz/5CDpMHcvZDQZh+pdb4O
+46RWje3i59iqdwKKYpZfZ21S+olPByb+WODpIeAGovuMmQ6/kp6EcN/yT7HxnXqzZ9VmcWaMy+6
XpOJoAbCE5UT4LOcy+ZqXWnMq6kQpKjUHOqpKtg3pE8klV6EjC6xUx5s4lDoWK5qfLl7ruoOkjCn
slUCqHifmSvKZJwSwkFk8IgvavBdkZc+Ppy9pi6nWOxIjQOwvnAcGYXkCdliiTlMRUKxFCBgPvGO
hyREFlZsiGi40aMYkbvfYPNwcdLQD1th4APh01KyT3EVDHjkrtroItJqqW5hMCc2t9fb+/InsTr5
OOCG+5wxvOoCIjD5V+nzA3TDg5vqYen42uBBWVWPw9Z9EshLClXL7hwaqeHfDpgNqSo1CwzTiYTn
niQkycDBcCJKeobaLy8bkYR0iX0WeooU2+D5wAYkGUAsRwfNhgEsyvAuSDXaEszAav9sdTOHv/yR
25yBxtof8/mToeUyXMVwhdtpGC1a+aDHspfByoY9No+YflJ666LwicsP9UXucTCrMlsCf8yusTLH
fVGn1YKdj9S26eQh/Y0awxwQmPuHIt6euUcLzU2tWZ5SSuFce/cuaMHNAvxO1EiH90TBwzaC8Hv/
6Y85ZcjPc/wYsmUPrsMJOXeqRtaJwfoVAfElcy6IhspvhNoGsNmibgFLG2mYN104EcUVAccA5nGr
seynrhfSFTTWCrA/MNxqKi+hmEzBpqzeg+1znIXvoJDAP2cUtGHbXnuGSFbF/HTbcT42iIOXUIYM
wblYBe6MasVM+0kBkdLftNk9+xoyS4ZQsjJl915niPHs/8y+/zAVJtEYDI1AFYdOzB+OAyZgRAMq
e1dct+y/VRv3XjRiDYKkUycMLPX+U+fuFyECDeTChorACd8MHTaYyYJb1Vb6mGc1We9oD/ZiVNXM
jK+m3hrdItMpH/M1DSNtlmAcqsW5ovao9umfQpl0h5pI0jCaw3gHueEEhd9S/5MbNhpPp4c5ru8s
YzFnaOuzCU5RfVDexihZKJJaZUkzyLzIiVVnuY8R4LAzBeKjwVOXavnUjbOt8COYxyDm5C0CbBSa
4Oai8D7ErBzFEYcdOpkByEbK5l0i6Ea2vZ2ZC8PJ25gQUxFQ/ONz+anN6oHVFA8BgAi4F2mhE+SF
05fCvD6apm95Wr4UIUrffUMCE8s5XFJmyOvLRa807qzgi2kxuiPW5MaiI8Hlc/CbIM3VSKPxZg5U
bO10oqTorVeQjJRBB94P+WUbh1xQFEAnxcmLoZIi2BZ3Bm28Zk/8k594pcz2VLR2KsLEqBbIIjPT
Ed6r9fUg710OACmyiHsdTRDXybi56EIKGZOjVjvXDV9vVJfcSnDL5ENSY09PcmMLB7aYKCx/Wb6S
rEZSI6ymGtlrwI0aXL1w+gvc1z2O/TAdCib2N2O/7DYLiU5S95Zuo23EZmE5UjOggKTgo3mGDRE7
zgoK1Cf+hL0lJKyz2Wi6TH99VmhywBIHzyo1A7EeCwOehogcrr9gWzW0xxrQ7xKEAkzeQHt6cGFT
OSAZMpRHfoxU1ScyKtYVvtmm0Xx7lXukFnGPYDMFKMB8wlLhQy+zWaEWhxlQ4Q+IxocPzKcFReXe
6K2V8oNREoYiFIFgYa1rRXcvJ3MW3BoGNVtL9XT42/fRp5mP6j0nNpPEH9fySXCM4i5Czn/DyUMc
SMk2YR6HX8usYbBarTsnbsFs6Yy+asrFLO3PeGKoEM9rRQVsTrLBdcemIyapDG92Ho7ZYuWaJ8OY
CpwTRoBKB/Us8NIgwCpz3ZZzcFospSO/eZnmmljoFwMhp0aCy6xevIFVjN2RLEQZ/YY6v7DuKwKM
flViDx+KAAg/NIvJ3dnrmFtvund73lgCzVRFx0aYo25VxB3gxqyumYrta/6X9/6I0xYN0qI2/SqZ
IBmSSsXT10sEvFMlzCk4OmzZTR0V7701VElxDTQjkELTVzpbSwLeByD49b9RdQ4wlz7By+rF/+de
1AqXnkss55ZBCl9OjnFPZYEN2D2JWPo8e47FMwVIcA4vjT0pBZG+mN//+wh6SBXm9p/vS8nbsMGr
SvTG/0JHV+chjzhdZ/Y+oreLYP5VQzYSy9Cedi4rWqx6qciwr3v07bzXr54z1WSV27XRBDtZRPF/
ucXLqCjuQhK54LLTe5HR7qnztWau1coqeaZgnxyHewiNelRwZWXEjaT01G7At2N2QmFbrr9youRU
tt5VMI0Pv3GpxHyEoS/sXvYKVjej5MA0u5zWI44oO//v5ZSI93rMopMApE3y3wOzGNKTtjrWfmLK
GIZnMpAl98c0JyDwVftFvpG01SCIG1ord5C1+htXmc3z4A16VSbOAQfXB9JBZbxZWcmYgKTHc168
SepDQ6p9L6IezXm92fmCNFFxtD2RL9K44xn6PD4Tjdx7+5jxqlHoaBo1/f3SIg8/lBe79UyM3hMQ
buupHlJ6U5BDvBK/pbhaU2B6lztZMKPTla10/2ks/1Ibcvvj0oNU/hexa3o/fMRzeDBHv3zb9OCO
R9AThPiam+PZnGutTSWxbJfbKyIoknpbqqpSgLaVuV2srPT3vU5qnA/k0Szk81SnuCCUf0aCwSGy
URG8OHx8RZeLf8xR5sPsYY7fKDEeaIn+LRvhm7cJUuSShC1lLfoK4wSs9xahb+hguAjMp+gYwQDB
KBlAli5PJhxXDqI9s8yXXGf8kE8rVNVvreMY5+9TbtI3OKWqyWe3Nt3A6HArfUqsG56e0t7VyeRK
y/5lLl9XL/lKLToduIUgIH7bQLwNZFlF5VklAqn1BS/JDIArg9s3MI77CPkGpgwYbQwJJv8dKZs5
sqve4vWijEYwfcQmc8lYYrJTDzDX8v6jxAGgpvNvxH7l2ioPjNvKa6/yyvQhlYd7Xei2WaWpfS5b
ZAVXnXiUTDwwBRk9PS3IWcaEgbpoNMNlhZL0DdxAHeUDdE0gtTMv8oOJQfmKG4Dnt908XInbQI7L
kkNw/Gl19LJqLJrrkLBxF+1h1bSw4i3xF0lnNUsOZXjAFrGcm7X/b/kj+TEX0LiOFkiuvqUOiJNM
f/civ6qFEx7x8mDNztWSWZq4goMP3z5HtHheKVBa7poSdfAdV+6TJkQOUYV2LWo4EY5t/wPo2OKd
hsSlZoi0lk6Pb8+YUoqZ11zkCF9WX1ne9XQarCEJM/1h25bu9xwjSTbJtLah2orQPdQfmXHkqlo/
NHVQMJLCFJYWSx3Ef2mdZnPXvITiCv5EQiWrmFNOHmKUrJQXtnU2Sg1n/bYcilaOo033ESQKgB3D
liVlLRNSFS5LqStj95Dd9KJ0J57ABAHWPcDF7aPX3dHOboHlF+tyDTWwYtuGtwVkLtfQ+UOTLdsf
AmH2NFSzMc1X9QGesdH+Ct8suHhdqm2N5ZYpA3oAvgxvakOKksLvmuFL3LFPb58E6mKApSUFfdwR
5Ndr68mPFhw+6dyrICTVn0c2LD08ObPasDCJbuUhxjDjPbmZoEFnrp6xKV9T/8jlciPraRiBUbtW
AGIRVc8cYYpdKB6hhyRPFwMJ4GEmfY6y5Xew9GSems7p6mJMOC6Hb0kk2Jw6b4SUCa5NrW8q/dEm
tp5kY/Gp/2pcY/nQQxogt0qo1QO7P8k14BsF/UHZdI8gTBIu0nAyPcHb2q0aehG8tH62S7nJdiww
R6SJnAMzowWVgpJaG3IgLkUu2F7Ri9LiLK9MTigPNe16S84wuSw4hholaWUcXVuVhzmMkkHoVBvx
DAmx33Rvmmb2OgdnDwep87kOlIJ5HlJTwrnhcE36wgVy+g3HzkpPpqplW6/Sa6qXI/UnB3tG6Hzz
ahaLfV2Im4ruuWeGgkKj3lfpHbIzg7uEy1ZCxG4vP8CsH3QJe/MSMVTY+XXbLEISjEK9Nw7Pwy6R
hXg7naNi3p25jzSiaZlTTQwG/tTS4Fh66Lm9nmrRROhY26rREFCM9BYGNJ8ZjlvMaCfZM5hwVhkC
Ylqn1tpk0NfSKwhaSPTJw6z80BA1zTkR0oo/h2tnfgExSCB3fbHmmeS1duAjOVjGsLot9MUHaGfJ
8VYw52kdbR4fbvpUTL7jSIhz3WxlSUkD47EbltffD4pcrV1w9FxhSCVlTtMc0uxgsFYH/Bu7zCOX
UrdXk+wPI/nwoIYoHXr8sKInp+eYDm//LQ7iX5+zCZFdtm0w/jT6rbkrCPuqWa6C8HJaM12q+jTJ
h1LuqRJbPL+Usq3c+hVivlUiWEgkj4+FEALDbA4zDBbwcXKvejiOt5y2o1J0l/VKfFzkZRvU1xPt
QRcrO/PMVR/XYbg0UCVEd0zfXTUu2/gKeJOw1RMBh58T3ktwBFQkKfTabjx9pctH2UYczF3IwlD/
szMs4TBVFzHZgvKvZig2GzILta4Y2GI9gkJ/9Xl25Q16oIlNyURf5caYsNctv9pn9m+hPhZphMnD
2QfLipRtNQ5e1Dka4cgGiOTPdZbrKWYdh4vK8h0PAn0JU9xe4GT/R2Ojh/wSL9ldy7AD+W+wTDoW
fakp+rBkYJ6CFZ/bD12X05mFzkCbDKZssVJ5seQ9Kjd9agIlMupHWHvIxY4aHB9J+b78IDlZNoKH
0XpT1QfcsxAjVz4tiygOyBYpslkQK/Df7+EZBCs2qFNawRjoKUO4tIfAN5YXy1Tm8Rab84HW/h9y
1agXS5ZSdBUhxw+voR67HlE4JHVcW0W8dM0i+KOxEqs++ElFYojRl5rMh1Y21+ULe0lUzIh5ljoa
9u9UcFYiHQENJfG+XnJ1ATXFbVX8xVsugCnAoFK40EOoG/ofNzRA05IRyR0OA4l6oN3Kfwe3IGr9
HMSpcZIZbBwoU/zQqvDBHq1GeiLESexWCp7VFb+JVGAcEOAFeHzjOq3erTTi1qRjvwRuc6jGJbmS
T/4P4+SsX2r+RUr8wjuI+da+ZsbugO/xRtHTufcYBJ0BnTkID10rzrGBsrT+7DE6KvzRQP0MLwH3
YAMXVreQc/2SXb7pxbEQ/ixOlS+a47BJTWQj4GdRHVOTiI48dsCA9qD3gArg3qkYaLmMZAXpNu2G
Bu2CaYGDQUui9eFfzuyfLGd7Bx/m9kKHxtyaIjOR3p5yYWKrG+mRnf0t07COToDNJ5UpTFGtqgQd
CpHibibb0WhtQnAZXPM3AnYu1UvfHFkKODJ2F8hpU+PPsg8rJk3XxyZwmSOXu+QueO538mmuzQPj
6/hsDo+SmFf6M8382MTcYgj9cbhlrz9yI8nc09Yd1+vV6I89XZxb1+Jftry7IqywwNfvlBPGMQnL
tiKfZLdI+HsBV4vFRBt5rGpyf4qBxrljf0QLTOiz6iEIWy1OGdHJjXQxqXuT/6I7+2XD7g5tdalu
skRo+Bf2EFAfFUzxXiuN6UQHQwEEkWJhsumZQGZi//XPU8C1xUe5p0UTzE+VWjpiYuoegz7OBRZ6
aXLmdE70NpQCS0o+w4UtobX0MoZnK78UDDcFOPdGIZ99JiK3zYnvWuwawMrXG8ipFfe0J2KhnS9o
FcOxAxaPE9f/Y6td51jhmI3nxXiI0G0HTkF1eUZLZeAfRaSdUe+C9+HjbQizoYKGzTFdibKzBAjH
/yzUXl04QiA0ND7zpli4VxJLiP5P9NCQzWD6Lry9sEtzaNSGagb/R+BCbTE9I6K3Fn23zcQnisVh
pbxyKZUl2m2x33dvPxViHNyMtP3f9b0Ciy7ZYuiHoru/YXrATZvznpKINVNIINdoXdkrm1VkEqnl
pUctNiJAJBsg/QX0pYuCvpWsGCTPzp/0g0ia0pen2HFBKgQUT6vWO6SNmfENjI/Svm2Mi/QnlpUZ
bWrGvsPyqrHTfhL8CDmY+6BRFC/zZbJzmS5ITzWmmGFRmUdh+NmF8trTpDVlW2gz3uW06PX2E2PM
JlAheRwKtZlGmZ/zV9SnRA2tX0biJKg7TrRaupv96eFfchDhId3zYau4NjFm802X5ogk2pmDYPF2
fFH52oxsMLHbSz3CKe30K8elHe+TZ3P495mq2C2d1DMc/qkEpl6FvjxD6wECvCR1KHfiPXJiku0W
6pKmDtk2tk08VU9s8mTMrOTtCxTrWYNeCXR22ZQxvuxey7a9q3HLSvof1UK/Fb5h0ruHD0LAmJLq
TUrN53QeBTpHzKP+6JBrGK6l2888BDdBQGhTq4KNI2Do78Exbx36s3sEwqwohQvKnmp34M/AeJFY
GrX8hazKjGtwi9K0gimq6kHWIgalV0o10KEzDjctQS+9jnvN/sEPlgw4LksOgNjFFYfCh+bbYaua
1/IrdJOGrNdjvatFpIxj8Vcz/xh3zdgl7a4acTi6kY4n/RrRxAP9Gaqo/GvisRvyUMGhzEPQnNB4
zvYKHS8xTO3sxA/Oq47qcERLR4lVVo1OmwnVvaiA9K8o/Q0BrhIUo236IH0zXzEzV7mI5W2hABaP
nGFsdxn5gaBzHWt63FfPBSQxVPEFxqtgq99fB8HQIET/SQc3MQuNchZ3LZjF+wMiMwp2WR1Le6r7
ZPD4Qkskg6p0xkUkZtWdhXys/mekmErIT0VHwMV4o9itCarYmL42CKEhMZgTsqjGhpqnxhypCFxE
QChSgzS5ESj2vRv5FdWNxOJ76mCBCyBDqw9KLIY1+hzjrMJnaegGJobz83W96p8ywqCe2fyKaanR
Fzkxh2V+0GrZsC/xRHIhKZO0ZhPvxGyS72aBxt4YEcbiQx5CD7ryEx3E/ciRWweU6/3kqypo3puC
o0891X7mWObTPLvqAnECEnfTBkRY6uzAvU5bYQf4XA3C/DLF8txY/WKYc+ibFcGu1Xaiis+1otQt
HMwZ3dV0laBgvBuTYrZ6d0UfdWS4V2O6WGMmm76Kic21TjeW52edfFAbDiFFi2roefBKC221WRIU
KZweoUjgkNuEGbByA5kdDOlJqiAKVjadZMOWAoFgUhpxN9B8IEXhNgSSP5yROleG6q9uSQcnl1DT
D9ROpnus2xh/TC88u7Jr49OreY8lVdnsvpnuk3kX7yR0Z8cXpF4GhqZZSjSrxi/VVx0qz/F+fWUA
56oTxWsy4nG+1/81bMOUfuOKqmgYtUimRAKlKp9B040LF2TOaABIMZHCoB8lfG2o1wZstcEdS3Fg
+48A/o5+OZHGg8ND7wdK+mbD1d+GmlX5YCrQZV2O6xTTKX5sLy/cmlEA+ONe91XQ+GvnVX3IQ/TL
IUDzss+EqzI/H3yT19VdBTMUyp4i6iRCsFG31Kd0h5RRUd2a0uFIx5LNX4oczygLhC4KnU9CBMTs
A+q+IoByTGXScOEVv46ffS84qSDY0C8Hng0QGBbxNqga7fuGQ4GKsME2R9olCE0HEEQ/7q4lkR42
2eWh4zRBhAqiP1+hYz0m0Fx+ksansFWE3aT3hPZro3odWXedBzUuW/xTdOkm57yOeTxFGV11hC6s
nwfx+WqsbqgBkhVPvWpDqt4HHZnd9f4CScRIo8DyENaBNyeXrPOqyPhIGKzZhDjApKPqth8x3aWe
OzUWLoynW2ZfMWsBHkg8Gt9bozqfa7JlkLH/Gz4AubeF8eY1pZzpwcmMnRKMzlgVA35KAWvZ0cke
QQEGeJl+zj9+oiUV2e8hTSssyk1iUyuxaKMbDOzDXJ9/QKE69OFNSm5o+T6YzaUvtUkKx3FpioUq
kUC8tcwVcemj8QkeKbD7Rz5lmcsbWAjRYucoW3ESHYNB2wOl2kgYhrZjPawgiQ+MXN8lDPhRNCyI
tIRAJ9kpDtFRvsr2hPXxyENm3nkGDcCK2/ltgKyPCjE7KLqjpIHHMJiAqaZRHKy7rVLYpJwblOEN
3s072uF8FwNU/4lG9eQe6ioTzpiQq5nyedGF1lj6T7GhVkE7vZ6foeKRfKEhq4JNfNGziGzgHtvz
1NZwaOBEIpy9txAI5kbIhIct8UAaJ6fDWtgZ3z/7mHR7oRkeSE0UUirmNPJKCs6bFlIq3mQRBVej
YNvJ2jL9xnFLX6CT49PBv5hu8Xz8RzOF7MaZKERS90LRdrOyPmej+J1713GsCyio22WtPYUH+M7A
l2lrpcTjfY+VxrSlmBpfW9kVBw1nF5BnSbPekdga1IPgcVYfnHjRFaPeGAr0HmExB+CIVYJgSYXq
NikJ2a0cxi7L9HZEsNxjar8hoXVGMJzVSqsXnnzmZYODFP0Pq92dSpl4+4F9Y+n6uaCosO7AdSF8
M3eesIyp3Z9Y39LiGy6XpuTfiMxvqP12yZNzud4U6ugouCd2Iqx+LoSn+Zga4qsqNr6ElpMT5NuM
wk5ShTHVYHO3qolzewHne02rJkxFumuhPISa38oFYAe4RFK854a4mYIPiyP56ON6Yupsowyto4Nw
9tSdEhNqBRVdJpw7SQibM/OIIIqtakHd11xlmRAXKb0aXoAKI/TCirLxnT3fJULC3RGfIZ/o+gRl
nviyhsAtLyACFDywOznOBBlkJwsZIRTPsE/2XXl3vtWvt7NJZl/9Yp2S3oR44OdSNL9oNXGjVTQ6
oy15pA7jkMYUidw/h8kdsPKC+TBrDv/zS0UvcYqSUx0jKrHgi8s+Nw6LbgSfheqTGCf+H0NUaqNh
Wp0YnclYoNowK8fg8ZeDQvoh/k1uQx+/UA0tnKo/HV/hAovQbr+CAv2FCg50oDMNW03hY9wxWwK5
qrUBMJF9+E+Ju+1p/cy8oDMngOaePob0ZCDmhIZKWG1jAG0dqd4uMDtuEd52pJEsKqYJ8pWP8lHE
aGwd8cOHDVAznZ9GGVBc691lDysz1yoaWNQ3hUGThAI9MXfuu5MN2cpC8Jf3IAW6smRtxrE4Cwlz
hpAgQt2JgnhMjFViCm6vG7hGB+iPJjtsrWL4rDp+6X31Ud17C8o9g+6L/8GmvcbdVjtcDyjzgSo7
9uqX0az1KUZ4nHd4onZds1srk8tLmXpO+2QlQk7HyLfj4Hbz1KSyGcbjxID4fNa9VTcDV49m1dpP
nWu7mrlErE8U9jK9m89yACX5P6xQGfOYbphZiWdkTQRbTSdTSn8eFZxiDqSjUEqpnoPV439zofVO
4AJWZ5XnrDAnsW+PiV6MT/3tnL1HnIJZUwBdh0qs3FBy7EHn1I7Du2vftwQaFgRTPqk9sSXQKVYl
MzHe1M0jAuCdHcvL8SgMI/qecENQ59naaZjuy5+s5BR+Qpo84cVdPLY9Y/bBsqYEiV9Xx+BIGE4v
k0TtQKkMr2Ox/bDqHyFVhzPX2E5Ccdfp/WxfRi+Fohi09cjqpuxETgJ4PtRjitsT1e8UbHfjKHMP
6FpOOrE++vUjnJjTRE6O8mW5IYFobVe/rlOu/7oShubpG7Yp6gKh8isFKrMXE3Ru9MrfmvGBdDCX
7IzthqknHsSrkEOzlaqd51cOSo6N6h8o3OgV0NpNG6r3cq00FXRwj/lzlQu0/qcMdmVxJKGo9nDx
jpWtCtDvPpvC1pgFqwQejGJ3zFEPpLmXlDWoInHB/Awd4Vfg8vKYkbQsPVidpXngls/OrPEyQ49o
ohHyn8reA42fDkc0L7McaA1z4YTLBICDMv5SJZWZGAVHyZPwVGVWmjHpv7Tt10Ft2AwChIOAqgkG
JNYWCDpEuOuByGX1m5YDhH2T2wX36vQG/cTzxoNJ/SGXvqaL8h+7LQJtgkKL+y7C6x30QWk6fMHG
wl2LFvMqIEV6vxIVstCIneKBQ5ewQsFPBxim/c1j2R3pwVDNypzOTkuB1hPxi0mOqOUksxzOcl9Q
oVZ/LsFOSttgfoUNvxMlbcniCD01cIkYsDTiRLQEQqOjwZAwjMnSbPJdigcQtDu1DY9J5+PPUH98
fa0hEx99jnfbXLYfD4X1Z0gGXwgGrK/l9bXMTHwP+jGdoUCmDe5E7QDu3i+nWDycTlHJsjU6gUN5
q80IKY6XFyuxq6VT93TzCWATohw8l/sbZi+GuEqAQuzuvx0OJEtPUPV3xa4gJ4T6GEaVxV+1mkX+
w7XyGvY0YdSrs+74+4gMg7Nug54+W64IoAjqK9XEQFgvtgMPIy+b1iRVJiubzVI39QVk3uNwmhkj
Ex0JgBxbx47EG/nLxDM2CwZZp959kkxqWrk0xSQpPGXIhgnYD513keapB5zcqCBkdpd1Kez3H9r1
Ldw88SOtL6T0JKCi8M9QjsTfbvdALAjm0tHpthZJXNtfAb8FNCs5TK6sWmVFu39fAadEeT7bg81O
Np39GrUc76pFmzth1UU6L69dUUKTuxEOApiZG+euYpIbV7SIOZrfI/2W+x1AvnkAQSOYOqpDhmCi
ElRdRoBSrOYdUzrMtiuWEEzgxc6ovEgkUZv7M+LVi56rC5XY3STz1AsbvjTOzXOBhn7aJ9OPakfE
lSxwtEZ5mKWyGNhNCcGJo5NLDan1Cx74ViljuRedUr2uQ4w7z+BASHusy2rT8GnOXQEQfWk+Yoo/
jY7dH7vu7W5+mA3sMfpmAXKQ9diuZh/v2ZTkQPKFepDoiUHczQPaolx8m5oX0iK9Jd0MGINVksYW
SXy/6mPFfhMgwLqU8D/YHnkGShPqgevlNgFv0yUKvDGBDX1z8DgKwS0y0fCdYaDNI67zhN8Ge/XG
BwwaTLq8gndFsqCZZMdbHycOCasAmP0+ypz52ZBldVvFZYqqtq7NtJcP1Q8fNdzsA13d478iJwPv
iydVvrLAh00mJ/p94INLER65IRRb6TBsILy6W+I4x7f6TYPCH1uMntEqZ7EHXYZ9tvHIldC2MyJ9
bubgQPMtcG9XRn05e+V2EPLFzzGp7r/An7wQWtBGbasFbseFyel7Ii2oAAjRTFK+I51PbaD9BBsT
VQ5Yv/lPMX6g/TJW6hErukhtbkm9pq9U7ENIzVeIm2yfZ/cu9hWCNNQwu3qIT7/VTEL4jZM88yr3
De2k3VZeZuDMkFys4JmadPtOGwKo/Q0H6n+nvGhUzGHa+nESNvwyHLA9aaHCj3arMd/e+lYHw/Q7
ALTcZX9TkPox7ke6PVqCPvqwrhNUQPIwx2VPgSfZpvt+bry4YxYb6T15vS1Tpdp84deC+jZ6s0NQ
MTuGRLHJWch0LY1IdkhAcDZvjn0kzUFA9qVZPz7BpVYajxYnEJP9Rt71j8WJhnatbXA480g7Qjd0
jeancw3/68TnkNY7n03/2s6sUrXGIKXC74y45qFq0IUHqwoJgy+PIxz5cmmfm2n5n18eEh3ojKBC
q3qK0/XRGwh7VwSfVY/sKKH9Yi3/SFQpzk6MlNfhXlpwuTAkv7XB93yLSDR03+rnHdYxUOmAsF8N
syVuS4SdXdvwUymCYFx5xewRVaziMnKNKDkp5Zw7T7phR5/JEw+xr32j0Qa2DqUPgMgyCFBGh/6l
t/KMgkUamvVif0ul2gcwSUfbW1oNHGDGjqxOjOlZxoePniBt5BLm2lrMoyBC2czm/BoizvyQtyig
YUXWcC7Cjl7En9sprUw7RHxHsu6soSpUHKrSPr5XXGfIHDAEXePOIVe5wDQOt8Rjmw3CyI1xwp6k
31NIhcVosplwxAAcnqzvkJF71YZqzQzlSYKbEx8aFfNA8Ssu+pBrgJLnbCFjqnHux+nEfULZPsMm
hTvdOOeOxdBSVByjrUYfXUlKhRKS1iRniYzgysVc5D9rc57/fM7aRZcqj5111dMzUBMGBYYdD2fO
a1vjZ2awEjrVQV+vLgliDnCUkUm6eigusUKdjsUuVRVU80zkLVFDAhiSxDtjP2LvBYIY2n8ffCTE
1MSCVCXRtu7047V3ZjvhJyEDCAeRMgGXo42YmQ66jcRa3O4QPq+oRL3E0TPtQC+fnzcEnn6YHyVM
OVf7MVHXebVgZ/M3pDHoGCy8zbRTI/4k3PaV0dI5Sx3gC04rn0uZZvbiaDK869RIeztkhgazFI2h
hTQL7BYOf6B7G3PvxuZjZ3pkQHtxCAbfVKzKKccIpFyLUlQQaWLZvHoN/Nv7mlHTMzDUhq6WH25C
WQ+vTWm7k/kxU8Z2LzFbsVsQRyvmj/WMNnQ7OJX6IO7MjX+Csd27OIad1g7UB8C83YnuBOGqaE1H
wEsgfUT/oKztvWgFLPfLu7KaSDz5LhXE2ugljwH8KLVmiOHPNpQOhvEvFPP0J/Bz+1a3gTbfBPiL
LTaSJz4J9hDp0euqSjmgypGwwOCgyQqVnWGeLpUwigFFkHb5FepdwYg1QkrIcIISlmh4ftM2Ug9T
U+iF84jpbEcAG3F2J3SaEO4Lj5rjXEN5qfklIQwLC0Y+999JVS3cuEurJjJTyEXvHg7KqjxtALgI
tEuUutZh2R9xR1HEoeaWpRw6s7N3h/ixkWSPQMtMKcAZqJ276YZSHW5iRBJ0+J492Gm2YO69c3dU
XiHIkNo+pQDlcCf9R5qPf2/diaKsHWbU2zVYK+VGio0dpSW3I3SyBiQQ/uCdUkdb7pw4HgUkc/SJ
9VdxiKwowFKsFwLfyNPvba7sji92VGJWgm2VHsn2XjeH+pvzdm7Dv6lEvYwccf8xqYfLylQJ3wJg
mKiZVAxJWS7dC+HkYZBa7l8yKpVTFviVCJZKB5rN7fnbJXTNHmNcax0seNRUP0VsxdZVkODgtNkD
Y1RoImI1ta/eyIZUB+CUP2TA/z+RRZ9sAWojFAffOeQcL8oj/NIui45JGtVm04uotiC0rWjDDtJU
6S3ux2YBDHKlox7H4qabmucdfxfwucaz2P3kqfchJu2gI5bXUO8xzcx2UkueCSSpoX/JqLx1k5RY
ANVNqYF3uUYg4ks5fGu4G0iDCVdpmlkx4yJHPvOBV76lXPLhcN6CD0Q3xzYw4ZJ/xswuK5imePbm
F9ncBISOxOYmn+LdCUoQCxHTxhJkCHhc5af6C4X0h5+GcscLMikA/FteteCN2wboCel+CkECEnd+
2LSp/NWKIGyIe9PyiYI+nm7dK82TX7Okbit9WOmsT0Uh1Qvkzw7+vRrhf/UghoVVg797IgO5qAzC
x+IQq4kDIzxa8f49SXXV9cZg/vxQmB7y1LrEbiiYDJC2Gem+nbqaSftjArqxxZIh4EACKFoEPRWR
ar0vhbYE+BddGwCNkQ1OZl9B8Wlgz+f5U3E/HrsxT6RqPvrOURstAMQ4rT8w76t2xww4tivhMax2
aq2mm4K91ZJ+DYMpT5A2bk5Sr89I43NfvkP9mD0056JTVUO0K7d+/Xwo3HhzTPDTBmCPZqFCEDew
OFg6k705PAb8R2nIpZcbvhC/hecQAmzpYqOu2W2DtN0Dj+rmnj0S/DkugZlXTU8/53YlAqCS0zt8
eUEbP1VE2e2B67Ytid3zLgL1sAvqkZndQ0TReVVIX5+ApNnOBmNkI7GEMJ6cVi6AD2LdQ9lty2dW
gY7d7rDFAgtZbAokPXUXdF40o+V5UA6v/GJdzcHu3A3tcTKGKcJ4+HmsQzxh/5duXZ0R1+617kIQ
iYhdhydKSM4WRqv22c0KT5/mbVchANP4vqZPjLu8/5ScAvQqgf7GXodn5yVvyyJDNxBta8wT2DBM
DTSLLlYhWkEFql2rghHElpr/9kx6Ym4z7LJUUHZ48hq/VT4tD4gYKFvybzf1GUIucF81BA++oNSp
P7aH9sop0LeK/lPgtWdEecVs7XI9S/Vi5aO79/QTHCSIgy0TdHFE6mkuR9k8LsIbWMZeoukLmRjI
ACX4AEQYrgtMh/uozUgMGpUNkmOVDZMXjY7QI6xjejp8haoJdxTfKOZU3QzQpe+Ts+CeF8AI/anN
3Z89pdw/jrNIZ0qaRWcDqhykN2oAOdvlJPiNPFrUAWDC3eWP7hurQsehCg8SrQV8I8Ks+nnmZGwC
0zjwCjD/Hi+0dbREj01LV76VaqRHoQmx7ZwCTzS4kDwdBgx8YhWVmR1at03dUV5HvNYVFTl1928O
8EjovUO7iVTFF960ou23Y+EAoeFHQqBpLSzUk1oCSCN0C8DufXf9goanxgVyd5NDv3hirALrgww0
JEWCithHNlRU5kLDtb0tGgUxCzNoUR7C87uR5KI4Pl+/YvEQrjNG2xoUkMKK5iNqhHw0pLhs2jAr
LcqFfSlk5TKViUwENf1d6zdEFL/zvkIKWiX76NwftJfukuP2yyQwQYDOOoXap1yw15SnuPULGSde
jD/IX/Z9HW/wAhFpG3yiRQmVnU2pd/d/HPJt/elUbmijLiuCt8QNqNSdBJT/8hKG4B8sI0dtd9Ng
MTYFGVWe2MW6CxMT5a2fZxYKrJVCwyJ3DMzIYbvOJcUFgC2V20wAM09GFasxDIT4jwkIqIAGQghy
tyrSnJ5hVVZnVYfML3mlT+dZKKA8V8BP8oQfCPk99qr+1G8heR/vHtzOvnw8nNquKFscLv0UJPsm
+ip3n7rzhPzzDpF8S+r4dPY1deg+OVLKrXo2QSgpRXcqHAkCiMx0NYyBana3RXhyXP2pudb2uQWH
s0oxWhA3YxoHaYr0SN0HjlfKeRCn2uReH+oee1utcXo8/p71VFLRkjPxPEjTiTgM5XtbYS+79Thr
uinIpYCeKpypNczRY+ClZOihgko1gwT8d45yljrFoXOASqHdt+HL51Bag8lSYLHOK/cA5byAX6e8
o8bELB9BX+sGaA1uWKo4cOx3CvfLWCwLeqFUaV3KiZ3AI9Wjgi2Hkftkmfop5QXyK2i0CJ7/q+Vp
cuIhHQXxm9A4+AlMnAkCXn2Czr1R1D3RlICYy0EbvNFZX9VkcPiIIpGP2zku3R1Jold3Xukr6Cwf
oiLB5O0t3M9Gp0SOYfgd6kI9294QOVpbtKuIDo+/Yz3+A92pmapqsimqsW8KTUdhVp1lWH3BpcDa
ptcUFKJPtH5WyZDdi343qRMcLZWYAp9L4fFxWpaCTTpnZqjVHsHTPvLpuNwgHufunqQmy8Rr/uho
/40LSMgyLIuJexCxwd4Ytxs26bzIAXJrOqgIKbjfJPsZQTc2NTe2mVir+mKhM3lS03QtV85YrCRQ
ahIN4C5Ag1I2dvVy8ET7jy5F9OudzSHDYuCZTsnRG7IWyaKVsJz7CJEEeGZFI6bWbpN7TaSFXe1g
Uy3x3gHTXbb5lPUf/oen450+0AIADXPFdAfeCPrasa6kU8MsfOoqwCHkfYHfrRg5kIoYsLvzxE8p
wYIYjdjV0ALXZ6RNGO7H2fplyLVR0CFOOrpQF5B6r5cOmHBaHqai2hIMPA3gNxJlshEpG5i3xQUB
cH82e6jV9pWbNzlMI8LKRdAmcNgrf5+9O60elBLmwUAPQKdWfft8rx5YG6HETRC9gDnk8h1rl3O0
ahKvoGCyuBVeXK9UhQyxufXwu35EYJqTS0c71BYjk9DDE3OfB3tdFvgGnbhLEIq8xcBTpzUuo/Ea
RIuapl62Rl02B3iuIQCXUv6CEh/uzCct0Cd4b/OZ7Y/v5h4Hf67GKgdV00O9e3/2tXoPh3d6xWV6
+j1zlvyuiThdn8KNS3UNZvmsFPUYOKmBZ0mU8w8FBR125yWsxpeBA7jpP49xSV+3P6qdld9V6ssj
Fw9eu5eNly11LXB457+5ChgShFsbz16lgENobslki3DpdwLwjrWt1bpNGUz5lxVQ1dFPP5BQT+Le
g/7OlxiupevkH7N5y+QLqucJAzsHL3jDb/0MI+Wkx47jC8P/z5yPhkb32uFhxhtK3qTaINuIOpJi
0WQYEhsEbgdW9YibqjhI3zx6ICfHpuNgGOKTMk4pR2lmiDBhEO4doFn0XHT+zrLorfCF2tleCjKy
U+GfJa4TnQL6uLx7E6FR+UPGEFoS0N62K6p2j/wuxwHQdnyOTtttc/QWUJbra+ZrMvPUde/urnUX
kAmffemMr0XwXu+O3wo3hB+0OjdNRtu4z74HvUhgz+npCY6dYiYTBu/zrXnJvs0tCYrBwaxfPtSY
tYQ89QyfG+W5L+Ijo8x3ZSxmVHLUx63SAQ1mqipAFb3Tw0KVogWQTjSSW5s/XxJH9fNi9suvKaBR
eKVP5PQ1OIMKTUfTiWyjT5MOGZfja1g2tzynm2N864nIv4spRORAySunRW7sPh7fPuVAN+XJbxVN
XOihN3lFbo1Myxk7grDcyR8oF1KEue9pKle8t0m+1aZ+ol7se21U+ILnQqnX3EP6JsvB3IbXLF14
b4lVHWdUV+rNSMyloTVtmrAs4LCy+ZIUXehOtASHkJUlPP2W8HnGfrEgk2BnapaozvosUEw9luj1
zX+/CnjqQ9WCECy96lBmZ0iqzIuKEW1hCQolBJ7aDMokVGOpGtsAL22oDvg5BrDH/ZE/O7o4Tdh8
8uFwlPRQhb4J42SptqViOgYHaUOeQe69bo9S7GdMg9adSELJzXLeQhreOjdodJruulbXTl4680Uf
U1slWLuqGXIbbXRD7OqolhG18q/mjOEl8D8ikmgOnDCQNQKWtImNbh9mUB+RepWXDJhes6EQ+YMU
ePMqdFXZ+UxhSi5MM+dMnXzSRvASOiEl/EDR4+THU7OH6a/uYn4XunUMYnxvM0oxD2Hca2jOHjE6
5IVDaeZmyuyhE7OoXSOyIjb/i9i5V55K/cZJzU+15E9Ggt46drHONk/5n87AjmFaLa6DLuHVCjxV
oA4EfzPF+QRHiyDmek+dvhMyQD/wfv9I1J0y87HbHMWIyOMhS3bH9RySE8OAnMF9rs3Kl7O+dj2V
19B6jFavVcG9p7lG4OYdlf2owsh66h75eyfhDNAqiLd/yNccqEamODwWThNdrhPrM3CjXY2563dv
a3uiZLXBeH4NVzC0ChdDBeVMZ6EqNiFwnLU4TUfRojc7zqKHyExEQAINzQCwAWsK40H8eTR51sue
WQstsNlbbMj0tqjPdW9+1GvXpyRIbA0Rri160INB0+CpQzq6tS4GjCm1FLvDtXHHwYQ6/6cClqPJ
YQf8EWCyHMPDeKbXDuZQLwHQ9FuONHRpbiPN9pW+QkvNr3sEk3KLKUiXHsYnNmQGrn/RhBSE9TrP
kW6TuuVo+Jb2oP04Q0gr38Kgh3umD1AaDlG9Wi+gRp/IyAjQGzdVTPechROn1ZDCvv9egtFmiXse
Jcoa2DLoCJHKnCsU8R344RZWtsyhiaRdZNRzik3o+DJ+vhKm1dXoDpEJG17v/fFQXmNagSo1hvTc
Vsaf3EtK09Rpijnrn5UwqCHiY6HMqbg5sFonMQmImzuc1g3lmyJ9ZlI80eIJvk9pr5CT3BGamnDM
c4WhQfMIytg4JjDO8Gq/pcceHyU8rvDu8rh73r2h/r6BlaMENNNeQb0iAFneoBisBEgy5hZIo5tD
Kpy3VUifEkWa9p1RcjW0qCpFqwhbvvkVOAoxKAeGMW1Nx18HYOn/mStg39NKt0cXZOvDC2+9eIsz
mfb7CRFgfEaYkU7+JY3ey5zhW4BfqTHDIwKJ+k9b7jXIegddvDMQJk6pPZZRikFxX/PRV9QagBJz
+QoXPW3HIXWHjwNruaEdDWLUbYPMdHV5UdDQmOE+XS4dorWONZuw0GiLWSp+1VBwytQIIvDH+AGT
hxGvul98eIxBU+SE1ZjFPUBQbB4Bf8UtK2efmNjeaXUZIFpyTVZTWnHc7dOvFq5DqSNH74az4lsC
BGf3xFipXIxAiO4PGKYmg0NZui/WWitDc5rAYw4Z8znZBUJWDOKclv4Q+XAfpzZZ0ioEjrdLHFZ+
xpgZReFHKxyDPmmXvLfyNNoVE6u2MuzC6zbYk4Z/o6gxwRSfqO/aLgKOvgvx5VQ3OHhdACJaaT0V
Hucs/MX6USy4TTe4JhDUSgTX6uzVFF9Sdy97ro4xxKsPWSWAI/WwmgS5oC9qjhBEr4H27gbGZFh6
8v619QvcuwkYEjR8zJQSlZ813G7kUNLkK8/7VeByAk8GNQObM//P28bTqIpkqdh3hCfw/TvSdQ9E
aLxcV/pIFVF+q8qTKbuGfwqyMrXymPzNjkfdgQen2tiuW5RXhOZH6z6ayGGcw1GBrv85IPfeYuHJ
FntTBr55e/HXti++8/kbpbl8Owsik/2n4wRwwQliepFR2kxzaIp5uO0N/BfZjE79/2B6BVx8woeZ
JThQOoIJqTxz+fj7GfIuUvDaJKdRkoMioJcU+iqHEnaaxnt1ml3HmD/o64JmprVLe1aIHsIZ0Ls9
lV57/Z5wBICzCIdSYt9uO+7rwFuI/sCQJWWADsrlHE5NLpbyXRC6F9eKGxE1a9oy+nbxjkn27jl3
eB7H1ffmU9nclRg+znH7UmIagce1UcPZUJP3rsiI0NGY61w5LEtpcjbqnZbocJHYNiyjMSVhiVDV
PktxuGct7kffR0e4yPTgnPSZgBBv0GSXj7HrJkmZdV7lpwh5V4+cRKAB/kkF31rXoSObRKE6i2MU
ltuMRMdMjIlvIg797qVRABCAnijaryHjx6QfJAFT6BIlZdhbFokUdJyy+uCdtjUwyri4h1xzy+ry
MdRLYKi2m+b51gIndDO1TpYNRIQEasNkVd/XT/SgEe399grke5EhbC1l3RxFjQtvLO6k9Re9zmxy
cRaemiOgyDeM+yAegNSg//9HpEvNixjt0YKclaGmxoA0uItPY1jM8jnqoZGs+VYE/1sD3nZx+TJA
32FUvS6cfTw/+Qp7HYaHDMRzvnNgqxIO5Hl1pd/CvY5nbNMv06qhi1kZS/8gSsIE7Y5K87axv42S
OmZF+M+QDYahCVG0OICb8Cj0yxP7XVe+B6ffz+X0rlw+tZ7HaZe0SR8q6M5BO0V803e8rTamNUZI
DPLN14v9NE5Q9RHO2JQz8VyqhFtR33ucaSNgxmbV06FjBFFM2o5g5y5r+Xtr5k69e5s0KZuNZMto
ygn7PXFCmjNwYnqI4IGPazEAMpBwNhelui9tkZ3iRFbjnxont91zMx24Y6m43pONV+29A40lGY5K
N1Ep6R+3usPrFyuS3cKhIXQRiZr6K1CZ09mzyAM2QlIzPn1Egb37MUZ7WIxoiI7D2vEmiu0l6v6a
fqCN3saGNMqtjxjZalES4DytTob6kO0NLyIb+8TKVoEy1VwibXMAUSjSc3EgT2AK59xmOAKIZ7xk
2lO8mp4wWguUNIBgXrENqKZs6cTFBBQ7SPoR1Bcgg5ix4JW8XN3pn8v/luGyo/dFFDkHA+4YuG0g
bz994bU0juyCQXssV/BZhU2xLCqFJbZEtcakqweVZ7/L9LEkdjJZagOtXrLtbfKjmZoAhG0kAXgR
Hjz9KoFUFlGCjogMUmNEZ1B+GHXu+DcdQxNxn22tgpacvO3J9TMnnfZIeSEhzaZYctCMs+Gd7lpO
obFx1/f1EsnwriC0E60z3xwDlpODzQp/E1sfVw8TQe2ZmlTrs4WnHyMdeFvxeRb4lZZV3M1BhvwA
uIDbZSjY5CYzRuERe2lRsKOzoYMJ4evCRPMfqsopDt3WeK+Kbt97OlJPWnDWC+7kqaKb0oMsFECY
WWdDCvs3g+vav8qPSUNEpW2QPcYfpEBOIfg863EcsK7hNHlrlEStyqI5XTQeL0Z9BzfDX1aZQ5OZ
jlNrx9DewrAH7ZcweExpr9broIFLxVIpB2MJMZ0IYdgCnF7ovK9M/ffynNHoB3Or1un6VgdmYked
HNfODBNoUTHnWyGNpwBd1AgYdn11MoJY5zFIzQGy6HbwyAofQq3ZUOc67VVibxoqmJOc/dEDy/Sn
7igkfmlUtwQRUBjlIoVTqo2ipWU+GZSBX1mFx6zwwJep+AimbaMzbzOSaS87kUOHM0EsGqRl5WUZ
yRP/0ZDLRE5NDaLYmDzPvNfGW3H1he53iGzErfZKNoOqBSOo0rEPmyE8Nu04bTgMr/iVqH/Yg93d
cgwVZYfZoyLMXFKABUXlFov8+8enEbYxh4rrACiB3krE781Fpi/n6G/4N3ZJMu4Ub9yfM5OvuvUB
FqshIspTobpjJF7hFkToL2+EkGsZHETneycaNK26vLGrO5W7sYty50iC6HfpC8Tsln0xG5Pufu31
JagKdZZ68G4abhJefcqZuCXasfz9Ccvffw8sbjV97o2+6122xeV/a66iYeLF+39rwKaib0lStQlv
60undAwEnSEiFQagpXZs55nrI3bhM7/1kAjGSHIBvUrIi3rFygZoDVc1rUQtWcm3oiKED3NlHWgY
kd/hurxBWXbnzRmQrSCdkWttFcn+DLT5V6soh6SGwyiyBFODTfri6qfdcuJwzU0Z6M4B+eEICmms
PlFsfAhdYY5DPeN7aDxf3yavv6GD1qOqj9ADCN/7jS/pPZK0crlScoe/J4WGCcpgHtcw4orxYA0y
+bXij51U1Uqd3K9s/+F5I3eaMvm824hTZVr1tXhKevaEuUuggYw4n+uYhj8oMO1sjkWnV6js7TDz
l49FJJ8ML4lqCAZYDA7+ATRCev1bZChe3AyKO8kX/DTeQVhf7nMC/qeOr/Fjrl9o5WiBW1J1bUS6
9oMJmyxJtOaAhDLhhuuTUqQZAPq5sRfGpePPT9vGu+00EjAP3HCWVoi5GrSRWLXDEksTHbA14JLg
BzaEWGshSsnUv02mIM8T9pmSSvkd5i7hgO1HAiOBq/0d1OIgct9a2h91bpZ3o9Epug6F2XgUKu5R
YvOkH/TDbIRKhBTDlKZD3VyPzTyHXczG7AJtZ/PsFgUzg+i1kcpkN4Ar7miA+HHN+kTmcl6nOFlF
3qot90Nu+SlGy9Lfb0bHC6Ih9Qlzv/DL306oF+ASTBGsP8mNEvoKAGotvAscmd+jBbzlT+PQDJMP
MyOWLw84YjJc58ERPbAt/XfGo7KvPQavfObBz3zAzbks2IOrVf2vl8YBqgC8k3BPPF9Kqc51HVyT
ufg7td+X+isRdGZx7BGAkDwmx8oTqj5U3F0iQkZUMN6n9TLgRN1onCKiYDX33ypj1iXfw3iEUxh6
IHMdE1ofhl/PpsQcLTrZaadglU2D0blrkG6QAPJTxS0MDDbLfRtOfJKzUkSvE6Sz3kIG3nIKrQLT
zA9KoqeOhUnUEN3QRLltDga39lXFn57pSb9el4hEfkjOHykCGjwb9rzMYSPcq3KCK6jsP2YLlk9R
x1GtzrKS7FUB9g+iWQhFBg3m0OVay5Reh7XCPNwtBm2/8rg29ctJOZ/2IZxzBRyHs2kxPBkgXgBS
QEfRLsDVU8UusU1S7HB6XOMmhROgy//m1oOs7EN1Q78irCh9ft/kn/XH8CtqJroK6y0geyr5DEpn
iSYKOvstTpnORthvYPSnYzoeOgbBlWfpGz2+TNqAeWoLxAUMhH7N8ZJE6eoodaS+QeejFIyqP/oK
C9E11S90/RPzfxQOhV29JgrC8tiA82FVQpvbRY18DA0i0sl+5yXbuzb1RJcdjVHkZJinXH5eZ3Ki
slJ6JZ9OEJ//Et1koet7QiwtljMglbbCHYOELOorvJw7/h+E5uaaIffZHBbiGLZp0Kvm/Seaqcp2
VxklRJEdcbmLhfxwBrSnOaP6jv6+JzO6/MtuO9im1rQhuT1/wO4Yw5fZYEcKhDVWefLPlCRrdXWz
DOQqTI63ehyIABC0l87EY+ijS8oCyEAz/J6J/015qGLobSX38n4Pf4jS5PfYPs9j71QwA45f283c
BZapt1YrL6EhXGXq93KfIqZ59CwpP/awZucD3U/VZT4vz+nzWUn5e03jRSluaCupldemEzasbrMb
Rw9+l9o2QyW1n86I4ymRVc7i1vzIkLKuT7wTsmfUTs0MUJdCTypG05hG74DkGgvLb6KUfvHFEqla
YBwuzhJgVFuVRoGNLeKhxcpwtSC8lHlCTMHiqulb7AlW3H+CVcGCFbHaDuKxJJed1oKdQiVSVQpe
bAkaT9unnQc9C1J+oC7Y77qnCme9DhV3ySdMGGGuTK31v1WIjLWpsNM62Z/aOTOpgY1AVz4wYmSb
rUukdvNOrYqleCSq4Ns3oO4h3hDrLuulwP+z3w6zUo1at3ZuFLn7YT42L/CLLM60pGWCWxJ2MkZm
8JsFBIqZEovVlPVQqupJmc901zfXyQl3r/XJ+1kxPsDXhjfTo5PDavys+WkOoqBCUqHrv2QSSHz7
I1WyazfaTQlXSbcl2uiqpqCZutEq+IHzt1FUXvnyB+UsWk65kj1TF97VYL3nTtfBB89Sff+imLCh
P+jQA5ZQIDzBijeIX6bPAdeCz+dUZoh/f3ZZ2FT1gd6sieCZy1f0CoGFn6teJdxmBEZGK76br6/m
rk+q7Qixhsp6rLUqGgX1oSjRWbREfImf3jwPZQIEqoGv1L0Rrzf8kLzGVKE9PH9jYhMgTltnWnck
hVQybSVHx2Nw/dQdt6wPyJt2hXSQY5QEUou8EPFcj0IgHMcUQB7yqxCyga2tS+Vz+nHS3cVFt5cC
1fLh/KcHLl0/7GMlNWuMvStQ2EeYU4u5zngfPLRUsp0Jh4T+Kgm4VHI2KemQUXV5wQaK89s3LqDr
Ym6DQ/FDjsL1NB0VbL28KkTaOAHAyo1Hi1B4etsME5Y6W75W7cYrFFQYtVPk6hDvIHmCrhWfTtTJ
2HoMmDFoJwI9dMBkNch6nHSvxx8gTU64YThIYResToc/AaRo5b5EoTVZtC54x2I9bRn6bYTWyrpi
rHY8zGW2QSMQQWc8q/Td3A/hR9HLM4i0/LwDpRav/7Qxh2JbH8kA9DF2B0cz8Hr+VmSXfcUFiPvR
POW3fAb627fCKSjhmv9IMye1oPwUsNt3ss06G2iirAAQYA7xG45kLIxIsq+VTRn4v2MHDYW2//lk
soEZyDiDceL4TMmrAnGHG1VSC27lN+bIjxXT9Ey3ECIIiQC3LEQwstetnOfVuf7Y1rWLtmPSSRBg
hLzvBfe9lQrtp5qGh8DcW3usNHQ1iX5jTNs3tQdQdEYFdILHFLvItU4ovVLokGGKHAnVRg14xJrn
SwblOnTjtjjNe7Sn1IL5seAO2Roty//PVtqG5pDKITyJ9i9p9a3zxvTwvlOKBmW1FcBgt5t15zmd
cFu45G7kUFyZXAgCBveZftWaQA/HbjV/DFRJI/HRtFf0dcQ18eedDvdFKBeNoK5YuvFzhYqg7Es8
nDzYPVNeDEUwaBf7/p45uKN9ZA+Brpeirf90kYjPP1zBgab4oRV6yglPwSWcLGAoPehP1GozzsMj
wO67FPIuT1LFlsu89qbufTfb3p1yhQ0GIEx7GW7xkoSg91skkB60+EGnKJOcuHx7AbSlfCxkZ5oh
bRxmEFDkFRltLdcTxHzW8xrEq7EkNrjV5ufoet7D58CAcsJHT59Z/UuuLBW9huPE2aFIpA9xalVj
g+iYVYKPKg5sebijyUAwTq5rqrSJSwkPYQfLn+0SwrjlAApmWuLZH8rMNEqbdIsQd1MpWWfMZx60
wxt6haf/K4fItGP1lLLXpDscVTa72G4w9NQNQskC1IdLTto7Y750jdDRDL6iB9TsCicd7CNcK+TS
amEtmSMq119BBQjszmjtOcwgoV+7Aj1kNXm/713XnBNafcUrH3Bqi/fafnT1sEiGXc21zHwm7pYA
Nj8K7q5zMs9OHCTPiq4PZA/axcIFx1wqs9XWuUGmIPpCMMlWQf5bCEH7cAQuIA2U8NpJ+CUZ0OV6
wkBxoVgYm8ecPAsQV/VWGzw0u8wynLjWT9Mg1uyB0AacrJgxCA80Dmnf1TnkezDxqzNotjwsAil0
c39avZJRQdmuSTy5CFz7kujYxKi2C3zS07m931k34nbYgA5uZOGU3vuVLfGz2RaPLbRBk+OWSBxW
cEUDoX6fC7JO7GvEdpID02cfcqs8cyI5VI1TfVRPfifKfuBY63kAO0visaIxzolDLJCiyzv7F2la
hk0aR0oPsEtmwk5Cdv38qi7KrVxv4i3symBr6mHCYNHxZn+UNx0b/R301hQsGVO1xo9jpgqX97G9
ehBPmOrt+l8p9f94YW42OI2LSYh4bcFapgw87iveGRJe05g9n1ROXjjxz4oHzXlZ9KTfXVPgX8eQ
PE+2O+zkKRlJEKMxTXd402xi+Mc8VQFzwT69wMFForJ7F2SN5bdqKD/IFEPCl2TaKZIO4/wdYP5V
ufI0g1m8zu3tFPzz6lem+7kRdUWEVV07DYjr7+zBpTSLasZR+uRNWARbfs6WKdxRrR7lic+h8Yvz
mmBJUPdFjZwJe53YQuVnG0OpEDB7kGj3di8NtMFA8BZI/2MeWNhaHcGDqdOmoD6MHSUi2xOVdu04
yv5Oc8ZJXjX7r1I5WUAnJvkAOIFuQFxZ9fl8hhzsWa+J7b3ivhAOfxpKDnVQWmUqM3F3RJAVDgCC
fM3NJ9R8QtpVi+n1f+m02jSwH2Vj5f5A0c8uZ2qsULj3QxReRd8LB/Gw2eXEe6gUFCMCvSEz8S6y
YnMPitGPKpJYRFXOB6wrtJF5F2vDpTE0XKtJk/eWHER60sJjpI/q/lIGLH3eQuoIgJHRVfgkr/32
w8318TIIVK/ST116oPI8QiBc/J1Krs2IZL0bAKUngHuhIdLSJYQRF+kiUH6Zia7egbWp0dRpCwKg
PS0MoMDUug6SKGUg7ZWCzxtY+CbxBNOP5utEoE1Y/ieOAKA2tfsRGVay9VyfavcY5xy3wDQhskR6
HyRjoqIq0D1+pi1/B+qrXqTWgNCuhqyHsWFikH/KEHjzu2k9mNzwpeRz0w+fzSGYlw0JiZVTOxX5
BbfuRu4BtjK2MTJf+DdO88NOQ26rAGsUJzoHSQxoyKfBb7bnwyOR6wVpdaKG7WSnXN6YfCy2Ce1+
odzKkMkasjA3ZbZeHvEn8PwFgztFXjCfE0+RoPj+gheIs5sEeGMTOEHbltvdRPfndZWItxrCYEHl
kmWpdaE0Rt5LqC8ypVtKnv8eEyHRs4digGBPWMS2UwyuQ+C5zO3AEYm6MeRncgcHH+sWTSz67G4Q
AjelboRSIErW9Ln/lIA3Rh5lQiwEs57ydSynogKxgBRG0EM5jzu3lluDXtphs4a200tsCCDLZ2iJ
KSUQql6Hntsq2wsZTd5trVv5Z3EV54DPbBb5Xou+aa7MGNHxhZZKszbWkRF0nHmgaZhrQpUlI5j/
gvQ8B38+ZgH64NJjEeK2HjXJ5RSVwk9a9GCigcsaIv7jydm3GO1Bhs/QmHecdcyHld1fJ/k2Ptrz
UeCtVPmMUcS7h1lLE3r5S4IKhURo6zuAQuE5n/TtyGy2XPLlFUPXLp1MkHDszbep/SEwf92vj2nG
EizabsK6QUHUHioQrPVnBX91vE8mD+pfuCaAJjU74/FB+RoOKp/EWn7g07OTyZ2lWMOVO4IOGHop
rJcjYQzZDNCDjdZ4JbtSUJ9BJQVGWzyCB7sFn4kiyFKC5jI1ah/6am7NKCNoZ9uoc2N8fPph/6V+
Zu6fpjiexolzKPApxlwkeq0/M6w28NQ3d+VZ8/3IDmSMSAi98h3xMjk0cS61RkS2AG7LAC8N3PsA
W7hZ9GU5OBHNCQXczf34iIV2WrPzgSf9qo/bgZx06ve3d74UjXYw+QwQO/8ekTyVKzWLwseGm2r8
mhY1eXOtHa0mFdA/S0K7YIhxOA/p7la+5NSpRtt1Fy1KrEmTQabLAvPXy9sSxilNoPwTHGhzvNpl
aSR5zmSo0nye0tqAsByvt3X4SQd3MFlIi3dryF1q8wwSa5YGAUAiRUxwgEtkB//qnX8PLzEdkq7e
nTAxlumeckSwrPEt/wSN/Hxnbxo1OdA08wzG6ZuoW7URVBTLuU9BzFvRJeNoviUyU+c3dgr/xh38
oor3CG78N+IK33Yz5MLH3rCmhAFfPgJgGLMAtsgSVcGsRKR9QQFpiLAxokPeJKQMANFNtPWmLWF1
Dzf3+CMLNiVAaBucKT4YHqPJuWWCtju5f3LDCg/8nE5H0ykarQT3FhS4AmvnXHPGHYXAw5sTTm/b
Q+iABX6Ai3UaIg1FWjbKaD3+KWM1MvwE1ikh5oHcVC+qFcN7KzwqF6Ealzzh8cEhhDoJhZs0OK4L
NNLvKIZSLFAESCxyFAcw3pL08timXEJr+AAofcV1tEgCJ3YHHDpkHhMn0T/l+UsLSS3NHLok/onU
8XMG3lzxPXohUf/OB5LEI6k6P7iN1QMe+Ys16nE/NwgKtPbkVoZ32ObKCJhmUkcbgL0l18ZTRwgU
vfqmhf4jIfibalaDUxHqb+xDdrOmfzbzLeq3Fg7llboQoUmu5DWyLC1cZyMt652joT2zwtQIN9Ra
50brT+wxGlGlFt0zJ/rh+04gV0Dt+LWfo1kIBUWMBez0RkEBhACl8l3Z0Ea8mS9w7alwtSiBiAOa
bZptWEauwZbS7FAv6qFlDZoZRgnvc+/9K8QAPcLzWvzdIJeXSTm4+ydfJAoDAGZnTmxos4FYjNAP
ItM88aw9vxcurI16BoXh6Su1SnK9mNgURPaAq4OTjE5Hefbvs5eMTOrneIzQbbnz4tVjoZKN14DK
AH46eg5DtdgbeumTvtqb1VRM711rE1iXD0nymGaxAHRjtlwcFA3eKg2OTcNa62QOGG1SKOOCqL6f
Hrwo7Jw1HuwwtNNhMd+i7nFiD+AOM9Bgt+ykjU6+VtvADHxBgVAMX9zM4gfKWl476eIP42czM7fA
ePrQUcPJ/srQQiQehPCsT1gQ1xoBngzsZ9FgbZE0IdIWJqgF5+hIM4l+H2/9vD+ovog4YQLu6JE0
tOKOlJYq/vJAGad8lS4jrCE1YZlM6YQq27c9+Yzwsq7JMSifi/sjvA0Yga8F1QeFEXcMa0+ce1TV
NOKZhSUW8j2O+hl+TFbgCzbeqHB/EmlXSmJzlGbAUPIKPzZtXvBac4uuw1REoOAxKt4ch5WwWI9P
vjATONR/67jtbnVUhZB+spPIKQDjWK5d+jLofwAVtxLx3JmJrQukQpqOC1adpU2aMo77Eu+RkoMI
ISPAfl6piDweUaPO/zwtLz1tyBOBqKjPLD5wrmeKic6vPD0txXg4yfW046EPr8D3wjmVDjYWocVd
xk9HcjJcDirTR76AbNIogSfFDoZipEKPEEYmBu1WIXufmGGW+MZbBXqZpzK9vZy3DJIRDwxUH/xi
YzXyWRs0dscnwfA22UfDXJw4HVDE7IgwtC3c5IixUS6JKyvC6SLirYxBdtXqnuZidDLbLdl182DI
wZYSo3a+ZZ8lrnzPGQhqQSgqiyMaU0k1wS36pbKdAqEI/w11OQ9lHqX+JAon2NsKSe3+rVgvJ30l
NgdZR9PlxYZ70uL1qLQpsZVY3PGePy2euAqBKc2PIraSnex00zSbWmVQ7ppj2kAd6wqzfSPrx637
A+Auj9rjACjSgMGc6ylCUKf4zENsXUxkF+VxeJ6tWOchUbPdVoIKmfUn+wbZjNuUCX5AaPPWVO6M
ah3NQjNDIBBR0RsaIHP3qZkv9YX0bwkcGxED5dHgaLEl7CdkcHcfYxlmFnXhitULszQV4IP8Qvv8
3zortHAzF+nZIMYRJTdsqm3Q0QpW5D66sTMFQ9KcOmBMQTsMv7c8MKiAiF+Q8mgPYRe5gGE5qcmr
5HhrpcN0TmLnBPd2jx+d3ycVW7anwRUsJgPLOiEzq8Mzmat/M7+XEEP7i+/kzZB4ch9A6o4HWmVx
qJxWHpeNpAuVQmFMaYsvVi08GMRBkPQiqTXLslxWmVkolecZyGXUyjin1nBxt+dSkYRH321LRui1
Nmq1Kvvj1QUyYu2ud5xvCz7q/LVkfHyatVrfxBOikMZwe847cDOZHmS61Hz0qBtD7AamSm8DhxTD
sdA2qzQjoaKK8Od4MJXbDFtavdy7czuPIPcRlDQjTr2w4cZG08QWncLqM0QaSaIrDbu5bUwd77yf
GJUnXLXpl6VFUHja2N9I+H6Ip7qw3EAM/28JeuJNjZh2BkSmXK1yhzhUSvw283br9vVd4tr4iEnH
Ou2EQ2JpK4Z5PdZNBDaCrkrFPlTtvtMVvn2lAIszTHHCJtQAihxXWPOcOYU5ob8oSCyl1wzmvf8F
8wmEM3Z9488y02lxS4eXNTJwQnJ6VjNhcpaTeBluaNolNrLVTdxmN8QiE5dA9TVnJTcNtBCbCjko
9X95UvG6JR4xT1IdSm9Umsk0gvj7UJFW2m2L1Ej/+wlZ4uG20lnbfX76Dg1FHekZKwZOeresuyjw
mwkKxyHr3KsDPLjXApzjcfRZAQouiP7v0pI33zvdIo96AtMdFwbZZ8Ujvb8caFo0Y6fzbiPI0FDQ
hwSY/5tR+ZQOe0z/rmInu/9r7RFajh1JomdxVRxfqeSxRC+xYOarIRr08AgYorb2g/PRRenFW+0U
bgpueQ3upwefQkhipk9/Gjy+YmKdc7NfKiDKT/HXmOQ5pcasht4lnPu/ukZNe/YNRQZ3DnB8wrSv
/nWWQOK5LoBgcAlJdHO1uSxzv0Db9Xuco0fGB7QRGebPumfBzHU0hLrBCceLrDa5vZYmnM7/5u1R
t8JDeojndu6fQzQDA8OHV8Om8qVwjrCrJPUAoccp9BeJE5Ue/wsbCp8ReAdVBNddNdyaRVJgxJX+
TPFhs4m0eI9u61JQMIBZiVNnXkm666kWduwpk4SumUxcZRJ3HyMY8a4QdN3l7NmaRkIXwddj405s
kvJ/cBPAdHLzC8crVKU+mAz2ulPlNVvLulC7DECl14RlPcZU611agsAL8rxP+kRyoVfk1vlyS+yL
jihwgRBkaprVcaKa6K1Kx9zazILt7VaTjx01e55Ld2oa8sHx2QV1uajCxE+VGSl4pmWm+vOFFJVI
YyVjMOHiBUOi/XGEb+iSPQQ96LoraDgcY7CTaiPj6qMa9+BfGSrdZUNQd2xNbt/2Ds357cpocEw+
boL40qwae2O3yiNk3LaEyCQqe8zIWc7VfOPI3SAtAB2OjDmc9bxIyr7ARCZMkGMMVid0UbH1W4ZY
58nL2qUvEeqGUcXzmJcjewLIVF67qDJNRZ4bONHHAPwE2qBBjy64OaG6ZOonQ9GGOFpBS7fNmC5v
UGXBYFtvLN+lww2m5MzO4tOync95O7TLa9j+RkoalUR+t8loQPXeToCgkQhBu+5kd0M89//6Lo5B
+eNfyisEFeYiwHdfjzSAhx+iYoGTZ7b4eysR+n090WWpsbhXx/V0GegIWmgvwGTcAHsDOduSrbSQ
CfYhf86+lUli6uodSIv6zxAjWN8may/UP7KqCYLLcFPF7B5H55gVoZmoYIxVJHwQq1+ZvUZD+LW8
wX0WAFWr5qBzolm9d+kyRdzUscik5SKKLTcs34+gKW4+4jJ0aqO9LU3PSABqyEkW+EsxNuMYwiso
fVZR8mWCgkErmNIM46GOm1TvWNsCWOY+lIdOjRpVymwanxIrAHEFRnSSDGvXHaNzxT/VLo1EsA3V
+vo+HtpEcRMtUMKUR31S5BH4WD5vvWesUyz0ImLvwEZvOTKzbAQr+b79r3w50pyYbWfK0CcwIhTX
+mY0TEf4om/nGLSkgOq1fqe28Pt1TEdW8Tv9/iimkgnCDXyfzAKlmEd0JQFsQqbtDdSAXaeGEYM9
cLI/hI8hYHio5c8wm++5bc/ynQgW1h7NoGjfVVC7B70OqczgJdb35d+eqbhY8Kjs1M5zFE/wCgVo
aEIwKJ44vSMRQ1lyNDefnUQLbN3bpnA9dbYRjQCyJzgcVP2LTRf2apgSHyTdDqXP5o4IC5m6pPbG
FEoUsLia68oVkcfJnvDNJIXWHztHf9xFc5PfEg21ZwqV0V6GDZTlEd7TwCAocsB0YQjTvJ2kpk7I
ZKA16za8s/Z5u0TKpjEo6xurPSU0KhviQTRDHIlEBBa0uWpq4BN+rkow5u3o5fCacm+H8/w3rRsu
KNoly3j9vzyx/pIHX+T+eiPpQ3ujOswrUROJ0M2XU/wf0CWhKeN9JnH4syHF1of62dG9HdCmcX7+
j+y16CCaaUIIZhxWUIRn0zlFguUKi6ksrf5EAQyDbrtW4Q5OPUQdf8+DFjXfvdD6x4ENSZeKmyCA
Z2cmbXlU92C0Bo6NIzmOOXeVxuhDTTa43J00cn7uNdz4qUkXukIXYfhNL5ccVs/hcvyQMkfpi8c+
VjrfxkKaKYgffH2Tjf65ibMnzPnzXKlTHhwroceiSSjnl1fmoPKZXXCqkaj7fGp/Ju/b6tVQ3wdf
OhyphTWvg3I9Hcm5D4t8ugj4CCtZJy7oBiZGvroDbbnb9oKlb2y1gajBmobHF4lKmYNpCsA4yC+9
lB/SrKEYLihOdjrkS2jhUZb7LcaENO1Czed+qTwludTH6iZs5W95ElHpKhbswtRqqf0XszH3sxEG
Fkk1Eh3gX5nxiSBNp6uPzPSxH6LZc9e1f0bLwQCcHMDNp+hI7WxpQFDzH47qbA+n3gbTElQ5ifSf
nRY2yyrEN7h2Xkxw1IM+fHmz8wacPOE313iXQtqdOd0/a/ex3dLum06kAYcFu4URiF3rIgVxKWrX
BssEVx7JisxrE5D5Xyt4Fsvw25x8AiOgoGXv6yB8PEiqG9YI7IFPjoWKHUfrRakJAvXIOYpUcdA1
7rkij37E1lDKDVZbegLvT81+P0WXfGzrBb3z3ibZMsN3j2IAxYqvbBhBYAw8mw+uGjPYmsoD8rcc
SPuy6UVdcQT46kDUFR/QNqySiV3nBBHjgPSU+MXhJV10NUprepJHqNHLMGkAr0DZ9/6F1FiwhPRm
uDGaSBucNBNHnHAjr/g7/zJtFCsm2o43kzh+p8ycI5v5vGVfIuo/Iwvw6/cmxbIP9h6zojbtxSlC
YEkl1YmAmj4YMej6wRcMPoppIdSPCrpzTDpGn13VkIB89MZ0EzOErgOPP780xJip6Wsh3cCYjwXN
q+yv+Sksk+soVJGD9JyWFb8hZXWdOgE28LPhbXtmM/jiVInF/OegPcfL42ipN6cilU1IMnXgXfbc
3crEsllhHmObZD6uQ6ahcI8XBxiaV5D0IYnkZuvHyQpFEoi6j+9wP43WW3IPhMhtBzqoMQ36FvC3
52oivWY2rnQLA+lORU+kPxqJBaO+aL0ueDA9NGCRoLe7lbeyLpQTw+JRKrTXOQiZlSdtygW+lA7o
tH547G6KjfO5j6/6Bv3gWdvywebuCNrbq0TYbFwaKU5XV/ok5hCRfTb92eqqGx5MRZeHrb+2QmT7
1HV3Q0/LTCcREeNLZCGLMf6mGAJaXqRyN+b7atWY92Z1LcUqiCAIUgUfBo2qYkoxR97wmetXqhhk
jw8x/rZBbWuuSmCWLI5ht2hfFlEx9JEEY87HcRU4zIaZhEwATM3zNFIjdmXbTaqrM2RlKDyplCc8
ApjHkzahZJHjpxPv2QQWHMNXufTuG4TKwII+ddh24L+xukyq2khvGfyiY9plby3AYAaYzD6WE2hv
4P6ht3s9BXRseOpUDTW1Af47BnpqchD0D/W6hbVxZ0BxFRoYrNHK9eiK9Er/e2GNVWlxZRHJoKDu
T/IDNeq/eVg/tO4UgLqptlad/bKH/my+AUJzLNXutG0v/Ap66Y4On7YJn7KJBF74LtBFIfihWKlJ
/cCcJEtFqlVffq6mF5+bpVbZiQmunUzKSOZwGzgLzcAsUSp8EQq8bjtZwgLiVAgTNO9K0xyWZ0kP
xitzDMNk530wYnD7QnFy6MUJfW8gqJRb8DkHb8JKqDHDugUP78LqhLhzNCRc7FpYsfbXVio406+c
p3MKmEOD/YK1R879YKGKJf8dtlDY5EI63B9Mf3p/N9A9CeCDHsq1nKowwcYUAnimIZXlQqeHo8Wg
uq+x1y3bxleip3uqEhrAK+3IFUQrIGBZBun95HZqC2DRjpTrCj8yddAYE/VHgsXTgOQd1F17zHgY
PWRd0q+JXP7UOfS/JNz2fs4AIZM3g2aB7Qa7fBGfC1HXTCb/oITgBBmHUEqXJbHtf3mc5TZoWoTu
fitJu4lM1snpMfu2254igT0QVnT89u/F73HpHZHAq25AQ76VJd/4o0Jm2mvRTOPEXm1ICmjte8Er
W6UblKQFqKkVc4C4CWfR4QBQsPpZywgkCyEs5Lyb+pw5Na8tBAY++wUhlKcjNzvyE7jbAnqzGg64
zx4dslxZnSKl8nWuPysMx1C0P821kR8xNCXrbFgtYV+89Q409J5qcieXPM2dbyntreRecpINjT9r
OqluGA2mSCpDJ5CyQa4cYjfodeWvE7B94thKQ+TB2Hj5VeG3UdM9t36nNHkNo0gTthHsMTZm8o/g
zcNC55r+iQE2wzT/BcztvBzDAYh4jMRGPRW7/N/lukZDfEstz1nvPJR7GsTqLQyrxNDe9TKDP0JW
8+LTzYOla9czkudzCdYnsEBW0qOt5Br0bm3m3rPXAvRN/RKCAdCMRGVpPWpsVGUWcU7LtEmhLsMC
wqOGt0bWry//h7keEW285wqerW5Tld2tMOxGYdJTAIHk7r3DWD3MuILL3G6qVJhJ2wZWf3kWRbxU
WeYTVgHm1Khs9XJCzOLopHpY3UE10TgPulscd/Emu3NCT6nmYdI4EQsormnWHjFggGwff4Sqv3PH
UVVVFpvsGyFKbRSOkIArPyjMZqic8NmCal5Ztx7SumdQUU3Kor+nySjU5B43bk+n2fpw6vJx/Ng0
sBPPOoYSc9kDpwdaAHtkt2Eb+LQi5toNNwHsrmd5InsAD4NGxjSlrcS/YOu7ffDOdkV1O0YBOm3S
6lb1pESL7/Fwwu2+MLK7aXqol+rbD8eY9n61NqeEcEQSTFXGQwqsYE7XGV/18XUcI9mYqR586hO7
58RWXxdhuir9vFvpNjgRdJaOOlqOy8cndxJWkBRLSBbYYnRfmUYwGAmit3o43+Wtmw7vm1CTgVXs
ynI97G8PmBwJLCJ5k1Ynijle+OAOV4y26fEX6XESYbvGIYTkYLzvo4M0m3wZ/Mvoa9tYpCsM6u8N
paYR2LhWSWtbOPn9zYHf9XN5exdM6/ZO8Y6VqqGuQC5ef3p/kr8febY4nuYJvTAMwYvZ2wYvNaAa
+96bed3KwMP5zR4ADGTnJD4Ywwu6zvLv3JaUzzsHhm7t9p2lTq+wObBJyM0FOjllPIY2Nznh3fMa
urUFpFf5cNqC6mPf/I92YNLKMkZ/sgOsR1P2nzXFJviGpQ1L/k9varam/VQYsrLlrhRflkj+iudL
oVcpHPDNgV3v/Vfu/uvg0B+g6Qlp8U2P/FbXKC7eQApTYhpxipLCdvujInurc+xiSYgWdLiFBedQ
1E8UgEQvdF/E7vidnjj9ERgDmMJgOtBi+cBe6qSUAE3SwN6nLzKnLdZ071LQQBLdAoOpZK3C7g1T
cczdg+8f4FpHjgHuffxSur9mlbnphjo+3WQ52z+cPXOKClMJAo/wAIWArWY4dmyZNLto5VHM9akH
549SqLZEVmLdctPb7GeWMWE6ZCj0TtWpK5+CoPPuaz+Wd6+nDmoOjF/IANqJAZKHh1muT0ok0ji7
LJGFjN5hA2wmGpTLkOxKO5H/5HxDMMWIZXQihg6exzVZ00+WGIUty6yJ58Yu+HFRxDIaS+mDuJz0
HZ5fUvvA65F0zncMTfyY1Q/8z4rVj1w+fHB2p1TpC44M35xXHj2WvBETIVz/6T0rbDkZdTWdg1FW
4GjPcXI/OwpqEBHXO+dAf8BqSMpPvJ0gZMLc2OnFreS2UDtNYXvCecgwsQP3K/RTQdC9OTdLRcyU
mIqzDBUzqCozemkMS19WDENnxEl2bKuzO1sQTZQAdd1TL/ZnUxOEF0h/4guD7AaRLK5mFsTRWF85
4RDtFDM6+YMkr+fxuscXPfHimOOPJvq+PVXplIviDPn3sPLKN0W7hw/9TwHkflii8dgp+Xbl3Kql
4UhCkYdM8L44IIFS8I3RDNnUSx0Plm60np0VIu27r5f0TG6kg5S62AjTFP566+vTITJXk1zxNKFa
8BuViBeAZOaR8FwdFOIzsSeFEbSD+SVTUaVENKYiQ1EKZuE97+Rtug39y5y6rOXMMs2no4ONrYWl
aqqXC+AJAOqIs5u42SVKUehguyPyQ1UMJwvaGgduDV6c/tgIwcwLDRbMaAiw/KfTjKPXB6ONOmyT
pmNy8ZIek0Qyvt9foZzj6Qoa84Mo0lqln794UvpC7DaBzLWkYpURlyWaTXEtJyq8cE+h/eluO0MU
7Iu2pCGDKUVoCwyjcd7pj2rxm8NrY10xleOiG4C0+fDoDxfuZr+0M8Wofow/DLoup+J2tqZiC7Md
nDBl+n4+FZQyrLdznsj+e99xjuoqDKNRdX+lg0g4FOoasgxbx2zguLavHoFtQnB7aXhQHlZjyaeA
1O85UtUwAlCHbtFSfQpSgVlQDNanuwjCGk6K1Ksch6tbdmQp/EyM0ylJ5TrPbEqS1VXfFLsdrqff
7i+MgawTXNGh95ahbofJvWW8E4F356rhWpRI0Db5E3oT/l5XIyWOMg/flJzfLdm+bRSAD5ZvoW7c
rVVxAPwmVgDW0JXCBJCtVRDL8gNQ4QlKeaHjEqFO3zypg8qaXy6im/x4+/Tb5MUu6qP22yeV/w6x
KX5PZ8stHr3Zi9B/8Dl2LrB1QfIO1hHkMW2IDlUpV76WLtEUcfkVtuEAnGCkNakeFJWjPOMOCTFS
FhlaIUxtgvnxsqoffAUTIrYsB/TsRvMsWJchggpAJbkhMks4Vjv2eXV3JlOk8IO4+A64wRAwXtsp
J6rbOe73lAjeBlIG93Y2t0PK+QgyedBGjoxdnvPwBiWhYJJEh0WWZJLx/ugiyEg4qDHSDPL2Lg5g
/d1FHVGlTXFuwAks1sT/Dxce/Pd3SU+qzge0/o9DCzWj/M7hhOt/j83A5XPJgneFt1VrY0plrSXT
+/tHaFRglXbt5yCsMYNYFkPtc3vLD3Y5Dls+1M0wip1yyE2JLzQmx/F2dRclMC9lCKoH26lua9UX
YyNpQEUHqHisSjkTRVw3OPEKPA1YlRPFRCSrz9i36EeEb8McXUsdaJsA+BfZd+CEMpM50z03drpP
xjrOsGXRV8BhBh3ZmkzLf3ZeYN/MEUI1uW35sxXOD7IrkIX3/YhTJ2U86Zf4KTmS37uKL1j84Bc0
ouW5oT9H1j3bhNAYYluGHJMj1q9FCvaGzECaZsw7oLFtpJ9GobEpDMwJDMFMQD0Th2Aw4VC94b4g
XfEW5sQiJbMJRps8IALN6sPZjvpp/QKcg65h1r4paoSnmqwe44CCtr0F66F4zvFskHgv3q+CBBof
Wg562xUP2VO0po5qVOtO0Al/VLi5bvBhVY7EN6aWLYcDMbZRDFxP8/ih3Zmhrf/k5Etwc5fc6Z57
gAs5HjDwe933x0JRyZJd1ByhT1J29AELU/N7aWF8mKbmDKSj/FvT6k/c48yLeZccgt415LMpnWyw
CgHdZcfotGstr36xKTxUamdhB60SOqz0YLzX49/SaiPRg0FXtUnhlkvrmnwUcFRdCG+7gY3ppoRw
xbR9BcmudqeTAe0RDzz3HDgC1eE0Y4usBO+ow+15w2ZxY2Fnjsp9BXR5BadE+/K6SbayGs9JP2hF
bm6sbZTB1AeBpLmnGTWboFk08zEjMk5deRZ8S9Nxb475nEVwPag2IbDGqlcgxXip3e+MLjrgxLlg
dWKJFtR+RT9Uw87LSYiogUZTDc8vMEHV59MmQzvTBu5aFdyDulsqxzBmU8LsGllslEnv17WxxLEa
65LDt4V789l/Tu1KttZtRFhZ3LtB4cNm//hT3+oNBQ87evlVkuKIgK05qzUiZiOPYe2Qi5YIQvoa
JmGb9yZdp9Bkl9anlgmJwuvGszv67F8O2Vw91rMzhHWOwdXi8avHvTGK3buJc58gxzTKRbi/I8mf
1es6IlN/gWGDocitBKOEa20qJOXkOb23z4Diu+XNeJ+V//7RoRoCmlLDyWddR6qQE3AC0wzELI6z
QE/dA3O70U40RfQbj2FirJ3qaWzUF1QR1DkGPx6/9Rc08F4/4kD7FqvQPw15yOfpCukTbNafZk15
/fJXCsRRullBOzmYrXO4cuo12zKU12SaXQfifwwn14ldFRJjdDpdbD1A2OKcWiWCNbhAG2nnuSga
+wthzeujboK3C7yFUU/V2woJ/SKUA6WBq/e3zMzBjR1LfDJhyvfVT8/wO871WWOFFBw/us6vdm+j
IvueiQUJj5+xer4yps1TW90cnV2RFxkwghmQF1rz3OaRaO7eoP26PzfOKx0A8Zb96Hnl4wSTwAK0
6q6qGsYWEBnnDIC55WOSOo86Qo+bOjJpYrl03iglwgzLMiXp/QDCyUrNIF2Xl/T/UK/MqPW+7v0d
snSN6lRAjBnSUkbRnt7RP+LeVY6GFmQaTvaDrVCNrCkjkLWTspHcasaqxYm6K1Lf5ZLi0qKeLXre
a0U8pQK4jJBQLxgsIH6JyyEXIIUjKAY4f+DpnzTEyqyxG4oAhAmy4oA96A1jgpNGS5NUKO01ziSO
hYuf/CSwqvG79rA+RghhZ+J9XW+PfLE0ueICOYhjeXs7yYAXoxNWxWyMtrADH9XYezoy8U/4Y0xh
OOK0gABnmBj35sNL/IAiOXJT1ew9CHwbxCY/ahX3eJx27fEad/R+3Pqx2YOJc2tJTk8xuJyb9LA+
n9IZIrhckY9DzvF5QmA85q+xwfnMEcc/YazVsC0+b9YJaQvqo0MO+y9tdashsBL3IH2L2FkdPeCZ
RibUnRFxxcYoTduVWToHlDtmKkKrocUZ9q+kGNQZ76XOZLan+GP/bZH25jQHyg0kXnMp+QW1DkvE
jZ0delKSenFelkXWx0hNLZ4XzQF2bG4x+azGtvSidCHm2hzCLBCQvSunupNrmEk2HY+7dXOc8fMO
aoxnyFy/e6Q4ULDufKgdW6pMlQc9hcbZtq1l0mPqaHErb57Na5M5NqMC88imAKSzewiSsm5rUHY2
/XE0irN2+lfNqZ0A4vuuqtYS685AFZ91sv19+gnKupjN63EPA2mIWeysVExAWdtuJFFW6e10JaNi
GPr8VKCguFbUt41A13rXhYDTHmz4cIpWTW55AkK4Cnfq5e70uOWLMLHrIYOCQ+9RxrNsd4DMzcMU
epcbhk8z+3jAt/g5gEbDGls94sjO22gAVqrZGqYdNV5C1jetmlKnLyrohGcEHc3Z8veY0E6ZOWZr
0r/his5Xbb8bg55QiNj1RVNNBWugDWvaRq52Nd+OQb2pM7ovG1dZa/aQ1+mc6CINPRIrQHOCYDy7
IMxDajgfOro1I8P5YEqigpf1YZxqv6qEQ8+kU+UMUmk7wYEZLag6fD54jKfQ+E/9y0q2GFB2gQX7
rC5Cl39GkFgpkKDbqOUhsRwZ4IYfhKo+cNPwyOFgkOuwjWpM/srJvj+jGVutz5fh48cMHQQnnZVR
r+bD2zc7FC9+k+PQ4ljZCrY7378Or3e5jHAEEEWREkVgJh2O/0WBnEyDBZrP6y/MHDogjy569Bw4
srLyLCIGpheKPgLg5fcyp5msjGjcc8ngqkSaiw149zB6qMDkhTuEQvF4B3J4sH15VcBasBTyFnt2
bLKG2HWFrWMmyj9xScc8bblhvbIzmnuD+I/tYjqeUQmzpdCDxXy1rMnLMmLtmxJjTpaG9isCDVjt
6ZhB1/8Zf/yrP1gsYgfe00ALBTjGrnxf3i/yxZxJmN9+lj3bvHW98/6xa1/TOzedb/m248zIniK0
qILD1a1Ej/A2ZucHYdkTqDIUz4Kyu1z33V8Zi6v+/nB5rAk41jsNb9ldeHwEso+4NM71fcsTlnkV
YmPfJjqdw/3C38tHkgTFa6kkaTay23T21ZKqsdRTbonQVJSbhE6eanNH2xrYg7YvO3h54gE7lEWO
UQqf95khclTPl+gxIDSM5EethNXHW6BYAkgFPtFBN4R1Z4ObEUJqcaowDnr/9CpoKo5Xx2tFKIDC
rfiOTbpEZQiwLwaohruMjzWCTCq1LoDt1mc7tYU7SWNl6FNDc7UNhuEV1lGkQsHskgJhs0xqu8Sm
nRUU41cZiqUfL2G6OdZbqeAFVfZ0RQ/v3oRVg/5z3QljSa+9j4S5mhXhYqs+uudY0RApLwcpNDum
IdzfGcotL8o+aUUNq7buYCgzoQO7RR1UaSpBwl7diG5bEzrC8dA2LN5QXbOtrlGmHRuOmirQoyrB
OOtNrDAB2MXwQfXrCEfo467eD9ebvP9pPN3gXEcfGuWy7l41Gzr0LmO+k75VX5k3y3FWRz0EB6Ty
MZsHGM4UARmI+zqd9mw+vPMjMCcykKCpG69b/2z3/zE/Z5howIOXNnTUUrU21UvoHDWfNKfdl8yM
0GIUd+LI0CtqQNOvKGkGRSqLMuNtVnPF+epCwf5OwEOjLZZ44c0ntHPo84CLdj/K4X+pVSLvGdBq
FgXy6b4TBjRKSBG+u7HCx9OieOs0KShOXv2uyyMugCf+O25jw5ZYpI9SoDqZwAbwxVPji5AXB6zj
EWxPyzIs2B2IYpsIQpgvVNI4IbfPVzqG5+b8529WE5rI0UkjxzLvgr02/4J8D4cPcbzhs2RAvVib
kErU5uz9NgiB5GQos4YTnRXrdouzhKAeg9O7DKiXVS2rjOPVJiOIM2CaQTYk7KAFtVfWuvvZ73jH
fQ1ItGbOlj4xD/CVX4bQD5U1/b61nR/FZzYj/Pt7KFQOcX+/f1SNq47ar8hqRT+Ogjwzu/9ZftNE
VXywJ7weEaw/Pr0jbXvfm8Ut+P7Dm7OeoXZe7A9ddAp6Hd61LdZh7tofjy7OfBXBbCaxhj42doWN
MkuIlu39ny6Dy7ae7H1mgfh/XcP6BXhuMJRCLWtZzKMJ+joefoNLrdUh0FCWiB83TCB0x1e5UT+1
SEKoGSqEy9MOSjMba/WCBpXkqYtp9yBD6mAgjlEtOZvee7APSlbxmSVyuvmn4LXYHOv7RPfRQru2
zS7rI0YsAHrBhr+hr61scMEYbYroh7l2CT9ZVDFoGaTRynOyY5eIzZdw0fFYChyA10o1VHEKaFrs
sBpEaOiZk2Zh6kHdmia2sBd86oWrshWvUkeGH0uUM7jF9eTytJIZCejYvVKRroJFFNVU+xpecQdo
LDaJHXNWAZe9lWrFa1zF5BaeGFuNnP8bkCai5apfRZsp9Rk123ovpF2hHpv21s3TLsNqlkeJx5NA
t5tuiw9QtQ48Rh9TWq2/53OPGAG9eLlZITmFvSS8iZjLGgPqdRx8O9wp9OxqzpQjVYZXkgCrof0O
px+LA8GfLwc3eRBjkpOJSBTwJyHrmju9UFyYu8DXY4iEA9KtZbv344/dYXLUPU3Mz+1D6yy8O0H1
1u+sLvOxXTUPG5m8BEhNKQFKFhe0ws/MrGe58p0ZJkqQNV/LN5sf5NrJztjdHccSOnq1uW5nkk6k
n7zHb0JTWi9nL4E8MdVacpCJNnqczIzvDJf+eMeW+RoeJlTEr0azK3PDbv1e8Gm/pCOz3kOdw0Y7
o8srAPCQe111Ytqzr6YAXNxtIyQcNZQeUilydAPoY63fdfx+oAMoYD6m0TiY63q+J6sw1psvmQaD
TEmY3qDrB/OKnB/GQ5Y8CyU0JFd3NDN1HKmhZvoMDKFYD+czteTLgjE7kBvrnj4dmehX25HC+AaA
+MbCY5Iw2053mQl6Rmaje61ge2rhN4pirwMpp8+DWZdRpD0oAXpTY8qIIqjABX/EQ3+RO4x1wzs+
/iTmByu2rqHZuMa8dX3dZj67X4pJBYzY++a6Vri6Ix9xugxdBgnDgU9GnDJMUQHGN/aI8/MbU02f
5W/Q8WhLZMkD2rtMnN6787W0mFq/N0DgABKm4mTHgwtWxf0VGg+NQoKg8XOgKYLXu9Bzwjey1erF
xHPjkTBvRBqXH/2QMDSmweEKnOUWrjQrKiRQYFgPxuE51XKrB0KbqZRRMEP727bebppHSpc7d0vI
/pmJlYqnm3iPMIc7/yd+I7d1zNUJ6AHL/VHTnQ/Dqbkir1Ym13QEarP03Z7LkQ2TopVVaJoBCvWR
jkbl1JF4OcKviNxkC1lyxKtLRLQfvWBmkpCcxA2B/Ws+HU4k6sCgnryisO2PJ/hVDPrHOT6WGvYl
q6Y7Gab2qtuLuajuPwUAt3eAoXKnDCQnzdb+QnHCfGvw4Qz2Zq0amK/r38kYrRij0IqhfzvKIXv3
jj7p4/8le5eZC/YsQeIZ9DAsaCnfj55X38/7jc+0IpwT2b1RiKIWESEuPWszPBFvp7szfQHq2Nmq
pAqd96Kg0mUFZh6PNuC/8vcIF/9Ju6c3ZOuvFqrUH7lqdF9hFHhcELGTtD6dMmxrr2hNBv956ZTw
ba7ZMQg/PeezinHnDwZLn8cGG4thCTjrp7NSGabLxfkMmztVtVM/uLo3yJ2dbkZbjwFCx2/0Llba
TXgbb9VJY1DYumeqxpPtU93uUEC/5JX4y8lLegKohghK1Hq9X3sc/qNnp9t5QoBTraHIsAyc+X/3
BT1VSHAx5YAv6q/8HPq/vZv8UHtZf/CzQpsD6txnRQ//G2BJwcXI0KmPGJlsQ5mLqVtWCCW6vYyt
2E393IwBrQ3XhsOs4mMDEElV93mgIOiNWnVmRWxrmpEsnp5j9XnXtoXgZM/nHzuluR6974QRXZbd
U9gd19KCwd+juGmWQ8TfQ7l29A/YbwuaJRVR1kzGKY3Gsq9SO/22PbV6d4qBu+WiPSnLkF+knHGB
8kwLGoRRNeicR2SpwJulVPi4uDo4JUoo6D6QYQ0YJ+EsYBDMBxSS2dlJ4um7+8ac1qITL12WIpzK
IqomGUPA4/p5a0EZHsWJJZ7Bw3ZOCCZkLv2VGqPqAyAdcnEYWnXs2b3xb/vP56I1ICieMYbGwWUd
xB96o8rdG+b6XKRwchQW6twFWN4HxrUFTbfgJXskkCDszI4NTB0SoAEbiP7SeGPeFKBvE2mP0MSO
Mn3XnqDXS7T8ES9iExBe1jBbMakH5ciljSJ2gyfVyndp0oBrURKA5UgCzcDlDjkMwwBL3BO5EQoM
9CT0X6imPIsWno8p8CdYyQf0xm2RrgPBYYUTFx4oMYrCODt1H1VFvYIelqO88jxRlNQq4djnC2oQ
nMzYbcoQeM55/X9uSOwoCUU+lkrm3y2NE0HnMm3IHWFuYjdl6o28RmuHv85F9mFAZyyKOGjgF5Qt
9ZwmddKkgkhCgAE3bHTdtchKCxZbMlqcqvQLhuCG7ol2HjfOX8wsYZr2F5CVjoEUg0dF/iqT42pE
OjCe/LUyo5NVZg7Az3Kj8vpEnVNShm5L7CCg9k7QsG1OIt5MiM9yfLhB6Mh/N86EvsWaBvD5bysu
muePo6eMvS3/ajoGR5bK9dquJIGL1b21l8Uhe69mEKcBT1NUJX4zlFeVLWUJOckINaT6kpuFaTfv
i80Wcppd66ClwfxFFt9nHzAxLQgBYXjtlYSM30X0xj17/TzQPTyK7vY4OzOVUC9F3272xWA0EbFp
gi+84wp8yY0lPB8vTc6fzWvp+7tmSi0b526+TO7cPTTmSJ0bVKoCsuo17jiBTzRGWWW/zaHYuj2g
EzwaPrL19Fvi/cSzQsjHagayc784TbjDmyElWY5DsqSAgd0H7VSLG5ErR4usUXkg4UclxXpo6LIm
faP/dtGU60dz9xhzbOd4rEWVcAZCINEgIxiKg0QMGwXl30C99bXQJIhf3OsyBFU+cwQI9SvEFHhF
ngBzL7E/g+ZnslPocNvyT8YCz4cwPZTLtpA+8fOBo60iWkFBCeaA57u2+l1o4BTD1Pdwa30cXdUD
EzOSss1AliOmEyZwD+CIjEG8mU6vIL9AUkkOwUHTfUNBQWTDqFmTBtMdziyh+OVGPLumGUlQaWsp
FBQ7iI4tq9kaOAzEFEWFsaDPJpqe5NMOzZ3Sh7nXwFNTKMotsXL9uyzt/4y5ZwdPQfIAVGVT+iUB
bKWu2t5vBKT671tsF11jpCEYfOxK0QK8wu42PnpPGwhKyGjXmAjVfIXNRnmuqow3otM/TSBnlD9v
ARIyFwDTpt+mPpnT3TpGHb2gdnIA7ocS5c/xbl/SmEXRC76WoYejbQ9md2fcHsgBBzuBkt0IpbX1
pDCN7WHZRZacdlMPWVRQmYzlWZx3PqG9yf09dakK7xNApX03nRC8uUE4XbDxVTJgbSnpJtc1zb3U
aaS/XxQibj/NE+UaTvwAiP2gWVsyYjRjWLMr4EwZEsdGYB7DNZri0fbsEYizXNPfEFjajLHQBMbh
4UnTfJ9yVeMVCIf4ta1yaSkpqmtusA34FMviLaa4MzgW+JYUhuWsn/AkHXIgxj/nomwdd76PDPYw
Cb5g6pySWgkuoNzFWqJv4dq7onwMlUup2sfExnVROLCcryY2wYtqzHwIgPibsBuN9UrZp2R4IjkW
tI/o1r5Pv1Fzz1uAhz4PssJDvfobuBUsyu4DZYGC2t2WBnlDiocqfR47SIq3mmJsCZeL9FOB1Zpq
kzF/cZx0rdPucOYqGgq4PfdiySC/StkK1L0Na/sQc3JqAGT3bBbq85pfniqGtnGTE9dYYGmwUSiB
EjYEdQb6LMbuGWxYufPTL2ziVN2kbwPVYhGwboxp1EXLBQJfiMQh1Wi+1b1ETyoWR4iLBH/CJgaq
Ru6WU8uO+IOxJ/ZFC3TWD7QNJMV9gjMzwG8Yp84yLyG6bpYwGAD2nKyRtFM7M+boUK2euhhvwu9V
DnaycaRrvLuNQjEUerG+ylcb3SkQuQ0do/NBUHFQL9x/4wPV5UOo1brrng2TKt/NsMgT1S2o6rjO
eeB2Ok3SD+tvZy26rwiK2nZBeYg4TWbi/4CWiLk9eVORmZ/jtOemIfYipmpQsnF37PVQN7ZKXhKW
MvU1cz3ktHOIIi1m9spOLM1aK5k3cXwx4lSOLuDRpp0jC0gVx1wi62FbJIhMeRlzoNHpyPuwU2/5
kpt1VNqIwdLxqaj9gJkrkZJpy1Zh9mZ/ONuUOj+nk7BP9qGkLVaazYmB6ojuU2HSNmW1LY0+0LRf
9UEh4hL3RmdHZ+aGMSK4F4upr0W0Ii71pGLAMsbUDN6bE4TYyS8bhk49qXcX4UN6drMxBWrUgU8K
DIxLUemkNb16MKOeTWoR9GcWyA8JD312f4Bz5k8tgzpARh6veh3bDNynz2nENyWTW+t7+jW9fetw
HCQJWtsLlZ8Vh5Ec0EftQoU188aID9xgWR884w2E8i3rzeW9C9Vvtf7foo/HQcJ33q5nsDrlemkG
RaRv119F7RvHbcRN4mCzZjquYLTS2qvH4CbWnr4LglS0KrHmvE77mrGo8y36Mlli5vkCtCwr7/Di
LSLZAQs5tsjnWCMyK2PJZie6lKq2psC3TtNxHlXdCACFr3mbYeIVIn4CsdMMmruxGfRL4xBJfKnb
Hl1ykSr/dOEBMXk/lj9/ucdJhdGqVqkLFdfUfeGmLuR2yfQIwcpb7w/ssK2mDJDSzcSAcxIfqfZ+
mPyu/tNbBybElu1cqeA3i0SU0Stme3t1On52a0TkCI6OuTzeZpOtRh+cMb/7W8j5mYYZoZ0Ibpsg
EJ6uSToSqbv6b2w86lZn47ioagP5GjrHJJbtrl3327QCrc9yl7ZnXV0CxZEGAVpXZEon5Kq09stg
ZktmyKMe099LYSiM6sy2wCoeC/xbHAP5YHsbQ4G1Uw3/ZpDu+FPru9IF+xEZVmzpuLHZnEwsmrSx
uhORIDjNkL6VCOFfGZAor8h1KLUo/gHislVoKQXLhwSdTJLHYm0j1NTiWoKj8TVPp6MLEVdUgQF/
QlT8cLuceQT3EoyyuJ034gwzO/wsC3Ma5emDyz5ux9R4DuCOoRhvecaimVkwTHoy1t+RTzc5waXI
1MmUbjC1cUz0gNgJknPFYE3X+MD6QGdA7n4Jcav4aLpeTlCnUElV5D/f2CF6/qw4xmXUkW9Vh0L5
QMtJ5/4B1htNSaf4YEo5LyzSLIAUNWNrGmUTlCvtQVdFomcKfgw0FzNLdDcGIXpZMjg+OjwIXVGM
kVtYv6cT+lUxzy+Cch/ce3M/mWoxIg1OPK7IZAQ3jEJycmtuoJOnozv2JH4dYwXPWJZKmjzCyKEP
K3uPsEqU2q+pGxpm/ODdScjVZxhGyxztJj3S932rEFD7ozOml5bU+dXQV7GzVTEz/dq/fQFnY1cS
y97T1TDhPQy+xq1O39FihzksqN6bLoNJp3G2v+sRHiXrgkV6jl+BRMEqnVuPuEj1PNknyIchLZ9S
zuJs5wgEW9ymlQexRygJPUH3doWlqSni8hJtmVUCZPFLHF6bJ2DLjK3pYcZpHrBSJcZ2Z2yUh+je
1Xa2rBQcsnRerED9KY11c5RP7+U8S7mQ3VgS96N2twHTWRUvd/go5Jpyqndt2YvIS17geVWnckom
lA/rhzW4oVWBqKpl2Phd8PQkgu6ANQH6fafFozq5EpPduXg9gjWQUEUfY0kkrgZrtAuDzfGpwwan
eQ6254lmilJ9n4EX11y/YG7xgWZ8rKJ4camBIuNvQaK+joVTCorJiTnXL+Cv+Yte1cEbvEXsv/Mr
d674QbD2GMgg6lMY6VnfQuK+MAzy7KX3nxZp7BodKl+R5L42iH3G1ZvVGJL4S4j3cepDiwbivlBK
pOo1WRAe1mrCOFLOxETtzEPbTYIrsjGSviy5Oy14RYYUVTakJR856IpxmRiOpxeNTl5e6GKEVfjN
Jx2xuatEopDIgGI9HiFmqBIs151VHvq7IVzB66QFkFLVF7sTwa+w4QSEMsU2nNlThYhRSxv+kVC5
GCu9lOqQwujFRSrig+cjKCX1ToWsCL91mvT0lD0Z5uoPkvEL/pEGjhUYEa519bRgojOyCgMMxxm1
LleYu6uFFeJV6EFoQbH7Glrm14s7oPlaTFj1RHqp535RGUCH5PZk0eCb+ORzvLZ2NWaArD/eHcbC
Et7kKu6eKSvYhyYLS0F6iM+duUWIalC9nS0YH1emTuzOBsa0jumTI4338G7xnfYWEcchzy8mMDNv
54hSYPye9AsJsY7SuB4C21ONgUBuu9V0+1TmrW0OQG1pGxQs9MPE9oyQynCsfJ3TIqqs2Xn2/2J0
FiwkpyCApk2zpl/ZmB0DcrY790asur70rktyifBE4gk+jIN4/nalqw9UgqwFUOabNhb0qkFAn22K
SwrcOTAuGa5f5QFtamwspAVDbLbOeBGfW4+nWOpvHp/q2s3+YRZjKsUm8YBMkVOztFzVzmxnv+ID
VoZ6nMGZLXWiWrqpMceuma9iiUfA1iyWvp43pDdwCt1X/AgNLsaLcpSW3P/Yhuy329CuW20zJLAh
5VGqjY8+CozWdxB+x+vU7SmkBZhlrT9tDpSZQJ2XWNHJ7K1AsRjsfc3cc2XX0V+pqEpfk/DJVCSu
PLu+PEHJgP+45GMQGg6tqPPFJA/A0YTzdrnw3b2uR4PwGGiH7PiRqbQTzEzrWDmsLM8MqerNSFjh
iMadjkJZYDDimMtnbBhCeTN/BDqZWz66AqJAnqErKd4TmwbjH9dg304Z2cPyAqFoY7t9tzdVdecf
bPdMQ5Xsp0Z3MdWksRthGWXy4YAxmiAFByMxpX6BLBfRxhJ9FGhfebbn378umeAAEgOgS57NNpz/
pr5Gai9aT40Jpcfg4L05VjaF0DdaFI9ECT5eu7GBCH20g9SqT5caDffb/OWdOqgYdHic4XYXKQBy
BM92VtdVlxi8ZzWEOc74mQVljXd6eY3XRll4vKcB3z1bqL71D5Gukzk3uOfq6ecDJ3WOsQmWwrBG
XiUrS3RMm+/KZ7PAOP3ArCAuyHyU3MsC8cyik8/symkWHe64yWorTMC29sQfUCytd2QCB77X7qDb
qDwj7QS9pNJxU3hhJf83LpiP9eqg//xt18BsQF2mUk8gIuO+TrcWekIRt4BRzZJDQPk8rocXpbol
5Qv3B7vyiszvrMoszygOrEVtdSwksXuzkTVidmMJ0bAAxNXU2SYgjPaG3ju9q/vjmMPSmWtl9out
iSNI5ShJ5VOGUEiaxgWRnYyKaI0vRdqHlqu/lCkiqmV3a73uTnsb2uRldS/Upf2uTcwJYFjCHqEd
Hb6w63zibM8a8bULJ1PsGYoL6/fmj6UZ+/ON736VixS4zadnNWn3LKdH5eYWEtCYlIJ8gguOCJwa
Fg51C9go3ewYOqA6HuAB7rfIvzq47GK+ZyVKzQB+SN/wGzJyrPuBGzWBYgF+Gwk/dHP26OJJc5jH
dwbt1RmFDY0W0sT5SKCKVeAsPU2pyb5iIsrhRXvseknQvAwX4RB/GameZ2AN+UeXVlpbZ2fsqsx2
CfVb65RmeBFUjy9xWIbzMSCqwj/g4nVXfY/MMFVNhswTT9VYbT9DrVWZJvYxiCpjQ2rb00KZ4So7
NQD8yoQa6YeJYIE4smXmi8IeS2BGPSWyx07z4YVDUx9zy4T7W5RL93WFOQbIeh5k5yPvqBobMogT
OICBrDptv0c9MbgeeQfY2fwcRXFpfrAn20akTjBuGe70mcncmMnwvmMtqgHsY+g5H5gtXQvFJyHd
D/FvlJuVnbKb9QFB28rSlJem2dYF6tOHlqsqDaL3ALhlb5K2/Redl4DjFsRjBbQR6bpGB+xQnaB0
5sFq0Ogjo/9BayKVNpRiu8C43bXDQQ5d+8H82T3SStGcrE/Q1j1s2xjvCQ2CmzFTRZJ1NNg4U5vi
veHyfewqCR0ZOMNNv7XSjSsEfz1OBpzNTZ7Woc0Tf2Ov0rgb8GSjWBMGG5hGub+mZIyCN/GrbYRr
gkYKsKnRmPyUog/lFIws7MgqAR/zway7VMWhYJlJbMTWGreCVb0I+NLUP/+/DwduCbkRR22od0PW
//0vLvC5qxf2H46nkpFr1gmLebfmgn9fPuwNUgCWzorYw+Qv3qI/tc8uD2cjAN5L0crY/Qbn+gkq
mre4l7w90nO6hKmqVPYdsbbBcUZkzPwMKlGwTt7TKQ1CnjlLvhbc8Zcie8fXm9WlJ1/1MUzsk93F
sSXUMm6DKOGp1+0/jE0jrm3C+9rvK2VsWmgCPL9x+bcDKDiXKEsSvevq3a2b/RNCOM7IKOPjGkVJ
Gg3i80b/Zyx7au+q7R2LvL8yAqjKm/q0TXIyutucxgD8FcLbKN5udbdIw4dub9B+hYzpr5Jy/6qk
hBr/kiC4THSbrVzNQPzzV5hbI+B0AX4Kg+Wi/b8/hIHiB9PoyjIaah/8VcXHpyXadK5BTjVs6sI3
cMqEHq+42TTIRVBbfNTLIW5J2pTM/veHwQRc9jGyK33eSPd+oeBJWmjfMEOAFrn9SMSWIgi82xzU
WbQuttAHqPB6ZGw+3B2vpJsXDEDOuNI1Yds7SUKg3pm/fm/2fE9E8Ept7WQY6GbZeDmHmrPUwraQ
boDP/hg4Zlv2+Amb8Wugznj4c8t7dH5HxLZIRsXzUdzEGtPO6rvbMjl1k3rYFNWK7GKt0lthH8XO
4bnXyeM5dnGBhkDj5FkiwyO82jhCTjetpJxdPfrc00QlPAFBKDiQhbdNFPKvwbCE3JCM5RD3oGg6
Sg4PS4QOY0Ru7KXeaoDswkoF7dF3cS2YGOiAWuGRV2Asm0KJHwDm4T2p1Jut/TKuPbvcAqx4cvWq
HDEYsWojyEaHxtlYo7XX/zW+MhoGAmA5KbozX140pmBMoQ84CiIxNg0Z1RPndy3oAqQVjt2hgzQh
uE1jaOm3Rconr6EYA+elA1EDKsis1PKR93Scpu5YRP5H6SOt5OmOpwHZIjPK+D2Bm7+fcqk6OGSl
TiP8/TkLQXo+8fq1CMQldgjRowVG/AKqxNceu6dYN4JoYGnGsVuZRutIBOj7QvAUQHK9aDq+bmmD
xq+07It1B2K5AB632xW6q4fBBQhbgJBMuN3XGwIUQdMoVvLPusdVn4uTsPYDJKI4GZokPLxlEPJU
9YqgocvR77Hr6zpyZkIytLDLjq/BJHI/ZK+y7y1Hl1iAVzG5Uo/OIv7Nar08CYCH9pT9tZ9NCwjX
KNx4Y+qsMflnnnxF1d63VBAByOSFzngig527Um3srCctnEp4eNg/ZPMpCeUA7rAhIBiYQH+4PA9H
YxHE8fN70oNguj5kUKnRwSY/W5VBy1wCZgkv5/SqVv5NDRwbFOhjc+Epsc6EqK310jCYLJrIubbN
ynJVhUTDKKNw7CsC+1FurRlvkqRWoF/9cnFeCQ+f9u8npZ2GyQ/vlv5WgI32j1XzCyo2x6SKYkrL
xeJigZstPpVcBz7B2OOQvaXng6t7ymKKHdkDypWOv5HlrXahv0vRv9GiDoibotSr549L5r78m4//
DUVE5qwbRFERHzk5nmQyxngSPc/CqC5JWwyyf2iNUwZY0NIQ9CMUom624U+9LbXO3sNfyJ6FwwIO
bTRZomCbrcfDpCWpPIiIyIS//Xx1uwjHlihnENRVajquZ+OzjEWCbgIDeo82Ed/lW+Wq6ynJbRAD
HQMf+9TlgT61I8aDIjk0L4QFsVRS5JKTYsuI31zus042YIp702Ip5ze0arTVuzM4rNLZ4F0SLDEG
PiQx++ifKUg+HssZn4LEl2QP/MWAr/Qr6WRCr6rxQ5zIn0CXATZXxg5Q/rHhRe1SB26nXaVW1GCw
X8WgZB1vhh/PlX14/4vqfxFtbfKhWzSG4YycvxhyElgOoB/IYQe1HznQ5bVcMov7hwUZj7oLfcTf
zYkUBsMRyoBK5HADzHOgUODct/k1TM92AogZQUVmetyaEnMPlgUnkO4HWg6b8Zx0vAXJ22nJXH9N
U49n8stcAbsxAxEYQ9DYmzoVSnMcZytz928VsaVB4kCPsdGoJ3+06r0fe3wi2qiXZYcDXmLsxOMH
MeYbGXLGRrDVeou6szmbqdkMqWdQHCdmA1f/tk05LotDd6f1jiaKJgVsTce43JBEQHTBbMGI49lZ
Tw+MKWLWUjOCBtDE+F4eSWu5B86zUJxC4smj72qmhMD0QBcZF8vy5+EfMl4Ra7RJJIoTHbiNpbPZ
qEm7TJ/hEN9Tgwi5Kils79Pe56guSbSFWD4KTIh9ciWtFZzzG3FVpCSvI0dYZuZXAn9cw/ZfAp1X
p2BWZ1IPDAUK17vj93zeHxQIK7WcHE3J76eYnGdmCIXNpYi+YEGAlhPbp8d+mvmZAUNoi7n6bKIZ
vpDjxRzHQ5VaI7xoPjEaFj+1uqX8YTexYT4uNksfiQ+CvZRHd5SRfg0otEjm6ZM9oU4Yt5BvavzP
7m0BJdimNCyRDHNv9HZfs+sFQFMBzw5q+9nYPG37OCA6W2EBJww0LEFJVFy/3NgyonOzwlq5h4Ob
HfLCukirIFTHdoGN9QkvADvVgh7F7JLs6WMBm6tKSPIYqzdMw9f7cCz9mPYhPsIeWyw5EPCPIUOt
5o4VxY7Fid0f2b9B/D8tUhvBO4oM5+gjRSdNHHXVm5rqhKbwKqanxHvMYZka70+trge8VhcVViIV
NkLzKF9/ggoeFdjID0pNqP1h2l1H8bPpUESUA7v7YPX8jp0l3IlRJdp7jfQrkvfkJYq5QlEIV5UA
CAuLaxTa4pqcIKIfEP7okZ9DdRjXvDV1ltwvNDKsBUeXZbSJJNrHVgy82MiAykRa7y1sRD9nYCbg
Lsw+YDdW5vQDJGJq2i1mftatTk6+2TW3vBccBorrxF9Ga4Ks+Tjc9R1RePzycBPS9TKK++yT/HAH
9gwj/Pun2AEN6c7qH461HP8TRBHBmXq6EYP7kRF2vmwicno9H4fV1t/GpNLaPzMNWy1qJgdZ/Z4W
yAvWR6LC4N9B246LclAmmavCtrbY0TjQoKbP18oF9wrg7BoXP8vwoYQ5UnJ9bEMPoaPUxGvOL5zR
NMebVoUMGBpogf4lvzLWk+EJIn64Gdo2Fmn/s9NJ2325UZNBbPXTl15frEj/lG3j7i0m+9RReZTn
xd+uJnvRlWMJD5enr7BykvtNpg6NrG5ND0dLOdeBeQcc+pJq6XJcJZQskX6iLJ2hLz0zldKQxR2p
n8xdC9v32HDF63DFGR4aGfP5vKdGflgydjl7uOBAldykMqh3lclU/ZUwzIaeOvqgATWG2Da0u5oq
0NYS9RUWOIE5ze62WFXjZh4LPkLUVCHFbGiQ0e+2YW11XQVhB1VEYOvAW9RlQ8SZdHqz71pISKLA
Oo0t9NPAP8OVXfraqsifx82zjPTAFLqNbAOJkn16O5k5Rv5QnutEmtm1Ealh2LvbaFIqjOj23vhU
3zvbdgXPyRrc18YTXTbMNENEEjqOU46917kTdYN2mioA/jqvfA33RM85uFhhEFD8axv4quI6lNAq
ZOWM1hqa3yq1hUbHyXUtprcnL13Dd/iYr0pViHiuDGKicF5f4qvIpsKbvBgw59nqByW4zQTV2vcv
HDhyUi2SLjtqoKmJmFHCLBCkRG9O1ksTbX0GseJG7xOAIai15WnttkWzPbY5QbWa2QUQVX270r9E
VQ08mWbyQ/TDIiNU53Ulw7W5RKIzsWYjWyw+7eFC/5pMAGfX/iAXN0gweXz+7p91V/BZVdqHuUuO
93gV5n8l3KY13PwMZUdptjhxHdfrItp2oEL1XE5VlKu2zrNIegZ78CrC8pY8hSOBxEOMmN5prEMG
/qWPPP4mqLHhJYQ3dxni6sQ2m+nt6eu6tF+cP35mW6Q/iKejHGomBCHC18CJ/cafwtLPH6ZBP/aH
QYJnWM9DNgORBcqScuHo1M9GxodARpHaZpkEAxqiyyYN6E7vdTjufBzAzIhr22diWj9KVX+Fe2EX
OW33pMl9oJXUOMiyujuBFeZ2kpenP5dn3pU1sm2h7Yh/gltkT7FKFjzFrDRlCVItzN6YUlPA/vBS
uFHldRdhWSqZK8C+azdyI9WOmKT/k8F0Q5186t8ik/g8M+kqL2nFL8d9HCce9m7GJm1B93CH+MHc
yczmMeclQyCbTrip91TCKChsGxEHmuy6guACtWCc8JeeZwFiYGHUDDx/6YDAm+bpJBTOnA03E7I+
fCnAZydy0cT1IiWtJdLiNbzFj5IRxUNGrtsDLQ7lrtCiVM/jnhcRF6yIg7wbxhljhHdreMYZNnHv
RSeiRlV4FqP47MdgalcQETSkqIQYVWIvzix/DwRibJBGuxImcnjWahzVjDpHYafJ8psAAELe8SjX
RDBzj4Zk0Ro9o40/fnrCMoplbxn+GbETH2GusPGbhIG+IyaJa9Bpww9oj+kQuDS0uVkWOM0db1Th
hHLwu5xffPg1r4SO1qPFfNfzW4PKCnIAvBMYU/O/UTmWkU6bhxdRKC4sqG3v+KX8nw9cMK9+cKVX
Yva3J+lq4EuNJBsVsVXiiFbKteM0Aswh7JpmMUGSa3itTGI6YyYl8WGZwIpSQJ5wOGcdtcvKEt3J
ojQeWK5XqUpOfKJT+FJiAaI4ULLdNcH7ztXtdv7YXL/h+IF6irOfzeaHzHztOpa5HouPsMKvSyAk
vjg95gUVUdXAOAZfq7edwVYk6+FjmUqMJ96pzIuy3YGkROopE1W2tHXyDwTFolw+0Qw+mklpFCoW
2UqxHTpnXD7pNYw8PApVQfzNRTZjrycoYMy3AsqzmHwSGpN5s0cQuDc/guBdZLlAJ7CLW4zsdsKv
vgkbp/28Uu0eAwJtAtdtvZuhGomTK3fJJP1wQnP7GjuCsurUXxidg4kSsnMfLzqZQWoTu06hTYqG
afXZibD8dOy7/i2IG9dyPwNIfouuGA168NlmVHPTAx0jYWwfc+oXYUbPNgNveMW53jCiO3M09m8u
pPef9EmuBpIKSVBufec49i3il0atsSbEVf0Iuxemm2DHqsnONNAZbBwN1c0tWI5vkaVgEila9klr
kf1OEgDq56AZr7ZPL5RXfUWF4C5RoD+XeJZbaAaucr9x4CVLjC7pyrQ8CDb6wKEOhXUEEeLhxCpB
LLvL7af2pDLNq28VOG1fTm5aIr2+IQvPKhodx+o8Shd/REl7my+jApWj22Cuc4oA2R9CloYmCdPA
028US3EbjVE9DdR7ft8t89UsKMTbEBRRi6dI+dVt9gi+aUotfvnSP0bf5SrU+W5Ukc3hcaUp7Zrt
0/R6fnrvfRQhu2fu4fjR6QBb1M3a/UmudPDcq+krhTAYMn2OWuUtq7SXiGwSoQg5syY2qmZOfTht
o20eNPSnlH+VRvjGRdDlw5MCAy/JvYFrsjy1LFhSWvBl4pcFiuyYOyNG2/IQrEYIP11bMPKsyLHm
UFTy/Lk/ebRWw02lkFZVN76Wm+u4NKUcuyJvgruUnQpuDbneKhfabLCaPnj4ljcCwJ3/3yHUYq2N
uLIowI2o6pl9dzHF1nONWFg9DS5gPO6g7w23Kcf65bBfz1QtWq+S236wz1siWF/C74rvDo0mZYOd
7YwZKc1SEnDgsh/pW5O38oJ2Mxs+XsaUiSz60y5B6+AZ1e8/U6vjv1yQNFbI8IHVLhKMMRL1cpVf
c4DkLriHdSkQjQ0Qp2JgiG8quGVeEtpaOC0+DK6faW07Yt9pTjCMpvHhvTscMxXF1h56FuWda+g2
olWcdlAt4OG3T7bFvw/Pahv9rZGXIoVplcEJ9PlMcdwV3fuv+LusJFXTyimz10rxrFjyaHvchTzJ
fFQRdM6VIXFVlp7BQeYUNFmrpqaJYZeS1L9zoJF1QU10Cs6lsaXqGbZS96rLIbGTHf3flWpTp8+F
dPiwegHe5r9SebJyK9mOjocyNK6gmpw8T5roO2Mzyp2xzd+GOXO6h1Vcy7dLWf9vERhDLco5kO2h
Q0tGYnbkGwHBJUSN15jCbuTbtcI4Ioyc6mrxZpK7g3TU21L7A4bi7VJOHmA04SecCjlxlNF2WwYZ
VyBrA8CwTwthtDfmcHAU4Zpwk5LT2KOB4/W4ATBlVb+5k8IsdcmbQDmYc4/jSEUgwDy2SlAkHngl
3l7vQeQ9g+xP6ct/Tn7rPSjsWEPAkB89HJlNyvJFL6OEX45luChvqD20rkhzr+VnAqXdrZd31tBd
wi08XvZ0mvA7Y3Sbmj/tsQPK8grNcUV2BxmAvD8d9J9A6gAuok6QnVziH8vNitVxLMK4UP6FE+nx
NtGjk4MLUP5SzgrVi8V142o7X9Ei5un22n9nKLHsvsIyzuld1WluWO2nYOJxQo3KGnVWXbbqjgOQ
bsLDNjzlfFVrjcVeQOrOp9OaCfteJlIJuXpc/I10xpr26iine38twRjPQRTfQMMj+lcBomi7d3sN
aMDj5ws/hSqZQF2HJZMMuXqPcASZnTdSqt6O3zpcFczkOw75LdcnTozOyysX21i9cKj5cVnErPEj
3xpc/KKmf+ZxdvgNBSs/X5Gbzae3hpm0grsdIqSWBvJbb9Tz0p6skb/flrCTMXVPeql4M1/uebCP
btxhtnjNCTrO0D8QlBe0ebjCBMRERH7uTgJgWCreKHurD3uJ2c2Omyc/cOFHo/AY7vPtQx/ZQ5hR
EQuPA8jfcgLqJDeTAmO1P39cZoTEvkorcNPaPokmpMQso66Lj5Ar2J2tJJC/+SkiwSqCY+CEDQAq
hspQW4Hmlm4y+4d9n96MIpQn2lkhUzs6A6YbEy3uTlFM7tP8/HyWh+ZpsgOP8260KmhcB6s9f72T
xlVjVV9qLvSjFIF3G6QR14HA7nxZ1NMbLYUWklMuuUy0VcfEMX9SlzWi717LD+C1sk8LmVC0ETWv
pglKNaPDX1gl1hjNOFH8fe8hZlVQBFZxBfN93ZQGQ9viYsgHbQJfmSCPJIvPjTAVx1y2DT22Rrjr
frqP5YuopbIyoa3opwUHVa17otriNvKL5LLJ5ckJ05t+ebdm/nvhIosG9ycv1MiW3Wy7AOstr/vc
aUppWuBiGI4qAZYsontD+3uXa/cy0RzY1NXmrXlhfidwJ+3lJ9R5hizKpd+SqgLAhexHehK5aJ1u
RqLS313q0eDvFnRcfkKw5E6sFg8fPlKifnxcBaRw0hZjvmgLuMIbMwVpmS8sJYKQPS7DHNVKuIU2
Mgei3prFxsKOWO3i8Juz3EM2dLrbvOg3lsR5ClsIJ7kOOSNQvaDpRv+oQQtXCr/lPtYBxL1ZyMFM
o0eRa6GvMRW5mDjs6xhVNHYNkxc52t5eSpWJLX3ZilXYxa0nS8v50rUKqvybdT4KYx9HrRwzMstc
WFzcqHo7ZefsiA2qcioHlhnA4lFiE3RInnPaZQu+OOCYL/kuw+Xg63a7f7lhkwU+FLsDFTSdpk7q
s0HbfpXfAD9VAMR3RvU2f9/0ON4EQIB/kxSZQK9v2px357vWgvtI25neyMJJ0dGRk1KuiRvKSIl7
/H1rGHwR0kfjQS2kafIMDkXg1Xf5E1y0/NxTZPf/qBb80M679jfxNYe9Sq38LtUpqaAdrJ8UeR5C
T4B4b80rOnPxYx1k8Bn2n5o+/1BKTf5BIdbtr+G71Ggo2i9Hj2VPfdYA3l7hYLn4vrD3PHIwl8WB
BpCfK2BgLnKGK6cCygdR9bzOrtEVZWP1wEgcmFjeADY2jCbj5MGA+gkQvGsqzZdRGe1q8fjXf0hO
G9DhUj7GdcPdaVZ8P8GIE+koEOXGoxqyfbq+fvX5NOvNajM/jtFSfDWdhYXztkNrsW44A66jdkI/
O9ZWPiWFeMkUSRkI2g3QSMQ51x0Hxa+Q4bGOAmh3973LPz/bIQeubgjFOGd6n0d8zgrYilY6vyFO
uDW5nYr9oiOgedXrH9g+ODCMMomTfCuBXyzV71WrzFUweAHDztySKJW+F1wceBrtqiIfIUK2TH3b
pOlf9KQNqUSXM9v5F/GVYB5N1s0tVneAUBaA1ILvF/lMpwI7BBFu1Td0zzTGiROVDszau1DjVFLw
Ivq/2WMyBAq85TQ2TWwd4J7mjCcWkTb5STiV2pf2nWK4baxu5ffPlxWWOlRYQ24tSVNYGBqDrWkd
/5qaIjKZA/8CE7iWo579HbGBvpe+n4LIYmJEcuDOFsBRmmhBXPXd4fscU6zstiXYX4PkR4JRVe9Q
IpCEYTF0kvvYaiMbLdNWuB/XuUdjMCHh6a0JN+BjCFbqOh/a1d2dGIob0LHw4IzRY2wiIynkeiIm
4bIz2tag5jE47lJpioZDPv9nIcc7FmuAVWi5voMMT/K7VCc5/y/YvUfpUrYzaFua+znxAShSCphe
eGP1uwpge16QZ3/MaAw7Uju5Gubq5nCs5AqnO92m89fROp52kleq+32+E4cEkpwaqbl64sO4dJTz
eImbhHUEmZP950riKrAmWpGwx9SYRUkr6NzNOJTLQ+AGw1Lc6yPfjYaKKSMJbtbHkKADOYHN66a6
teCyJZqXJ3PuVNOJcoqkAn/ceC61Yjvnfo7pd7M6YtGpPkqBhR6JkmYauBjfPW0bjDjtfniKNgsL
FDj7C5m8Ct028+abhL9DwjMJ6IECvItX773Y6fYKiLKcwWBebGSm51dDycyeGld/JgzlyLOmBmVw
+/daY3Zal4ntgkPN8+3Dt2CLZpprDZqb5SD/kdZoRACeUGdjMArsim6W6FRElp42/bK0syqqPG2y
XCOVXL67c6C/Zlxiy67VUNpVJacpUoPTzpnUHgmsMOdUVYFISsp0mUFS4qSGrlzT5VlSw+vDsGQb
MmDuaxo2DhEeU4qPDYQEqmwZPKfpDzaPuvsocMBx+gVUQPEfEugYv81yhBzR37zkp01kxXKFI2Y+
H9ncaY6Ef7B2ZDSsJOB/w3rCVvhvshMNnmEdPs/oL3fLNcIevG4TYc5HRj0AcNWSwlYPG2Ggb8IB
cfbnzV/OSFLUqzn+ws1NjUGRi1Bhnbp6S6YPBHhDX3gLT91hWCKKoX01rT9Ttvi7JzSFYegFkP/l
6fl83lOhYx1bO1fByqYLyxybjZO5GnUy0uT1ZEKcN+OaS5V470Z9YYQOTs2hTGjIVmE9Tp5li3/W
8USzTRb2UzPCCJSfEUultvwMTI/egS6zT3PmvKLI0ALVE+7E2eoEJPtiAKKX8WHWddBiaAA5+bJ7
y7kjHk5bwIKHhqjPnSmthAsNTtfxB8gutatW/bp5aEe7jBX/+ZlnuxDa0Gfg9fatLiMOAgzeVI/H
aYtD1xArkj8fYlubzhrAiR7IaXa9RjuQgzD82+vVJdtfuJ24wXHJx3glQipogMdBZRsbtPJsNAl8
pWMZDfrA44s7bmT4oa79hWCExI6FJW312G8lgh6wj3z9beHT4shNvVwziSmh3EpAPzF/YsWq7CsX
H/pKstmvXOmWWQ9S2O4JNUHqvJYryrj2fYEOxZyCogkvEM5d6wDE/cvr8VkKkLbIEjrqegmzaUxa
oi3DjlgTwMXDnqbuEa9Ihb8o5CA5btPQDEXDbJFY6xFZYyZy7DgQLEo8EjGoWjbn6zvgv9hY8b6E
TjhSx/xrIdQdcEnwGs0aDPzUskZFX7gC6NtUEPepMQc9MpALLe2qhCSvjkB5K5VXB3ePCvGsBhQJ
5qq93hJG1R2FPhrCYRWcyyn9600oBRklTSy3uTy2Q6a3fscBj0+QeCPnmt2x9RceEVZcLLhv8p8W
0RMXWGvB/64I5iq+bglJOPFj5/Jo9Iv3OIDB5+O0Wo48Xj6gPsWB6/i/+ZY1ph0WW27PapH1EuJg
LNOms/XoQ1kruJZMwIQkFq70vBieUmFxKrvyB0G+2a+7mYqsUow3vxYlM6dBexdEQi7i66vQb/gd
FW2M5uLTx3/Msa/eIbEhFgoVXci++1mVH+LH0aI2A0aZa0INJGAUirD8pEU3xoEn5nh7cl6ENILH
vg+qv6BJXdjGEbrBgcbS8+A44jcgbBKrAGgaMLlH7H6g9Zw8ZHYEFfO3Kvl5DhJ7g+SGme4pwakA
RFWQ/+j8jb5ZWbioxhaPTEwajUipTMpXBWM8Bsua2GlOYy7zT/7Zsgx70SUS0fmQ0SOzHrlr0UFw
uDYBIMxZC3lsVK6CmX2/CE5yNOvQS5I3dE5ucU3MUovEf5MFTOasE5IQNtD8/fmJrr6YE+N+iC24
l70YZPvxDKZ43sxnj/ewfTRuAbend3qI4JgzFNVAg7mQinpuHGCG6ZUyzfx4MnVtkM6/3ah96ce9
QpK6OptbqDdPcIGJcBajOrWMPofNmh57uNu5tKgHfOHQPzgDCa60BJ9jEGOCEF+GIEhmJwbj9557
sQU0DsIDM5covpo3gtO0IxoPTM13SG3+BugpyDzuDnu1B+osDCXlHSNzbgrybOXpz+zQFdoJNFDh
l2Rm43iYvet5j8y8/Fpe/+L9PPlFmSNTi+L50WhPzuqThouFyNee6uqUFwkjN/8wyqMNPIq/N0hE
yx/1zr2ew2AQ8hj8H7JWnosNoZW7vr2G8G2GatlGNBydLo6f+XGVTiLePa7FwYRI7nqSDnE3oZYQ
9gX/dPTJzJbnhmD3DFW0/5b3Eqi4r3WMapXtgsTpxYshbQeYJ8YBYLgaulKEvCslt2UVc5lXRobH
eYsONFaRiGsCxYofuynliqDp2+DeqHMjTixZHXyS43f7ccO0czhSFfLgSJtDS5/l7fEEqz3RwKD8
xdFbbRmaphf6OnQnzgXf+v6Q4CiEM9f+/mqaKDYCRLjGXIrRHTX2R5jECIJTKPEL7flEvoQwOk+4
AYmftnlHihdQvscPs9W3le/FXQrfxik1ZZKYbU+8XduR2X646QCpKJWb8iOLDKf/zSvLwDDuh5BY
ynaJbEcZicAdHalrVYc/37DFIjpETFWAFPIdwECGhCW/bRI7I8MHpRv9yJi5I3AS6wKE91o1fUS5
1P2a9hmhvfmBuRKUqElymipl4jMZMqd7/0Fd+1BRAYiXEMSWdB3cU1H/q4UyxMH0aVlOkua/c+wR
fUdF3QsQg7w94oNXP1fScDyVei6qREnXxWDSXCySxMpNUHwxBf0Xox7gS39fFgrW7I6l+rJKrVGu
wiB9z45nqpBWbWu8cUFCHGI9twjAiQjWMxDjPesChEhlcRdZOXwuca+4Ct2YtDJOpGZmItUoLSmk
I1XNOQMu9+n4CWuVg2VL0h8aqYT7eseuIz5mVRWCO/E50Jtmt/G4v99sYg+MlJW5wxqS4dC2po5e
nPTdPgLHN/1Z1hC9wXok2guFxjaEuAkxj9hJs2PPFRzm5vLK4tqY4eUi2MP706a4Ku4cj/E8y04b
XwZSv1WsbHgN9O5BoIcC3hz+cbcLbOIpIL3v2DIwyUEX+hsUcS68NTf44b4MvgpmiltJgLd+xOZl
UABposCrlxJyQlmen4oAjW3ba4jHa797G+IItOVdh8vGXl69YMwpYDCsaumFEecPJ6N54d74k/tI
EyjN2t8tEatTZOnCDZXOIqOuMZLjBUsnQXfBpgwfh4ZvZgSX/SHJA8lHKclYX791RbPgR9TuobGk
OoSoxChrM949cBZ7m6ggbxXZ1KN6qTvEcdV8p/y1Mnbq3nk3IT/OvbtE7GmZVpzafdCZunMivrma
aESrVtIwZ7vFnvGZyr1rbkYi31XX/q47nUXA7wL69KYzRLK9E4DdRYbIfQ55hlTpw9gs3RVD6hyU
AfGne6BS7DM7gYMQhcseJi7ZPAOx9ImDNP20aR7S8WXnW+a1juP3LmwrpqSpUuMZF7L5y5aN3M19
VX1Oq4qHwQ5d0rjs53EO0J5j3KPMZ6orcpnvVXAfFTXis1iM0AQR3KhrYLJowscrhw8pr98czwTJ
udp3Kb7Z8uAdc0QKgQ874WeyEt/472whtFY2eVQrKczIX3/bAJ2A8BdLnIrIBUOY5YLzPRTLLd0s
5yo9XViFAuIaB9yHz3h7iKoi62kU/MkaojIwc/wsbdl/t3XtS6FvAVyEaoEDyC8T30PnE2UFakiO
F/EySSHtL8EIgFq/XjnMrlwacBg/FAY7vlvpYUosn2637cJATbo30htJ7OtRFMcwdv+fT3E3L3lk
wRA5aAD/OW/SOByQcrOnQGB7AUMzy+STd2FM6oYg1DdtzM8yOYpFuMJR5jDVc2FoD03ULuZFfS7F
nWEh3ny0YRTMlSOg6aY5UkprXbN3VNmhnA8SmBQPuTHjggnMfGNYXvk3uSQ05jgru7YzimfYEX3c
atRuW6JcyUu5RE6zZyNT8QruHMzjkP5EkOkdYnDh5bCFxwu0lvxgKJdXxcn9j+9jslwR9hRS79Jr
8+yXVkRBGPEq7riTTKV1HFoNWz7AT8ZEQhGSNMlNgDbYIRYRA5wjaUopjBRHKj4ESfTBbglT8H+g
20vrSNLE8dp7fML2S/J707Mvxega9Ef1A4sKs15QHLBwKOAsFkZNENPcBGdG3RLzVmlnAW5M0943
y8nCgNBFJ4wSqLzRVfdM57Zx3IXEGpJe6r1UZrNwkJnOkmtMOh9B/EWpsKzw0nw2vu4LcQjiMI/v
yi1U5fS5ewYoBjOgnu19xiNGI5UPqRgVy3TaZ2XAQxjtrLp7StRC4lYV8zJUor0zPxK/EaFqJleW
qujSA2YjvF6VWlQhBJRD4ZTeuJqccT3J1mvJfC+4K230CI8bdbG26eOBla6/ZQ3qANgRHJWjEYnN
6A5Ee4bi5eMKCXEY8ATjT/kyCUTf7hykPtELMrIsqd45EHkYFO4TBtud0w9S2pw8Zz8yWqdGpTtt
Lqp5Pf9iwActuBE5Kg3zDL5bFxrkpIy9GXq26+XOlByfOyBwGr5auamFP4XDXg+eJKRjSFgc5HjQ
n88+3+tAqJklp03HeHMM34HqkK74vefxtu8ibQIvd7ffXaIK84Btzuv0ratHeqrLv8y20Mof/rWw
nfCrwLlBEuDDqvr+TwYW7pg2c2HN8mvEHLKOQUjoASmIVT4lRWmmWubOCUZPQF3CV1GQpZht9uvj
57kocPsaGyyyQj9xY1YnUciHylbUdARTbHQtaBuoVd8q+Ym1A/MnXUFB2uNmJudXMSfCcwIelSKA
76d66IAUEoUytvrJtmfSqE0DlVJozRkthJEdaTUwlylsiqI1HELya658A2vciqUQ8HciKgAu1VpQ
Ry1ObGaKmhphGUuVYzE+5akACGJ0hJaTXZkDR6dSL8klPFiuMGsImofToAX51l0FIpCVGx3YHz8c
Ml9Cox5WSzBAIwdt3AtCmZ39UB+6BI2NSq8sZ/lB9u4vlfnZMzINEUi6hP7uR7mgIcF0lDEMH8v3
4L3TL02EdSFx366egNEsfcUnWCfJflp4ADggPnJNoCCCAuMUY0M6xqiAnVoYCbJtHTVgQSwUmCb4
1jlr6Uz6j5rnllpXUu+d2mNj8rCJtwapHEOh0qUomQ4LagnBkBeh1Ky2nmvtLWSDNjLhQs8840hE
dIyhsYH0kniTvKodppnyYOOZTGDVCXFbHSc5AYEOK7kdWPyVEbHsutgIummwsDsvX/CibZYbwOt5
4mnuVY7h3YjMdF3hOXgmJDZjkSavOfA3CQTHr7CLWElPERMcgoIPH0MalT7CxliueehMCYULwri2
wwYZy1stjx+QLbR3g7/hsQoVdtWEKC/pSdC/gc382sN+5vO/cMTaGGK0mHODLJbZ2U0sJ+J9A6Tz
rA589g9J3eeV5w2bpmdG1yUVBBJg0egRhp+03lw6KAsKi8GZgufVXo83vH3l7zHbckws7xx2KkIs
1dwlXACA6Nz59zW0k7elbxMUdXJNmM3d7TJH6mXoGQliOtw+x/gDqJVYTJOjengRNOu4Apt02k3F
hweGVt3HdEvGfwZ2cocc6iqVF/jzVTC8dqvpJMIHOndBMNCZOeeGO1ZNvYUu70PnGX0pvRQDiP/D
7ggBO9qV6AnRopbT72shEYNudnAl4VOtBTHX1fJTFu/kwt1oqDpeNH3fq1p0wcsDiu4C3VV+iLtN
UFoKeFWeFb3JXttbbPwxZe4fTBXqekUZhT5t25of73KqVwM8mupsMTz6bHfOZzMVHCvlrcVroyl1
xs8tOoKo+PV42wYB1ciVH4XM6F6e0PDMCzAel3uYaevgLriGNcTXTVWu+saz92SANPMES6rvcmKC
unvtjJM2am8IxQB+1nRcUrr66CCR70IrbSjR239ftxaER2+BeNoivRrmdk4biMNA1bxoMXbSszAS
Q7WdCzQC/1Bfh9PGpCn46vXsxi4QRyvLPWd+aBmG9SOebtO30Tqb3MadPcxeZxfSfKrKA/7/lYtl
dPk1q2OwrwBaj8WBvgs9dEt98t33EpIpJGV8NmqQ7yOQ845z4VFvm/WXFQ1TsZVdgMORpyGakX2v
SyrpCbevmGSbG3CiKHBCbV1eeujUq6Q/UFSigi3vhdT/I91oezNjn43oN1fQFFwHYC6YRTedPtMA
gm/7UtHITMftQ/pjbTukVoVrI+/XDu7KiPyO2Gz7F0aMiC4jFe4vsaEO6mrgfxWAThTM2HZPJbYY
UQXc4kF7N5jZWe4zs0lZS05Qw2G3SXa9+Ez98DY/QfxoFTfIIdo8n9KKeEW1Mmnc8H4pUXZGJM1J
A/rwn7gCk5eLB8TNV4LsofTemFHZ2cE0dv7xyLuk/RyecxTm7U7ZaIuypt6eRVu8wtWqj3irNG9d
xh15ehMDv0Widoyu7Kd3ST9AhyziqDNoBoUUZtpxVInEWvfEknm1x3IBd5BF+/e90AVTuAwe1Flz
f8gUaudImIIpLxem/oT7blRKglW84wXw/ETkciSB8vFY5n/gTdjY7D87UB90SfAFxdD5xrmLNQ1/
xbRg7MA/Kk3UgjlRn3z6H+97xb0Vn0QDsRXmlORMZToV767MtNGhjrvt5fX1+xQLm6FbhBCyrrW+
6++vCtLJq3YyVyR0nnYLb5AWSCWiDFcCKgkGT9hqYvyuDSN57qV0FhhjRoOKiG+DUhYzj1wts6cB
uEXPPd8cftTC92xqmm1cAaOs6MEzT3QP84y4YatrFsf0VTAMszmr4ydprR4GZwrUCDoZ3PeZHLMT
BqaueW0ub3vzIkQa8uVJGpaedhk6I8xPxUwex9SjXZGjyWBnfnX/dZr3QG7X97g/akRo1pL7Pofc
9TYC5N3I5/J/JYWwR1iiqmnOVOgNLrS3hc+v/p0O83A/RYo6qg6A/awBiiS4p5V/o85Tp97vi5Xa
DC9DGtSBmALRB+5GoXEa/5yg1O7kHhB72YDxT+1MbSfOesFJRF1GA7KzhYAZnYRPSeyaG9jasOPB
g+SOoKxYaZRWJtDB3T+kNIhlUbQBRgxa4m5HWD6CKSxHArhDDqoWamZ0CFd8BM1UQp7HfDPjCnIf
ggeOV6Bc3qwIQEgx04Om3yrIJSkV8FaISguLUMynW65f/jmeP5a2ORQmBEsBBoTCTWLiuzC7YZp5
2iS2yx5H6yryWukZvUcFNogxwPSdOxGv/Pg0km18oUoAMxep32dh5uuOGUvSXG3gYPkj1q93vwCC
zxG70ddoCc5WvHDFBA4YSHdFf0jFU1LkOwKLEIkoD9ZjiQvObm6Vyas5/TfZjp0BowI+D9xaXKO2
CvhWgq4RjwdJW5HJUYm3mYQ54XRKJ01+h+VYsq2L+JQmKLrPilI6DdBfdWEtvN3CGjvpP1dCKS6z
tY2gCN0rLkTKUKwJO2bdag0ItoY/ASFU8djsx/ND27NasZOkMu0u4s5kzDb7SWdFUhr+JfK7l92H
gyv1vMapzq5zEjONXVZF9mVaQPFqSTL5mmUZd0qXPhAbIWMrVR080ecg8vW/AICejAYmPJfLw1E7
TZ7qQhvRvRR3ru48lY2mI3kyIjbnkRawlpR+Xr5M+jmWH5ckHkKypHkQ/Q6R6O5lwrwgIBQlT9Tw
mSYQBKr1vZMRattU4FuJtg3j6ThYOy18LRdCHGAsw3FAlgsizq+0DGq813gopH4yYZ8iITJR/bM+
tKB01H5Jm+UIeftTqqX7mrpu+VNR/s43aCPK7fZIZdUieaAIdRXR//nizCQiQ4U0rHJxUnT12IJA
r9ZZ4Mn+gBmrtM66Rnj0Nc8CFe2rYRORiW1ADMVh7eJBxHhKzZRmaWdtJiH7ikUNSsla0hkjN3NS
T5tJngKbow09tG5dMcH1iBRjRf0nJ1z9vTQuHawO74UR42MbX/EewvBIffk9DoJg1psSkOXxLqmz
NATsj0ugjPaVbaN6WwHSna6ugGBoKPH3GGU95p94JjHTSxhCd4y3V+mLBMsq7PgLSxp0m27JmGpy
rpf507/qxpc9Rgo38xygYz7idDze1a3n1+m9fEw7IRB0pSTVNZe9m+mpcgOHYBmvqyISGZW0R17b
zPiD0XYo1/BClnkCesVdq4ERhoNwe7DppzLQtDtrBJok5s8ZCfa4kT/gDuHkQPDT8zFSV/WRElsM
9ExZ9tmXwEOlZa+hMSM1gfzKiKKiqRWqE7vC7l+G8OeoceDQVkYHYl/76xfd0VUKvJjL9h+kGnDZ
tEfhAE3MN85slp9LgXqroizkAzUuneF/zHg/jE+oUA/fNUFTcaY3XOgHbFDSqzBvdCtttR/8Vg9P
3QSAuQQwrnYCwMaRVTvrubeQNio8yfanDHU8YYNPIY0ne09l/q03M9Ozky66nmytF7uOzoCS4I9q
C2Y5SYh2FZnp+hZOfapmJOUBJ0IwZFkgqpvZKrS77rC7sjEqAz9TBHTUAfvLdT8OcB//ybmEzBIr
8Ov+ng/O0YPbFUC/7eZ/bHA1D9eznWn1PP8WwKnq9DnTdXr1lxmHKMfp/cj+eVqN1MCiurkqobe/
Fm8Ip24xP5FY4u57iYFXwfJIS4vGfOZltjGW3aiqDPhdGLcJyo+N9NH14GIvwJHlWUOhAROGdU9O
7uz1Uk/IQ+Vd6QBe1y0p5rNJnL2FoDGVryWOMpcUV0Xp14LKGQtZFn3fX3Js/FNRWaC0OpRgy1rK
hXj87ogjfdJyoxUGLIGZi5xM3rtIuHGmrcMHT3IPLct4mB4MrjuaoSOqsBaH8Gx6ng/fhOgdgNE0
Wap3Rh8Xqe659kfGSBBj55jjbSoRwKg9PRsBedam49FNwXvmJLae8+oYNteqPcanOlYXHGHjfo3J
s/wQPGmQXdj3X3ljMVsE7BcLCHikxMcYzieCPH0vMZoWUiPgJ1S2ehxUbrfw6lxxzEAox9vJcwXp
gcbxvBa0dKBA9l7Htr4bMs4Biua2Kkt6tvjOT9e5+FocF5Q0isX00CEHBlgXeKyHLQmLJnMvZQqM
Hbi3x3OWLSejyZIMXqFtmr04psV0IQifuWV2PQjvPv93BvQBAgV6NL5CZWfXtF4rONnDm+tPiTwx
5+0kHd962zH8KGmlAGLxlz+CYKwLy2JfDiP55kMlNt0Jm4EWy9Q7vST/ET8UQvqCczMcK6vaYW1+
P/oKehn7cTRwYDzw82ptdqE6Ob5qvr2OdEz01Ya6sW0ennym7T6XYAkGh2SjChoyYU1XQebRNLbl
wQg8LyRCPIu/TpJkIoIRg6MeV5Zlb26AG/z3D0Kaaac7HgSqvA7TQmxAs+R1qx5F0jdvYjJFm7Im
inDl9JUbAXlqW+QbMadMCQlnnf2yXv0qCfYoxKhTcOOj1Z5RClnJ55Spdu47YMC9NRLPW73Jih/z
HJJzqwLvIVK8O7vVWiWRMlku/CDGqwRruekzoqKoGt+EO/jf8dLEuQMW80FWcXgoS0JNLeDU7N9J
J/kN4A+1xFWfEEibGrIMASXhuE4FJD5Jj1AlqwSZrRq9fz8iKb1YSgYJOxdVPVNvJYOctWblQdKQ
QbnqT0OwRAjRu/3AWPYzXi/7M10xcklrozMJasIip0otdOK0NrtVYtXMqEfJU/ig8pQKbB4j+oTi
dDBiO4eJcX1jzg7GT+rmfO1So3Wmdl+HKzsclvUKSk8T/KHvZtIuWcrKlHq61DbRqpM5+PXkaHVF
W/J5QUxvTN80c2eb4PqRUtSBUUsJgbG9WEA4VdbXWTNvW8/43xRixv0xu+neYXXa95eWVSRHUjAA
cbgiWIRJRNFRCSE9+72aojgL+YnucgqcgWheF54udAXUnlnklpm+gT3JiN2aKSPi68YTc0e3J6Hy
bdEUIbC+2Ze2nb7KW5sywJWJ0SYnp7WE053drd0PJ3I30XZsqtHrf4PO7ZOe9yejY2wk6Z5NVmq0
yJWSsrgzATY5znYqSLjYXYHMGf6mD0+QJgzCm093C8wQhyFjuU7LJNE/lS9gbezZ1vkem8X6izx0
amYSXt9W7H4ithg7JBlMVWXI4WI3csjGKFKsoa1n/Xl6/VOcL8dRqZuaFvjYsfCE+DsLtJ4WMFTP
4Rb8uvCARj/WrvLhi6TISNtdKF5qvxK1UWkIHfEurzGgHR2q7CwAK+elB5iY0P2llPIAtYy1WRds
SUabtHUDpUiGJUdjg/+YWw196IHzp33RejrRlE8yvxe3SMH7nNFaeH+ggT+Z65LhpTeIBtckG+uW
xgLErRYJPOZ53rzGmJ1Ah0zFNCLnFaKZFQ6MYWi8RDXOP/YlNV0MymW7DO75LZVoHiOi0vnUMp1d
YBZ+9Yrra09tAvUxc/qGr7L7KuPXXcqGZzb9OTT6manPtYLkniOolg1wlFBFyTOSFq+mauv5TO4B
bEVOmrsTbBFf+mwAlBLzJ0tS+cDwueD5sTNzG0IoKbK8my9BII66yoccvco07As8ZK4duRbbAOle
GcEoxZk5K7eoUlmp5w0D3natW0QHKkGlu3AtGIHQt157J36HRQRGdvIoySJwQA97X4BfPkQ5UAys
cfFCcwSuETAOQPsL1ZtbMLUFNX2CZEgV+YLQwCdgSHLE4KNBoWNKYVDdwFXAspcuVnW/e+i5vBBv
uB9gHzudDGfk8WqjGGMPbI2kJv7EpxstGrPNAfPOjCNQmDb8yOB+lDUTorqsIZEhkYSxICS1HSml
bStoKXE8QC/LB14g8uuypALGIThwsvmxp0luJS4VM+cfloq52y3RsRgwjm/uRgF4K/wN4OOFftST
vXzYx/QJm+FLK4LjtGD8lmJJBX/XJ3kyJrviBYSPOeqnAftt8maZKJGOrVQjOUXQCifNzSCiHND3
Lf/HxaKZzq8HfD+WmxbrMjTvchkvsVkmX4e5MIO/W/MT5qRx8F4N8JHVdBGCzYjhWTHV73FoGd8L
HTjXTEnfYcZSA1Ji7FEzavtXCsJ6CDFitC6GR+XxO6uJqe9ez2bjmePZEhkfxfkbbVTfiiijh5BM
2EtlSigNtv5CSIIC3LRNIWptMwtoftMydfEe3JrfxPjmWc230G+RZah/hdLnge/j5TjXKPk4ArJs
zN25L5AE5TvHkmEkUFpmhEdRHXaPYQ5/NoP5/Hlw7LzhFlPm+5mPZK7VxsTXdwlgD+zLq2XxtNYl
hqZddAd3MAElePRQ2kzhI27eKZSjRbyWODfroGbCqjNr3ymScIe5mgzxfjl2iPEZWQcoyJSllWwI
u5ol8JZPyodmpiyH46DOjtML7gHew9+m7F/Fdz2/TjZr/6VGuYvOAc8RPYbZhIFoWHmL80d1oOfW
aYFJPhC563Q0whsYJ7P09EWYspIu3+On5Pft+XZ+ERjRoocvTYbG3SmqMnci6tL97XmPivxHB4TB
aHYxYus0HbvJ3kKRWjXjIVecRFMt0vviyifNm8TPwr6itCsjv49dUKzZ5zuc+LXQQdL2oCdh1/dm
YFp9I4p9lGNlzNtAwGs3Mr+X8l+6ByzkzS9qQ7c7DpYc1+9YG5HzLDfSqwdzEZQoahZzXHt67SMf
oHIWJcyDn9lT9vB/RvpmulBIElS0eBS8HupjmSobNWorDjQGElvZsH8RmydARwrH2t2MRE+l611c
6CbEDs1kDl5HR9ICiMBaDcwbxZqyeTJRKAeVviRv6K4olueuaV+dC59w8LLj+iu0JcRzgJLEG/PV
TL45m2dWbk84LhY2ICtwpaUuNq4fI3UtWFBMdJmA1RdnF6k7A7n2xFJ4fFlR+ye49vXB0q2XkwPo
c/AJQZK1W7mPx+AVJjvruMLu/STTneh2iYf9NK/jX6/HJRd97xuEwPcCPn++tAMxbv1qQ3s0flMj
CZc2YTf4T5Hs3CbCh+IX9b2yAxPTaD9bfUNbIWC9bbqU8Cuk7QXHbQ5fsP0Gam7/jDn17ePSkdyO
HBi5oxLZCMUtSWJxU6EYZpmW7UgFHyOtEBav/iI2LHYC8pJahwGc8BRI+Bd2gcIlbqR1ZzugtgS/
AQsgrzYPii+81ExsyrfHXKDBShnwviSjet+Z2gGtc28qoNZi1vszJXLvSpN9iBADULY4A/Ux1UYs
KsXlmMVURfG1eaP2B/lWNN9IVD2SwH2VZZGicU3RXZEjfMtolriChym77KO1rIQJfNcS7XHWRIGP
OHcHru1+sL2IfoHxx1GLmJfhPpXoCUMqku7CIEENhKe4L3KVxlkEFUJ1rirkc1QF3W2yZWwNDEqM
+5AZYFVGgpW4RIoHI0FAGjbfggjK1GEN78mW95JeqpVx/fTRnILcoQskLi6moXshxh9hbIoX5It0
vhvJ9j61X68lTWK2cX0I1S0Dn2i9w80/mosrnrbDE8xP/0aT5ET/InMTZawfP5n0W8X1i3ezNT9Z
SurNYMBj6ppLTYZjrS7gCCqpIUleTYz7lUJRi5dTBvhrjLmMB4F/OS1VnXFWGbiRDxg77h8vA1qQ
dw3w4ya0e5qra4AA8+ui0ohF07UZVwpQ54mGKLNuiyKQ7q5zM17QU+5xon2BjwcQTvsNtmfrkyQz
BkNmNMB1SQXQUF4OeWQjjrgKAbfmxsvyU+vWPSdpzRAgsPfD/ZvcVuLkm1ZG8bc14IGiyZYFQDvA
jMDQBcymFmp04bHqB4k22kOmBK8hhf75aGQpy/JWM+6GSsdpiSGsdh0iKbX0xW3fWQmnEdp5Oi6/
AKd+MB1QBhRqbxL/HhC/sFLtWzB61Y0qX81r0axmDQK4FxJgsjsCRRvXNfJApP1yKt/ig0gC8XRB
2prcPj8vld+FUlJs3M6TcbUNXQyksN9a0SN9Tf+IywelGAIUMlt6hEt5BehDrxmpAkHRBdSaavHf
zcar1kpmULpnDa/AXbvROZYAc06dhgJyV7c+NPAuM1eOlgSMC5kbqqilJ0CZoxSLmIKcDxHJSfk4
TfaWnpgIs7jVMUhI5OSsRUwmyNQUDi8kIRp0QTVVcWAGA0vPjH7JVMqy5K7/Bhe5qPxcGG6vWJ5+
tOXfX6IGRPNtHwsdSauxmKGUN0XoUWuA2jZNShR8BZrSB226qtsDKZCZD0MccNfP7KOJcz2dlOXJ
JQ8Rx8+skVMKJa7NXO1lF86kSwDQOZeujUZXib2BvLrfvn3GLiyOJotnZsch+tC1268P7/U4B5Sb
Pb8k1dbw9zjNtNclT2QhhV1YT4OFooe33enKpnzeFqrZ1ElDEq4KfM8mMPzRzxB3T5HiR8AGnuQB
AwDRr2Xy9EsZ5pN9xXRSPw1CQ00oSmL/tKvY8U7WehiWvyNOXQUSIJ+2vLm6d4VcIpNTE6z32PbM
H/qSf9k4FHe7KJ9iM7KFzfGAncJTIG4EDuFqr/p+rb/aYwbOZp4cnKYLMT/no0oea3OBa7HGy3bX
HmGHL5ZU9k0jsCO/1AxMnC4FDVaHyCaVMLaw+gtlBJ2Tn41+dZmQh0NMyqQSodSLSuiELstJv19n
2s8WjMHxGMmYghkiFofMOcJx8cCEreQTjwAus1lj8M+Gy+8F8I7hUVoHt/E6v9ZD6TkUCth33pkI
FK1JxNcvKpCOBK8YYspVU4Pw6yzvanAwPNFMqqtIzn4AFeXykgKem9Jx3J25Ngc5/0ECoDo8QEuM
i7N4MURQjO+s5zNPXrgIVBfuVPxj5HndKSwPZJ+vLEgrsyCe37fgqDW1oxTcWiATGlOGAKEayy6T
29iBSAhwJyYzGEBwrMO5V7D0QKQ1sufQxggbrcA5z4UD9TWcxqorUBCYDG2oCiS9++91jKIEjNwW
E72v+hwQiOCyv+nhXd5YnbWbTzR7WKtGgkQkjOgGByLD4kFENj3wVEP2c7jUNYtfw3o/xjIMeJhK
F9QbHstOH4ymgjh3N2pZjOkmeBDPrtoqNEVJTKecTZXoQI6PMDACLS6beNJjTcZGvpAlCBLCuTKl
hPfu/riQ1C11y+ODYAHqKKtcNa/RLOA2EchHdE4cHWBJdghWrZPqTQj3OpOYVq4bsjxjqF0BHlpf
M9bxKoHWwbbvgjlr7UknYn3NK8FWBYli8/dL2P/fGuvVGtyaY4/50+YmgIR2fHBU4NnF1kv4ICo9
rZZewsRPf4mPOn77HNBiz3UdBoWVt+of2lGzu/RdIfO2ff/1retNaLwlUpEKLbOWvBhpH9QaLddM
AwxSTUxUbrYbpa99W7IcW2NbyFK7NGEiEZdA9Z9fiJ8zfzBGXE1UcU0VVvmk2gRWxsnUsCu0urIl
1udLVawUDKsG/djM7YwASBXeZYDKgHpwjlQSugOvd9R+TM9aDMTxauEJOtILXUjxod3wzUtTfqz1
iKqLsAchM7//3hJO/ZMglKtqpKV/lX9mPbZtqg9qXr7e4fJb7T+cBrYQ81+Uw7oGP5+KI8Ata97/
q9UTbysJTTS1txetgM4M6fJFl7ZbYoKj9Sd++EJxc+tvRXi1rdRcKsTwz27f//DZlAfJ0CpPaINf
hyDbfODQrnVgDG6qGEFA571fEw9J6kuEQuNUc66brwccu9toalK17OW6bPYSKVr6uHK8KPD6N4Sr
qay4s4bJ6bAwg8dr2WUFgaIqFDfd/6VJ36DaijvdzmulLzkhfSGA8zBVILuqdGjFt3XLTykiAIrB
hl1+FQ6hdvMb7LKZ1C5tsJy7f8lOwbEnvdbwingT0lE3c2sh8VoRqKWrdYN7bJG+yyfHp6GqmF4+
qB3ICmNXhoPzWFWxxTQsvpfdWeC9bSNuQw17gX1nWPrtgGCGnI2+SYWn7g3Z0xvfjNOVu/P7D6rN
hQggiTvgrcBU++DzYu9AMtzZ0o6lA/d77CNKa0FPf/RapJya6Bl6mRCg3aVYKAk27TU4PAZpKd5q
eUSKyuuWlqx5DYgwDxttJPtik8+MpJyS8199IGvM96TsSKpHh9jQd5lUbnErRUV7uvVzIAuxa84B
aVzdAAdPLv0iIlpBtkIjHw1/FYkDF8kzzy6n/6E4rt+n+Xd0+AtAN2QJ175vrOZ/6taCY8wKWI51
3hCkUem8Xa0CUPhBXwGn0lKZX1nhJXY631SUzLDBD7z8jMyQVViarZRZfFVSM0W8fFboKVNOYP9y
syZisKnFIhVVuUEVuoSQzVM9PE2ZfAs2adrCi58VewF1CHVs/gfDUuUMiHfAGD7BpsOBYiJD7X7D
Uxctxgez2xnuIu9NYyLcMaP7tvnUy988TYaMRRkGdEHIq3I1idUsG9gYM5Z7AHcHZ0RJgrY+3U/0
2CfgiER2bKnvd9fbG92dU89qYXAWIEBce8cuEub7K2HPBVEcRXmhaFjXL5qtfDw8pF8i6ObRBDdd
2o5r182JxXpcjQRKLbkQvcx+bbFzdGjMt882SEjPBymhz1mr2qZ/sM3yymI+/t5Lqs8+PFpKDyJW
oT5kVpHhjss4nAhet9Cn/MY6XK+oiEdpCSm1cZgue93oFpSHiroK6jDPJyjLWqy2/2lOkuofGyZk
NlzYYU4B9pXkct9N3k+3Xsonz3ca3AH2r645oj+RrvyKZl6EZM3fzl+plA+bppHtqgScLZpWALKZ
sWkydGlkLfl/m76id9LlOk+ne2lPtmxY1w0uqL3PYxih1k82arAqy9aUSFd74VHnUMNePzzZy8XO
27lDJ21SuaT5pyKxsADlvk7OMQkTYQHlumT2Q7N5OQfymYvIc4qrAtEw6dPp7Sr6Psel7oYxeFzV
Mwnko6Vc7sFDW6C5PSDyzlHbadhUxdL22TfxxSekJKEA1V7J6ii9ziG68+2Wihvkkdgaxzzu8mKl
DvT8Bc27XiY7t56gYEPDIfcK1XMi1tySi/8u7XQ/7Q0r8qIKVSGE+XDrnaAgs196GnDDq+1/oH11
57pqYMNQLpG/od6OW78Tu0BzOXCnVL4RHhcvftJA5KTbsV+Pso15UEUdU4O4KiwCTaXE9hlEec4K
RJnSS0id+eSMzL2oYQFNyehds3t4KceCDto4PrF8u7nhvCiBGBBMsD2koM2QgnqeANR4Z5Npk1Ld
KXMD4zLOVslqJAonjqgg9VEg0d4KtryF/92Bc0HYB+S57SafqtoS2NK5U0ze/P5OcAg3OwWTiahx
VSOiLzF1t+WZGDKifBTijoMu2GXvkRhSQtBKgJ3Wz79XxeYebpy2E1iSCGLOipk+0+1oc+6AuVyc
RSvAA9PefIpp6mYKl5pZ6fkWaLinLt0o0YB7XHOqQQbUyJLC3OmYpSDlmsnZiJFgIW7M5MxP60ia
9Q4E2FH2pFGovXDCC9t/Z423zlrr8GO/A8N3MyGAfs1BzwmA6ca7Vydm1flX6a4NzTpEgMec1BN9
gfRMWMn13wv30uSydk7EZ2/NxdWJ958jAsPoPRTgvNaATwWO3brRQCuyqA9FM1vbNQDkvMMUpL7j
tM2F8cFkUY23w6FMTte7IQztS4gYG3xJT3yRmK6vmhnyTUngMwuMd61nqvM8VBugAt/xQLnWkBcM
7Qli1XiH3tbRzBewlutcuw6bqQCwNNjj6Qp8JLlm27dOISWcsJyQqM6a31USljVGIeP09rK5lXId
2G6mgPTb4oNIrckhknfesEoo5+WVlBhgGD+3FPUHizq48S0lVdyq3lUOxdNGQzXdSXOhM8SqdNvX
tSQcN5fedDVSpHNDtYvR4Od6NvsNN/NMugA1WOCTnSs3O/CvkvOXg0E8Qs9IqH9CPKwFgCP1fGHD
I3uxkiLWjRiWFneN0hWZE7B3hAKehZU5lFwfjfnsyJ+dPk0q62thFGJSUQDUnLb7wNk/EIGwI/tv
TnjWdjXkGJ1CxDzllcKTag7CA6Gklv3nRPzhtSX5DhUiiFklWFfvkGvYf8YFmJ5/qR4DsfXei9Fz
wM1oe4H14xpv3DiwHAgb9qBhhEOwObwVTjXSB4sAt+1qaTLmEdwNrtaryuarp8mQ+Roc+LBjQjcu
e1EZQji3E+6L9EDJf/aPr95J9EM+F7hlT6YVRoa7i+QhxEkov8gGhF/GBTkqizU5CJ18kWGh1DNd
JGlJOpXsCBWLVF3I6fVP/4Vg5O25+7trKL1kUGUg1d/84N7xRgorxlHeRbDt7upaHwi4RoTwDuO/
n/0p7I0ptngi8qPnfp1u5Gi3iLpzEplhsYY7exgz+/a0RXQUHr0dl9PpEXtuwiKank9haaADRGMc
EZtL4YKhWWcwgFxwnDjFu1lIAXVJi2MMGliFsq9TmXx9Oy8QT7QwvKaN50Gy4P6M/Bo2Fy0Z5rus
jP/iptWbnzU3b3volcbIqCh7RC4xmZAmEBD+ZUf/DHlXhwWrfagU2qiGgd85FPYlJR+hk8IlIyjE
LvRxIryU5Pyukdytw2i+SqwBlzRyoHwTovf3qQOc0ghstFEZL5YKI9dZMsLorVb5VFtnLpbMPsYy
n9beoCkbPD8pp0gPDf7KuGouK/o00tX2nhFlCXt8IO2zCKP/+JGwdCsiOPvQcCF0qH0C4SvPEYLA
blNyssP1fAYfRkEa7jWDXXg8r7U3vKCX5lBwkbk6bJyFXxqPnoVuZ4CSqWau4BYcKc9mJCV9K2mh
zy/xgMF6bU3Hd5k1kHknO3ifMkTZ4eQ5lPcvOGS7AL+jlV2sVJadIv0OxSd+MV+DLd1NYlamam+H
wEE/9QjI6m7tqoHWfAvXUizPUOI9LyZXEMo8eox6cHUi0yyrnk12r8EQdJsFvP1D0swDb11bQecn
RR+oU0zWCW+3XWjbvgmOWZxeIK7ryWYqxJUN1YUO8AE8PAMjnOEEE6mFv7hHwLPmIiqNFmnBDfuU
ZEnBSJN/pVEwVdGFKT+OcWSXatKPVb0chUVmSJ3PzqcTQcoucVAooh4F4J7vGdZCMmWGxw0apYJy
EyriVtSJJUZR+IJ8eGjLJZD/sffJ9IjPJpkZGxk1ZgIwrftIgFZH0DOCcdCERz5luUXEy4co2A3g
2bjXyoPhW1HrvtQyNEdpKR4Kd9UK5/5rxKNqw3rKtihoh/rukF2yRVZNpGt6WOPnek7q82vzSHcL
Vb3oLsfh45sct46i+umAV4nifict1PR2G+ZixGvLCAuV3eCL4BgrnlblpsshQ+HXeMcRGR0Uc8Fy
eO0/XCmkRolH5Y7ATDSrr3ot1k2C5HXdRe+58Bbgo/RZUS9oC2kHfW9v9uh+/Ig0EYcCJ/+z8NGN
BJoPOfPj0XEObDWtHCaZk6e9jEDpgGQ7V5cMCLP2qu2kK46y6kbdJZ/xZZPd9TD/1wdV1Bysm5ik
vrumEsjjHMI16K4q/pY4oZDEQvAgLcovtEfrPPal3QYF1B7CxuNLT9AgpeZAxdxiVYNGC8R8U6DS
+Ih+lr3PPuuyjzWmyjzgZUz4FgmEOcWo9xZ093rABNwKD5hvF/fQrG0quyFZRUv2hITXrIfwt/k/
mSzv9BlWNqW3bCTGMwJ8875HfI5YC8ExDRiya15+uIt/eSJesFX94prxDKtesi959taNlyiPTdGL
UTYwh8/IJ+9J/XvGgwO9ST7MuXOgLWwBzSyKr0w9o41LrLaaWFsBb6ZnVfPhAbuiNRDH9cYBP/tr
t4vC+E9PnnJB9McVWBVTquxs442R9pmUkpctdrXp1tRag59zwZEo3vLInjYnlQM5i+djQuZxNO8D
oUS3cTWFNMNC8zAlljUzqFx7EtS2gCG3QI6H3W8sf6LtG7hTWemzxhdx1z2IQ2pXmy/vGvXvGvtU
L381FIDlHyNgaUmrJNqP2B3vr86mpttfw7hf72mHGprSBj8w4p3oFisz1Kd/HEbh91tWjG6Dz/KL
NHWYhY7DXBT4/9LGIKLbffj0CvG09MjgE4ph8JBDNKJCEArVzaQr+cqPAzyphg3ApfP2wt2HEpK6
IBh/jmP4ygmrIyrwESrLwtiTFdka1OPnMbm2/Pk/aYXqbsgB9yC7RNjk1bguIPmBIsOsJfGyVwxr
p9gYewsq/FVOKswJPCN97gUn3W2NmKYewzCrxIvszD59QQAR0RKokJ0SeR8WNE0gip8vg0pjpwau
GgfFnvpUxDq1UtybLzzyEPAYOS/7HAGf6n+XXCMU5oC7v6hv6a6p2miRhZkbNZHprVTKhW8yanY5
0375A3UwTSvNMPG0r5sUIm3r4AtNU8+WJaLvfl/eSi2G/4fYHMLqZo5LZtU71gmRt2h77ylNqoqj
BaDaHYyrpoz6OvtpqgdCDptTTOa8VlES5pFvO4NpWKK7wrpZkeh+MMEsqcSb6ZCanZJBatxXTLAK
k4X9MJocFqCUdFhn1zsUWiAVisa4Gc94YabdlNhpDZgR32gnCVOmNEC3aqUgW9Uch9zCYxVaWZF3
ZAMxWz4j4pEc2h9/g0e6FFODGRmcBr8mUJuWllXnXvWDrNZJHd9y5FXKreD7Zn4uhI5JFSQ908HD
bs8+K0UTOFfVz3dCmFGieHCnEsSx8Kupy0WSjRfKdBPAwpz0w28Y/6Eos2X9HK3OS+ucXEmWPveI
vVB068xvKOX3Q3zVBUchmEnbiKDrYsJ35gk9omJ2SX3j5G70qtaljGBam6aMTREy3+uB7qNGv7fu
Y7yqhw6eMPVMrQiej0tretqeme/m4NCkroVdYWqzpC/+Myd/hESNfmExWgQiBFYCmXCHMK+ulRwA
NYZShMA8zQAtoQMa1ezpQ/JX/kVaQgKHW27uScX1CVPszyasRvqawkysB/v5yvG72CaZ4C1wWFuV
3TdL2vaR3TP8PPGnsMi7XJr4+v9Hf9v+mM3QXk/HGU0Tu2wbjgGMzXYBc8jzjdvHoMegs95zCeAd
Wx8+JsgdJ7CEnkz755OGYY7kTkEDu71ut3qRSt8g6xYOZuVKhwdNCFjX6D3b/Z12Ok0uTEiZQinL
ROhG0ca66qKDOQ1SsS9S9ptqw/JxFJkRYyhMUpm12E2/cGyf1hoiY5SWUYl8XTXhmEc0+fAoU6zh
3FBl5AT3nWUUyDr2bKcyOC1Pvl/8yAKyI459DoYh9NjYMkZnLxJ1itLeIZuX2c50GXtUl73ibclo
tsE40HPSJg01I9wZbDoQ4C2S0rc7No17K5ugjaCzVKczO1w9RKT50dE/DXjGjfRN6oN/B5XLz8yT
UsO2QeLMBV1AOg3+3wnEmrwecGpMrz7OSM26tFdYfBstTOW/xK0c4LYuHOC76r/d8LVr5e6Nw2d0
MFq03vvM09KV4yjO8/rj0/TV0Xvr92zVKq4lIE2BKx29GdDDLdrWrboQ5gl9ouiZwlMnHfDQqouj
8U8+XTfY+HGENKVIVk3YeV/SxA1Tg4/MwXOfpSjyzpHPeNG/jMyZ2dbKQhMGPDsy4i9jrxVWP7j6
oFdZNNxYKdRFJfgVuCF+UPTiuTYyKbmAhmxeTRm0CJUdLE4QKDsR3zvPzr3v6AYF0Yw+i8pWFvow
BX/VQ/f0kRAZ2OItJh5b6tfJoKRowNoKmz3ZJ6O8VGYFdb9Gi3Wptb58t8dRUuT8rApp0sTXdrq6
uT8SWg2rKZTWwjEpMsfH1UBL7HJOIDrV6/biQXpo4PNfR18g6QqymlyGnpoXh4qWYytXblSx4Jes
vmAuT4m1TUfwuTF9pfMgUK1nob4wZKtNvUjy6J1pQJpiAFyA39ynH+yROfo9kasGTJKH5hRAWD3d
b8ILWry4W+no+H6qp606fTigB2apZt6Rf6X20+b40sx+oWXJrN+vWaIPm/s23bUGtvEvPQavi7pD
ybajRsmvjsPpnUAyaWTb0QdjX1WcJT9iMUp67bUkNuFv+99wKha/nhG4v1RrJ5/j+6zAYZ4hZiZn
2PytSuey4L8wdtcruv3pvXaaUWuWFuk3/wmEhggfkEvdhWvaTiDSnPZzWUyr4q68RbYFSbGU5fq+
D1Bne7JCFPUoZipjvYVCBH+k5230BurRd/VYnq6xvDPD3d4N5h35a5PUdlMeC7q5ljXfe3dXbmXt
Z7QOILjEzb4V2+Pk88HYXqfgKcZSrrv60WytSHwjRvY3MkCh+EmJqh03tFkj52hrUD3E+KGmIFdM
Jjy+uLvkzR2zokiPs3BfrFFGWtS/pFf7IRDjaSgBsSUzOxCFcdPUl98pKzTAlODkIPy5AFEZtNvL
wMyCW4MKbBFoNHVFzv/mm0wt7iL4wUV9j4TVGJ4E31SBAuqZcOQdAiHI+7GbhSK4tN30if28UiA/
icBA8pVCDkKmvoHt80DBy7tlQ449mwcEwrgvg9Filmg7zxnrG7TDAG5SE+emiidUZ1tV42qofuCG
WW4xChgdvQ8CTMjAq1IZi2cTSrTrUXAUgxz/zr+QiPdf+fhReQLTGHokbryCnFG3zTzN/yDMmWkx
H3b4t+oiAG3ltExIMFOgzjkozvwCUG19AG8ahgU3iEedOB1S3jkjszxvmJXwsPWGRZ9noB3IhEJ1
heZHm4nEKU29l0tXmBCNlMXfepLFr7QNKWmPIXKy/aO+8Q+2BaknKPwRvkUJta1piK8nzELRyhKE
sc20VH/89uId4ycz/oOUFuw7MZp+0uErW22Bpi6yuBJ9QMCELmwDkJTdI8HgYkMUuoTx2cT9mWik
7hd8vMlaxvu1bEjYkOAlx/S5cuETTfdKymFlm6luPU6nDvfrq9+3AH8IZX+tI3udHB/pqM+3QIVB
G0/6SbAc0byXHlzQLFqiU9e0K21+HrXI+0mxVhF6KjxjlCuZLX/fBxaGBlParh+klQwoF7Qqtx9S
cVLDn8kKOBqrEojrZnZIaST2Yc3w7SOl1+MnYM4Dw/D+qxRV3i6B1D4VpVMDEgjm1vsMHcb+SFQ2
g1oELET2Id/fta6KmCYDqJ32Vw+OXTkvqt2AnCXkYqnOyCA0M5GEEmglN4sPRzwXO6QPjxGNuZKg
XUUlj3zv/1Ar5mQ4RZgjloks8lm/LngIWOA1rHI79+PRUSmhnk5NK0NisQF+fGyBxcuLvJPX0s01
WQYLYBaVEscf0UuPl4xnliyFVVOZWya64HSuEm2v6qbk69BsYCgmevunOC3RhyZzaBd+1bdp7P5c
/5zu3whl/msQCEmyDfYhMiat9WI+LU44FJHCQxSNU45Szgf2Jv1adDZdgGRuceaFa1N6lbtjOwss
D8d4FNfeLHPZlbg2Q6IzjHDDZ+3BQWTM76bf3S9Z/AJKZblbdN7UwuThWf4J5wORnc1xCZVKowB4
9V84m3GS6XV9hSiOap2JHR5ahd00dNociw/3feL2XpEwWBQ+AVM98xsmcZ/QSdfGd2kneLGEXuu9
8/6JVxGy0u5MKxFMzaQv7EExeapyqWefIpUtNI0EnxM+6rkKuw+cr8TccUb2FSpvu1WgcXHkINS4
/fe5iDTEP7XQ1ND9pbTlFsd+bM6kN9qGFFNwEcxgjw2N2iy+3UpzMjSSa3eaPB9slj5bVu/LuKaa
0YkjWP72zqyszzbea9hcYuDZvT4oqNYIPz30sOWvQWMLU/MB+1eswZZEfa3PZF4N3yi4SGH3g8bP
PPjMoW7lNhD8AN3ly70cIwZGNQFIdKqzCwgOt+YtqIX4QhMMLVH8cZbaqeF39OdM+OSHNzqKfftj
7m6pZjsJboHI3q2uniXkEbUhCOtlghEF/lASG57DOHQinuLPL4cJ89FMGQtw5ganIE94kN5KP6kK
JG4R/GOVSJQ7WhB3AGQdEnj1MwyHWvm7uNPYN2MLgRzGMVRnxDr6zdnuD6wV++EUUwZYCeFZye3K
SVw4Dm2XQ75JGQGWL5vEoZ7yAFigYWQDpcCzFQTXb+scQY1i33aJ1R3edH6NQfHN4zynDzq6+14x
UKykHfYCx7/AjBic+Mb2qKhKhPldQ9T26cJfCoPWzp1mRHmlzVLoISZRYmyZJd8VCuWJCG80W+Ec
ZKJ+quaxi9JsnGIJoXO7zhV7TXd2rbEH58MtW0D33SG1w7H4Iv4whTNqcsN+UzxgDoABgPAvv8um
oEzfG4BjQMiRECaKrc7HSGauOrM1lkkmigIGFelgHcl7BadwlBo/CWR5Ku3Dv0ozRlwogZwzEeZY
Eoen0Ctl2z/tIi2DDm21f4i3YxzIZoXOdoC1HzCNE84F2mxULRgiu0bx04vNmNja7EglWgjw0fnw
yGTAA3d+BN7D1n11rtWxOFQHP6VPbwq17J6Z4/BY7+4WrFZP+epc2EFkLVc6V/fjpSO4Hu87qzuo
66qZA/o13d8qaVAxc5dHwSGkYB7NkvSiEOdVE2tsRz9T3mEyBX20YpEfbsMC/x94Nbmz2tzLVZkq
w1lLoX/OTjUAuI/d8VVeurqRApvo7ayy3+DMjsxYwXzEtCqqCUaqxQJ2Ck8fGzapiqDYBFlkav1F
EJuJmfQMUUM/Yvc2oFeO/D21wKpQfmi7RdadvjSAW6pvguvUDUHdR2FtVdXUs/ckFYCDqXsoicUo
UA4fv5u1W2YMERcFhuX9RebR6CdJkeApWoXGCuA5iGcxphpBSxtJU9ZjZLDXRae+kSS90WRYI2BT
vMFbt73RIwN/EDemFQKEEJAiFZTxgUza+1X+N+cWvjKWGz1QsLMTTUsWAckIN6YXGHcddK50pPsp
D89j8s+PirR4U5tSSCJZ0mPuoAEp1d3o7oi5V3QMySpWXs2ii+rPHbYVhEovRZn9bMijQwqKMGJa
9nn30q73Thm0GDRasEQMZhqMxJnG6Cw7TXKCd9RjO2THCu3a/XBNw3WgU6ITKqmTCOBDx1gTslCq
bp55p/O37G8DhaHC+Qyqj43cHAULcqsoRSqKSp0kySIqBbVg2a4+prSTFWUDSU4qoQwlc7VqjE39
0m9+X1zdwn4q7EqcP1R/OMZV8wgAQkiQgpACPTvERsQN/y7kE/Maw26S+KCt6lDT7SjQ5vwYHVfW
AWBqDm83iiSRM3HAGeSqo73inUYc0OQDH8Ds2zhi8SpgVNHfajLU7nyI+DwZbRsThp0WxORGwFtG
3udOk6NWox0xxsTZuvZbnmgtSYNN3Ls1OKSb8zu2MXOdJZAxXzjtQ+JhN2OTpF5D8rqI8Lu7mb53
aUQvSqSmhhhj41WZpRv6fyAffhvRKzL7IJJtJTFONOCJqpXbKtANtSP8Uur/HI2c8/YgRHyUlVtn
ISPlHt2AoiE8V5h0keiYYRanoB3BVv+bn5N9Jt4/TJlDUt/o2BoitFrYdRM7myg0ZVu2iQdmsxtf
xMmK3RgjvwAoROi0lt4+8J/nUGMVcYbiUvXPfCBily8ta04nVpp5wd8/+U9kjbA9/GAmC4ezmyg8
8k84NlsYKV3rBefYvQI8c6pI/jk7DSNmYQ64QiSg01GJmk3oayfsIcHrWz0ybJbk8tiPBiQ/SHT1
4G0Dc8XVt8MD2IgzNpcvOSO2b6Siq32dyCy4s8bxXvG61tQyXS8+leEVrJJSX16vxy3uvFarn6fg
YjyKey/eT0y8Ln3ugayNaDVVGliKuYkU1IpThaXpTLHYIaZhv2HiSWX9IevviJYudFwjn3+JIzaE
Vu/utvwfpdE7NiaU2PnCXPFGz5QiovB7bhK2hzpKMRuC9+VzlLgseZ1wnO/mN+FNZDR4V41g0Ggs
SVaWowmKPZeWFahrz0+Ksw8WAy8tcAiZATGXwkiLCFcOJ2lA5tHwZZIOw3Txw4rtv61jwfWL/eAC
7JwLzl6kXrWJl7ThuCEkK6UtIfM9HzcD+o6EX+l6RjrOe6w73ltcCEL670PyFKdkkp5d/87WeyZ/
77FTv7lhRXRZRd0FxPTqHvz7av/vw9BVOkWki/5vlTf+4wURe6/1M3baJghrw1697ikdijG18xN8
YqlemLrdVRc6XG+zXXwJwhqW90hNfPACULKP33ZZQj1mMULA5qpJiGB4NSYNEJDY9w+gDAg2VNCz
dqYNeRXgKByh6ORgsvcpaoo6xWi/b//2PvdBBC1gwgCkWSJ8WZLnejFlBrDrfIBefQzZW/NaEiFw
UlGx95eBuBW4hAVQxxfZJ5Tc0An9YUTGHfJsGevFFD+mLmig1snp/BiyagMYXT/3oC/UHTGPbWkT
pzV08i49I9QNzosLRSMlFmXhKxraGvpmWJplufz+j4I9XGcKW7DzfXbaEAdE3o80/ncFSNjmV9Ok
l4G9ot0pv7nPtZJqIDwc/m2JcY9iAdBXC5o2QdKl072yZrwIQkUmKpdRFKLuAoAUlsNvsp6dXqPN
kQNad0X6z/JYfZLPzjt/HbFXGAVeaPKZo8SLUctQlMsWzTDP1Wj+DzALaX3gYcJ85ZobGxvFBdaE
ajYZCqAnO6bWm3cbTF2rS0wad5TYZnyDR8GFp6mwTDUi6flz5/z8fKVxsrklnugxlV8WCg+/IRVI
PHtTLvZ8gPwvTcfImEzMkxKxbMnbd0aXhxRPLccIUFQStD7ZVejKUxpQXYp3YswGxzsG46iY0npJ
xr3vmwK6OImncNxXyNtGcpn02MGgzZTwby6BneyI4oUpgXc8zbyvyx3UejQi2LCIMv1dkSIPAsOJ
e37BldkYUjLM4mWnWwMrstvm5dfluNFXgIQRyIoNC8ITyeKNLOp+vr9kfGJS8B3K4rm6s56ipjkJ
0G+IcqO5pDFmKM5DGwtjimPd3stj9cl8uoapG7j5v3jW+LDGh5ZwkjVmb/MtNUg5kBKlH1aKdT3c
HU6o/jFmU/reP279Yqu+d8K0vDbsI09TR0EqUQhXSrfD2dyqHbpKdEOljbSszLXulsygsFBV5rzI
TB9gzKLXkZp4zsNkCLT46zg0RqXSC1oKlud49kwuw2Dr7dWNlJ4f/Z9NnasykA275wtOaOumYgDX
LQnFF/0oNNNFn7TIbOev62Ohy7QR+qe0KbzcsS+qdF8FRvSUcm2oiWNoyydxzr3W2wc/O2desF4S
GZ+ESr2k+LKzoYSGHa6qvXAAkh0zAj62mkLajX7Xv8gGCGgitEIT1lkHQtZ86tQGCDCTnRUN5EjP
UWjnledJv8yQuanBJLTn+iwnqZ77w7QC0wPDmmIQOaKUzGn8jjaTVPdDLgXVUkUwQhVczTIZj7BO
D4hmn7YAbZQofeoAn3w9YKude89yfV8VssHQ8CD5aKsX4JDocvgvuzbnyY6YmlvbYtNYcm37wpjf
9fDziYptsdmxYkaoZxeExvfU64XY2zP8ZVr/qb6mBZWEsmwBY/ulUtQjUxJv/exWtDFbtNEWgRQc
YorjHaZCwPErKrPA3zHeOdjU7T8UdVZ7R+9fGysRh5AhRWtNCvKFytr46gvCN2QHTdqfI3IsO9sB
XdAhaHPh/rzwKaKKGV/jDZMwPmXQCso6jAUros3Zeb+DEG16lc6qVNmCmQhGqanCn+Aq6qnnbZHQ
Tjmc4UgxUPUcF0vOwjYWIZiL5fr3wBG0ZQGQ6zRa6aNRoo7jd7LJytxFOBsjfE5zo3OCLO6NL7F4
I31Ho9tmFRikC4xgS1HnTA85RxaOhxAInhDwcjxOBRAeonvWKhuqdmVmtInYQXmxaUJ3l5iuLmRE
ssfQzhTZMK9qWPABomzWyzdFWa9ftubt6V79IyuUWQWedSridEqSgkgvHxzdUJ5HfiTitEUBnKq3
5sYTDD1CmgKD57UShVDLMYI/Rkvp5gZbpSknUeTnPIei2sIvLlqpyREeJdmwDlqiru4mpvj+XfbE
gdOW+h/ZoBnwA1JDVSPPrGTaeSfnUDa4eQ2Do2hGpI/x3Q2bZ7ZPcXblhQmSwtLZ1KsRdSoN7HPs
jK1Iwn+JUfVbT7sO7mJPYKpU2SfeWC5EoIL/Uk9aDXjYi96UFx+kmBawGHqzv8vgHVrk8IBY2E2/
1F3gwsieRagJegEen8vfmNgnHH4bnGFexO3E99WxhbX0+g4GKJg1TkZSEf/iRPXwTrrelWIZvKzR
rvreWCqHv/a7266yl2oVNygufzfCHhi23/X+e8P0GaTtslF6LTkBgivqh36eu+vdie3J9VnI0VUU
+gFMSbYi2hR64+jdBEs850+QHpbJ/tXvF9g9uK+IyAjRNuWp7pcfE8JjYi6fXg65V9JDlApApWe1
cLc5aCcbO9hehpCLYbStpvi9Leb3ErlVFL7Jrn+dZBGE20mFoMi5JmthC+I/dYsTn/+Jduf33NAp
9+zRtsX8dabpumOPwvlVzFcTN6RQlY+WzAhVa8IhOkNKpneutD6cQ7F9IeXXTJmBRQ3gDtMWH1FN
EEQ6tUx9r1JtgTREiQJlPKfMkDwAz9LP/fvMSx1hOOh1QHy6iaQs2DbV49pK1MpS6tU7DKr8/Wvd
PH+EMraUr10SeOuXNeYxBr5MSTwIGEZEcihVi38zgjQCh5zNPuNbEEHT0ep1LUwCv5/QNN+hdKnz
5iSmEbMY4v/g1AvyeoYIQGvu4b2A8yU6J14YcPokrL7gpm7LMmUjSbEveS0qrhYF4qvqK38vbTk2
DAs+EUjt5kTjFNGJzJYwubFGO8JHGzXfNQN99DhEMWsHG/8QgzuSoHuo/RDPozt5DM4/pdSoMGvU
AF1ZvHcWsScJasGuucVKEIasaH7flidJCW+DADgAH9UWcaU79krp4dXvdw5HpjYyi6IubvNzv4yK
8txSB7lCKLx4FvbS3GU4LNCSz/KgBSKkucU+eHod+aIWrt2zxn6Q+e1RDADyI32Gn6UwY+Ts5ZXF
H91dK/X74KnXc8LRzLffjlvYz7azC5qZ/Wk2SxdcaKJ+gJXWrrLxkb3xXmOvIFFcnFEMGcbsrVOQ
rMmAVUb+44kh41gpfBBsCmjTgF3CpMo0pDLIlBQlPBIWcDzPSpkS45Xk/riOzzp9CwgDdd1UvY3/
9/RTbLC+UrheW15nqM+ggh7lGGSnQ9Mctez7F1mzy2RW3Kwe02uYM+64JmhtPutrIy6qYHghNre5
u2jUabd971XduHG/WYIfAQ9GefjcFhkvMrdsld5ITazkplvPtNPIe/f+5GtivAFvjYFnHytkT7VH
ztXD/oCcHbpltpYg+qpDGTPFXrvU9Cyd43WgDAw/ORCTorcZCorkky2m6i6CAqX1pWOgrqseR13s
A7moEbG3GdpJDjXba1pLL8y7AkbwPMFdXQRAQVwzDOLWX4t2ZYAcljKbiREKy3PucjMQSnRKBxrU
XRZFiQk2Rwg64qyziFjOUflLoCNq2sPL5pf30OyS4MZCwi1IiUKqsMCJ3E1sMnDj5c9FlZrYV6Yl
IWRrjfG1RVNNs2UoCOjIZGWbpzRnyEyn7/XdsmpQKcs2sI+fAFM3ao4A/RHyKMEAEQ/K4GUp5+OF
8k2Ss6vom3CHPIGfmVYDOlu6RbcL3LwEa/5ZahU+1qCjudSVxK52TGF7Rp3FaM9FXMuWoz3u0rrS
WJOaet6HjYNcegt7vxFpC1qzwGoDN6sUZ4h3XBPhsGsfMVSvhoNoBgDzDlPku4685H8xJrYL0yyp
+drdJJK8w5mlnLUo0EcAuh+RrZB8G8W6JOrmD6ySSoJt5zvt68ky2sRGwsMx3BKOKVOciKTNefS0
q6gTn9t4OIF5BviO5oY5aQCA5konHW3HiJNHytkDpVGhzk9pIn5t5bs5+oXF5VFMWmG499uJCYd7
hG6ZpiNiI+5zIFJcasjkkZM7KcobjCwQOIHRGVBxCBZd1r4gYpsxhL9BxYVqT3NinZjhMBGO4Vhc
1ojhTrLZKt6bOPziYmQJx+pFGPVganCM5JARva7+Z6005Nn3qQXan9KqHJSc5qNXDd3a2j/PQcdO
ovdqpyYpAQc7ZMzfgWib7d6VoNqhHSHM+PPTrWh5P0oltmGxC679y7/1U6v131N6Pz4/AhghiN5h
HXve51ERBaejSJTnR4SIDtb91DcfGYQEJ9t2trNwiwpD9vxY30/l4AqCMg8xXfHBqr6Dt9Zv4evZ
uH7zajHFThJmzbCMx6EcMiqyTimAh8aVE/IERK79Gi7HQElzcDNEE8xUN/HRq/1a4kxCH9H18tf1
whT7j9W6cLqv4vHQVYiEtcmsONsq0+6reUZdMnB8yL0lnphJxNfZdDdxaNDXe8FNIcIkqjk+c1wv
MYRxiO3Lo0n8kE4f2F2/swrAxbzvYJMLK26C7QXMPM1+Isq1koT4DSq16BSz/1x+filGB92Yiuvi
Mm5JEGERkEd/HbUNjW2gTNzNXriAAdFFPxmAIjRjtSig6YkGOUJsgB9KAj3XIE2ombiEIsIw1e1x
VP9L8rMgH3N6hooj6nkG2aF0LCN2PI6Dhdva24gYUHp24CgW4Vf+a7YM+DeVaEVpmOAi2gjUYdBU
N+49Gmjwsey8LaG+ofGYbiqpE+2LwvJyUqXg+iO74NNxyKewAv5U5v7rgmQI9GGTdvd98YP4foH0
T7ovYQbitL75DRjypkmPw9Ltlf0SG03mbt3FCS5vGIXsnXAGoZUqjKQfIFNaFtP4YOMrzwYokEiB
qyfB96c2wrkkD8E76SUto0ASGx7ahdsiNTNqSeESQflmYainOKN4Tfeb/thkQkfRa1/2CNX2Sd1W
wGwI5D1A53Ure1v8k47ZY6idUouHfiaecNbBmihhjIK0ixwj/wJVI6yJ0lfkNzA+vfGWFFiGwaNr
NS4WTu4+19iRx4woIVnHooW80MeuUgF4xXVCKq5yJnEvSXudOhivhCFIZoRapvwx59CIN1N4fZsJ
41k/hteGYwiJBMahkadHN/ZYlhzy1uNIiqYDJ7tNalHzxd1AinM2kG5Rchhdkn73jVGPQHfYZyAm
Xp/+M3ZDdf+djhL7kv3brROeegRB4huzD7ZUALqpu8hT+aGz/ic+mCMiMccTeS8zTZ2pq+mhdtXr
DPIzuINezdmb6FE+t0+/PfOAY0cz87EsPqZsDCeqz0sw/rsoIVC2cpr7e30h/aRJbl9LUKeskIHt
tXNNVNs5u+Rkr9Wm3P/VzAjgyU/uJeP7OxBa48W7JQ5nx/vQ3XoswQtdowa+OQzRw+DKLp2Z6VWF
+9WZkptEUjZjlSPnfR7dT9Iu1HI9dpJ9c13ExJqSUqEiofomDCvU4y7fYpUxtJQKavpQAxxM1peJ
98iYAA5fbrTYVWTWGXM6H2YNbKwkipyijEI3zZaz6VbuZWSSDb99Bcgo8u1k7vTY17K1espNeLf6
aQHrkY0YrcRockJ3mtHEJBeY3N97epfx+NZLEjKxe3+gkwOVCeZoD+gYymLjpN61ay+BSW+TeAUx
TLyiRhmBxDiwRPnr77a07WUyl97kavPWoJ+c8xK8QyWfOUbyHymvCHQGypJZpixJQOdZQuHlULaC
l2lYj/cv5Lj+S/lCI+uOfgkPhEKpAGNRVM9MpmbSj9O+V1USTQ04J010DkyklK9THMEzPRROPnHq
1Y3caMqQ8W6LHm4PchJfXP062Adff/SJGAWGWjE075ZjEyM/cQ0BUOxxihzC2a0TmBWgbFIC1J4s
Hk/SnuHvnBRbJedmiJJMVpgpOXblkTpUMkvOpLtvC4VkxFGw3c4FeMWlIFqtUrs1u4PgQXrjAVfd
vDYGKogWUROSyT4oUeXE9BHLzL7e7X6vBfpBpfK3Upy16OASJQ9FqKUFtrpj8MNTEtgyKl0pIV58
x9SYNz6TxGVNW8jznSB9G4iPitEm4MemShJkM+vhw7BeQX3fdcztTQUuZQkEL3N03IHLGmLRcCcx
z1x0JsQIhmCbyLpZx2C/sA7P07Wulh7GaeXvIMHnJAWtpWhMQEcUozr0MkRORGUin9oFrbFNZA5G
6GkanKkNBy/cGaHqWj6NcLQK+icSJ76Q95RUNWHePsyuaIfbFIacwgbvqE7sAikeQNTEhzMa45D+
qMQ3jS0PVPm5rkD02Nd9NuUrwKKFg8QhXQsWFffl/cVmbW++K0a6MpWkw/40r2eoqxqREfTlXZy3
pTidWjHWi/8ZVcUnSocD0FQL1o+TpLItTpyDkRXtJ7RinZWcyjWSevZOZHGmNWfAAJbHsGu5qOI7
jZ1D4zOZ7IJl4myru+u4hJEXwHziWZWhprUUAu37rUCbUHGpGG9BRL6OxhgVirZfEBu/YTRR21aF
Gmo//kGRxj1AUJD0aVGHh4kM/YEVs9KYicAD3M1oCc3Q2ul2M4ALUGS4doFbBZnML+IbnsOtK9LQ
PFmLt5cNN22Pc2e//eKuLcag/6txvFz1T4lASkuVX0kj+4XpaWz6iS5UFuF4RGahEcTdJ1fy4hbo
4yKxojFUGa51pElCWgZNRFdUn0MQJ1PP8s1c/Epz9JI/br4UZQJOex1+yS0SXP1apsRBKOCLEllw
wKXfzhAYVhhu/4aOg5F9677c2CTBYrI5IjxzpUMpopNo7jJKGQ/MQG9VAnlXO7ssjJHPaP+tV7bI
nWTOJfXIYo61rm1UN9LfiEPausB1NwL3+9ULsINJydxVpRgCv8grwjwDdjdL0aoHSKqX5kiATJ/G
OPd9YTUblvLNcDJnGtKQFXaYdHUBznlXgDe+UJW4oFOXhVfN7Q0hJhqCsG4utiH1k9sRMF73B3DG
Aj0syP0z159o9QcqJa36N+t2mgszivtNl08wKCWlop4z8REO8N3lGyHctK84SEKUS20TDMry/DT2
/9lyBqCg6PnsquMJwLbJOewhGK/+5qzXhxPM/vaHRgd4zJBX6guKtotcmVSRuURZM2baHkDiv5BR
W0SkZ8GqpYuRdIFjNyxRDG/bOa7v5MwkuqYRqzBMvuVLw77Lu9/lLkh2ZhgjWXg8tsHLNoYDqi3q
afHnjpkI2MjdYUTRMMSN/au3ZtWfNaaO4wci7/0Y7wq843iPtehh2WgVo55kvNEAzGXe2iDnL+Fi
+dvB6Zy3Kz4qZFSSHpg50nCHUb5Mm5tl+dB0DJL2i5Pre1HhVnhMBer3OhJLwGpImC+FYPCoFHvW
9Oj1VXYHdo8X9cdBDQhpbpQDZz2r90xiN6/XauPFC3L+6AvR7Oorma0ZdmY/LNtG3leg7lLGnzdZ
urpuoc2PMQry+8Wyq2qZb35HD0ZWeiViBHL556Tvgx35zU84g/Shcd2onhn4YIpYp8+HOZQxJDS4
0rw7JGfwobpk0VTIJ6xWMe1J34lxOMbqVhuH31hPKea7BsOjRO+dbvUo3MC5cl0QyP4qfN71SA6f
krMAD3woHoH+gABPwoGO32KITQJwnEgmBOrAlDf68SLpVkLKgJZqYqrawFhXTdytHCihPa/yZx29
QuRbQb+Rax2/YLxc7HvGAcVuPVPprroejXIP6QQqjVUlQfKVtXF4b+Kw3Cx73TuhRh6WIZV7E/Pi
+OJ2Q9INgrFTzkUwB9lVJo8FoUQaPhqGacam1nFU2/EQNNlmih2nCpNguL2z9PyCX+qNPq9iKpj9
p0V9F4qcLX+QZDGnSsaSmGiC8nFsbEOyNB1RlKCyuWF1FPIyGszog+ufL3fzZObaX+TDjlyPUvYa
dBAUGHNjESyTZhI18dk1udv17qXFvqyMAcT3dtyDJR5J/ojtcveVHDwBBWnktBDID691mh/87X/J
N+K5+lGZV9AscGahVsXlAGxn3LJw9J/NBMGKWpsnZQmCC8hfy6eFSItsCtUXH//PknsTc38faHrl
WgstZLRpy/Z+Xar1XmRQwHd90EutBlFBRqR1kc6eX/1zmjMnRLS8TYDS0dciB53+KUokQ/TcP0yz
2F+mZ3KRfKuQhwPxHCSE8L6/3md+ggS84CW/whSerKoVwwXZUbWOEhVqUhlgCMbstKfCuYbI1UK/
uIrhH6tJ/eD1E5WblnkwX9TD2zB6x7mX53Rx4TFC2My9VUNtGaMSrIijFjHfuy9LIj3SjdT63gK7
bJyzKrhEJiTYERn3igzk6CudnToIdx2Mnu+hcmxC4PIb/FcUJ9UlflWT6bEzebC/VMYXsD5SZ2FJ
NWH8GIE0hd3uRRBpUWZiPcFY1nvv7JoDx0wssuI1c2WTAlxoUuqAT6hSlAyk29Q2FvRmsJDK70Sw
3niP0rCRfAv5OTJVWAT2lkFIFv7OCq78v+7ep8AjHRc76gZwQLhr/Vb/lWHFyZqWaRZxagDjOoFl
pMOJmKqfV06f06kF2tzrWDZgc2cdW/EzWTaM/74tGK225HJMgps//2yMpyozFbtRGS6/iPhjWCYc
dnFjWRxIgYmZ7ZO4Raa8yp4nwfLe0Ie6nGuaXXyyIihG8z+4PLLcm62mOKCcYi5J8ZVGIR6LcEBf
K2PWxT+1+5C3q4TXQQwG6JcKxuW1ep809DsS8HPX7xdq5GlgN59ZIvYAaIfocpHgK6u/I5laML8z
My4exJLVt5sHga6nZrnLMu4lVnQNoEc5fPJbXJRc82hPXRTP9YYMsNUBZxfjLxeHdsAcPSnn+j9U
8y3cZKSICxT2b+kIF8MHGPjUL+Khg0FEIY2RHXAsXSWJwmN/2s4EaxOL+wvqYsmb3wtiNYimP+k4
UH3+h61UUg+YJI9/Hg0D1sv4em4Aiyt1Gk2QLCKrqbT6DlaoTUZvBik495UHfQReOBVE7LMgXTP8
3IOzpSylHHXyqTRBhIDv+B/pH5rDU7n3WJGFecNG/yvQiXoK/StfZ3rOQDCNBTFmLSQ/n8mfApc+
Xou604phFRKj0Zv2VBURMXgsM2CuP3gMC74nyd66p1fBTx7IvxN2uag7EGGmbR7RPDlNObmzlyUc
qk9Kfdqe+x5089ULQeiUclYvtmPjrbD+e0kowqTOzWigThaonvrWrCsCkhaqw/lt0ULVS2IfiOKH
t26RJ8D2uhwFYT8gFKMEfx4GEnNM0o7x6i6rMDJD1xjhDEVrO9lpEmESxKpFPX5cGfVi9y8N3rtd
uefwdXl3l45lwd1Z7yT4BGRjNDiFyjejgbGhXq7qt40YNrkT7684n+ecoon2OPFLBWLu0Ao9Bgcv
22PZYsXhidZJQGcyXk9WyzfBzQTyXmC3mq0Dg5NZFsrCVChkE4w3xcffCt0BZ0QWK/bhkksgf9nX
/YL0ZXbCWdeQ2G9fSVkLNIhbYEtS+W+MmE0FwzwD7MWHonvKJaKdXqJAYKv32m7OwE+73ZoZl8PO
MlRYqWtIQ9KgRGA+MsKDOkaEo5GavHlp3O9tXQRB2pCq9+kSm6xYDtBIY7rVG1mJoaWt5r7coBlH
CDej9OtOt8bfuYQN36bhy7Jmy1/JbJWMGIpM1aASopfEAyGUO8a2n+oetS3FUg/gtDPIlor36AFC
gQT4eoxCB89gFaEFvAyoDTVUP2yDAsbEun4tZU5Up1OuYNBteMrF+rMYtylfEaC+lQdA1+vCiRNU
krzGwoo+EelEZA7w4Ri7M3OxJn/x4TmoSAaGqLfXj6pzON3eM4HlsaFMDMyNECnkjzFvAMwQurWv
iJH6TW2qNY2WWAWLbnwf6660FJ2ZXhlOPAoU18H/snfyGVFR2hmvmkrZryr3QCNUmaQqVdAmTZYV
U4Drr3nRaVgfjxOeIQW7dq/8vjS2pzxV8ICXuYSwiGgh/B17no3pLwFYLYcElCaeAMzJPp8SUbkW
P+GW9zwmyU0lAwrKLLzM3ji4PrnOcLWvZZkueD0EF6czOWKh72kPndnOF97l27V7Y9NR5JHzy0wk
D+/C6PoiYb7rDIc3t3V+eIUVa9PaPDyhg9wIxCnDcD9Tg7So3hRNkUxzzM2gNuNC2ftfyx+jhWGp
FERBDQ6YkkhdRhBk0+dzeN2iigni4764wGyVFaIDEsmpgIqL4kDzkdsGsyHxk1VA4M/ikYD9lOK5
qEtL/U9usu+qdXxFvaMq2LIxzV2I6dL1AlhMtBngUqP0hEoMhuJa2hiPEpq+jJlUJvJMT+5Cjv7k
QAn/L5AZ6sIjLdKeaYYPV7TVZKfBtIUOsoBjkJNZJ9hhKoO39KVhK1wuOxJMzAwGB7H1bMRF4qi2
9m61c7dkccC/99xeBnwnCpORrc6jr0HtNqv5EAP59lf8H29jQaS4aSN+B8fbacHIkxN2Mwhkne/M
zL5dNmTYWtgx9auym+VYdefF8vXttgCiInAkpgaXmfsiUNav1625sVqN0c9kF/JDzQ3idEG1tsuJ
DUPk1xnyF/ByX5Zz1zoQ2em8GbpWtWnOgQRBB8fuA8bKo5dwaZo9oiahxgdE6TTvrIDMUiqtUjDv
3Zdntgu/3v3quVgJDsWHMJ74w6Fag5bmwnI727zgdB7XrO818yPDC+gDxZA/UhZwkOEvnq9jPTAN
rn7/iAM0n3Z547sJ6cawg4kzT+mhuhfOjLqJ+13Y44Hxvd4oKhMqStVVmEP8P3a2Oj9mfSum6aiF
wvC5HRCxfJ7ETQNkWyy0lKK05bY885iWcWDVOGgWwhloQBSkxZpOGUozIp6MJpIkUtAVeN7iqi67
DPEgQPVe44nrg7cvT79eqs2qRKz0XhwXRh2euYoKM1JQ7/8I425618QbWgDPL3ixvsfvXPasvc6J
igOTbvbL45Ldpg/6jHW/pUkfhbkKMcnn3acYru6bzjhKfqZUzIUY3vDF6GEtCUtDAek2r5UKyC40
YMcGSE820uePaKvkJk2m9iYYSfScCmmt1pLShffyt2xAakFJRKjYN9HZKgmi6hGgPEvl+kJsIWaC
xjKxUFID0np89eq1i/UazSi7rG+BwIG8r/YM1J2sfmvOenefsSASuZl6O26bpLsNvFw7744KGSr5
3dxV5kkNTjG28WcFM0OiciIycPO9MjIa6LIF04ZI29SVdaqoGhUQLcmWzyt3VRHNWbLKJDRY7UOj
uYIheGfic4kIMsTPoZIN2lJAFFqEG5M7itZlvxyJ62k6RtNDzDCh8fsU56Iab6ueQgdRDsdPh8TT
db4V8ARIgKIbhD9xjNTMEL8yNZsWoYVndADmoT6Fzprcu3MWZ/0wbLt/iifGe1mhRQZ/URKBaZC3
tMr1Qe0LbJ7jO4w9NT8SOfAvR7fDXE5cEgyRSylkFwJ/en/TSpmf1AhAfAnlAPu2xFGRko6lPJ9K
mGT2FAUW6QHnq9omnhL6qbh/cA6twRECpAczg/QdQ0Z47uuo87ZCnnMvdTZ+Wkwd+sLanttvoHJ0
alMr9NBAmabRZbhLAoF0whOj4+DI0qOqvIhD97pA/MvwLwzFEw0Xr1pXLDjNmOE8O2s21Lsg2fDi
8kW/Qm1fZqVtWEgxQ6ZPKkBYZq1owLg8uj9xAUSlst9vFqPnD/yAXEgAdYmphjFcoLwe97lKRtBI
0KLEv07Irh+z7IBpJTDbH2Obp4j1QJ1qvKC8oidIH+TOQ3x4lqmelMpkC7g0LAayrmo1R1dt+VSS
IaPyCYsqYiOr+tOte7S+R66UpQaeP3A9yVWJ2uIHudVbydGVj+8JTSstPHD0g4IHjhJ2Ye25ZE9X
BpY5A8aV8lXU0oGqeDI6Q3k+K/LfU+1mv1kVTO4gZKDtBFds55AG/1P7CJmN3un58Hr/kb4QaNQo
AINk7VW1iRzQRd011LY50jPcl6L5muu7qHzoKBoaMGm6y7eyuGLEG1xYvoaeSpMX+qtEFphHwB4e
sH855j5AbXYNqQLE8HiqJPwkEI8RDnlY4UZRhiRRnka3cNLAJ3kPfeBkjgVeJheT6286dl8XdEf+
kmTb4EeXCriRbgOL+KDuUQqNx3eEJtRkgjLcX4RQrE2irKronaazaS1R0MvrpSfKKsNmAmTa1hbF
3CiyOPYBQpy16c09hMViXCBMSOMreixo3mu4Ox7dLRZaMq6/6P2v2blI8wyPGKcWuYj3nyGLJ/+x
ECm+xLYLxZw7BLIAebHGoxaoJgXEeCvqYsVJKy6FInb2lK0qW6XpjdgagwGX4TW/re9mEnU6rlCy
7jaxZA8WaRIWdld8B1FDjhdAj4V+z5kpeP0q1zUnr20T9dZFELjSd38ybKEeZ1hdkm2u5gk3hz/S
o/HL5FV6573YZ/6QYWsclz8ty9OOZ4O77Rh1+RNWocyDxZlltHrwWISWqBt4MCLDZRDYRfyoJKMs
0r2Pe6ppkg4nuGeClH8Yi7vNYxp69e/7Ww2WVZGl2m8pms7SAcGiqauTndvssIQ+xQT/RfejYxhS
Y1w531U6yYqZxjrri/nW5K8Yw4c9PbFStCZfCJ9Kv9H6uODq+x3bGkmuE7H0+FxyjahwK/ZIPyJv
120AvlYvWDEg4G0Awhd+haO9ep7b3zhnDUr/fDbEd3VNr7IoJZG6bqCWM3acAXtIfAwo/heFGmj1
Gc9FgwbJ98NujIzmUirF75g702fWv7sRAfwulMh+VnYtAn6y2mIfsBMrn1M/1zlGkJd+mjiE1dK6
o2E9rJbJQBh1w09kwGOn9MOgj08Sq5UDNugay0cD1Gzu4JH1QSt8lm3ngw6GWMFYltyc4Q+gnCEd
Q8Jv8MKScJ86kfRjAGgZFQtEZUWrzfwaFcul/q/8Y2PJIMPJpQ4OtI2W3N70gTukmB+J/QtmKxnX
wS7Ou9Qai38CeCHZlg1aWI8dkKtMai9ledQ+Wc0KfnPVb7Omya+kVHxocb3DvV08f/N9QBdxZsJW
euSIUu8MrV2EoAa0kIfYSvsy+aOOHtyUiu4EOdxScqAh4lE3LGokYA5flFrVyE8InIKl33LHaElW
Bx54hwLAAlzU5ejjF5fviX0R50XdUSrcAW1kt+09MrQ07Xad6LB5HNUb6GpfTlJZeyOg875bfKJP
2zZ6vk4sry/cyBPvB+L6FcXhD6X+MY0KdqVSznLXnY3Mm3gJwCju/1oGdZRPgDs5tZTj9IUNm+PW
gGInQLv2BBjUpansinq7egiwrOqRFPJVvthOyY5y3Y60ChPqk3cQigMnwKlooB5PN/+XOMBG9U60
K1IweDLvcWn8+toT3jq1OdqnI0g4Q5483sAvdWcIlIjOicrXaQF7Lt4C7GQbWoeZogexyS/FcJkf
kEpQa1bt/byOXbI6hQoXVderdumgnxDsa0i5foAlu3hZg526NLZMlVJQU5AYKnaffnP+NX0c5PU7
olA1/EjJlxEOHDZm6VAomWyz1hetbWohRFb12ywatXmrUUn2PRiycgXDMTOnM+xpuPoxFV+du9IF
mGT4zooPYRomTDYwlk64eA6NW9ZJnH5aFOb6WB429Q8PKC6Gm96K9YTOajLMvHD4GgI3ieHOigHe
qr/B4x3WatC5GqT/3ZbRjwe6imuc1s7leSOaswEX24Ipby9avo/sPJUeoe/URNlO3vxecVPW70p3
34hBKTORkl8rSgABXXsnB4LW+90w22a7l+CMTecQ1+LL4i94cPGL+tBZyog5baWlHqPXi9XUE5MC
5JUnNKnmyolBgoTFYEfGw7M0hcbqPbkw+w/2dx2ovBusDR9ePmChiwACuP/zA4D1Afv3HUv78vXw
atw60ZkBck6MO+Dkuc3tja2UtR/e2ZAQXi2SD2aiLkGZk0sr6L3/GZi+8AkuT5pjY071lgVtOJsZ
60Mf+Gl1FVN+1Qj84Uku0IPq49oFC75SKKMQQvwgPW3E7pWhmtxekVLJmiPqDwEzax902+Dctd9S
gc2oy9qz9ZP9et+alwo3D8vOLFODch6KNnuBWBvEZ2N71I9sQMICVHWyMq4yQ1HewaBkiz+6GwDa
5W7ykyN161yhwvYQfPevrmAhb27sJIClGBtqpVpMsX2eCfvkSUlX8UOsf3HdflNhSYjIeehUmn8Z
EBWhnGw6XY7HdgirVhEhk+uA1eVvZvJnaQeAYEBiVaviyCrVc75/NIZftrAsP6NF/5CsD6mhcSuJ
XofzcdHmhyU56EyX4Y3lEI4V8j8RV2IKdabOK2RBzqTwjwQ8llBXqaupyZEBbigE4Njlcc8QR3Lq
ps5IN22hW+Y0Em29QeNJh3oEYdoqomjLK+SN9W1YrUEgvPGLEs1SzDyUM4arAqXFurv19ikLUZz/
ENhoAXcnKyfJC1UYCznpgokKkII2S5y0pKNjEDDSGsBS5aQWMpYtPbJcKX/4vluIw9JiLkO6aX/P
qsYo4QQbagFmxRrJ6CssPauhF0t8Ue7Om3CsfjH2oNtc+Txa/e0F2cTtj2RII4kj39wvK2gKuI2Y
Ii165/D1VKWgUJ1+zslPmVRXD0wMNGm/ROD0odKiF4qSz9+X738HpzRFV+wXAmjhuS113r/XKPvg
zAjjBtc2bJSC9lsQkiVsbgU43r7YlClALfFrPBDduMSG+DWO50alVflT5cNkcnJUQ4AISl5jbedW
dcXruTZWjDqzuPnNZ7us89fZCPAzaddRovYWzyGkgdSwLEeiD2/Og8VEu7vxdQXkTTY2Uuf4on3y
1wY2N5TuIw/GHddw5dX1vZw9u9bUcU96TAZ9Bl5cQH40hj49nhGmtakByAAMuBXDdlJEISkR0rNq
x5pq1FHQ7ogorECxk3lppP5d/hlinw2GnerXHLldxMy7ExUvfnj8WHJpBHcqr9c7cB/aUiRKjeaO
sk4zldlzqnerfmcUpAAR9O5e1BD0LhMaFYiqsaOQlpW3FydL+66WJQzrfucXerWwsVExQJK6yZhR
4BfnwQ0yOqB+CkL96HBSPV/bA6FrI1nGUMZunjaK7xTzQUZblX6Zoy22QZH4JNErgyIsOzWsmbuL
bDJLSvB7OlB4eKktyZ5nLkVU7BQ3HRpV1MxcA52u2tE68DhvtYc8vPp9gCyg1tfxoz5PJgFFtaf9
7Kcn0RpZG9xH4HZp0Z9yK22dg+EWciSk070IzdljrS8+0LLMTHcbH6yY5lt8NhLG/wOy2JgWsaWS
Nn7FobtmoKISLaeENIZLmRjpAKqsncIErojcijg3aSVdvsGKy4I/6+XypGjko0ijTzfrf1pRIH3h
ofR+SZbGbon1ZFdFoTouFJPNXQ4P4DEmALuOVvem8C1h1lugTqziAp0u0mIW2wfXOOAz5dWCV5qn
eirJTLjDoiVZ5Ar1KB/+SYmJN0j/jtMcXbgb2pBWu3FbNgHXGKeUgEmsN66g8PsZOrEbwMT7Oxmn
Y/1FkmQ0aixCobbDAmhAlt9bBn8MaglvAnSXRXhZ71NTKtobMRO+y4WOIdVl//vTzd3zUwiOvHw0
1AZCvN6HwTT+ms12AMk2a/JRZT4wLCRYDMMBsLvoFkNP0KKEil95MUfO6sWDBhC+6282cVHynCv0
lj49/tkfbAM2lvZ5tbix0cE8H94rDop0o1lcmMpxrYzx/f90ubCB8naRON3vMxHICV5UjjnnNbhC
eu2BYesR0ro1Re/JTZilILH+FwIGH6mxMXGK1YAX2HcqDDVgvuxgqmtgytYPMT3jVbKlexr5quhZ
QHhbLa8AnCuypPM+2y44hWrGMC/+HkyFYsHODMpinJ0OGhpLxxWmTlGEDW5euPG56xkg66kxtLYQ
FGcxhfOAERaU+gt0d1VtV3ZWMQWVAsWbbkSByBI8TAEEmD7qBebpyoGZCWh0c+/ZHnqlXY8o5J6r
ufn+oqNaJMmahHp4Aor3iltd1YyHJkDXG9/6pDGneZB6j07Jy9ZQac4bheKTaltvNVBF/ph7DQi8
/+yDNSM0pfZZvA7Pvz7QwwsWHG5C0MOC1g+s60Lt1t0Fe66ekw5HHkG+lMjVMfNjjwHxSpiaEtrM
ZJevwPNX4s1oEMTsU+4H2RKZ3+ieO6oBUeXgoMdYcKdI/6Uhav8rCqZuqzdq8ERiQpz/ebeh5sRt
j96Rw06qlsEb8vcoVZQU3GT72hyXZ+2/b87/vajBu4uNvT58Ds4yO10RtdAX5pjFWB6uW3KnI2VC
LEHDIItDhqP7o9kQuHd/QLjXFERIGj0+ZHwssTX5Bhokl2jwqHvq7u5UpC68R9fjkRTOGM0wP9aZ
wbSxzXEk1v/tT+Ytxwrz245EGCoioNBsNCTQcrxX0FAqdWj9991Uu8lrsC4jewHc1IkMvpvTEBqX
ahv5+8O6vjyhgz7r/yMiZazHFHz9AcTTcQniqHfAi0/Mt53p+K7cuQQX7e7kZSnGfMIDumOYqRsC
EYsMK3tSx1xV4khvOSa7g3DqVJlaUa6GahVCFALYHvIrKU+bjEGlED4tUVKd76nrcjhCHG4SqIhK
GxpTLjeajTxxjfgkm8HrN50PEDkEODL++7nX1Q/aV1c+IMqGPmgIqkL8CG1dUzoiQcuySBhZa3jj
xo8k5EB+TxtAbRzjc4bZTNW+BPqMRndUx84TZF2OdOB8bwHEgeNCkNML2eooajIhDQHHMJ2yAcvj
xq8gYtJLAF7zdOENdqMBC/z0eB7JyCfEpIw3V0lJywFTbFBA+5OBMzSQ+wCpb/twXGlGS8+60J1r
xfvSGeidsKgRHQyvx62j+rZMn4mINDXMnGm3y8mb/nB1ZewAHyiXtAcvHbGnjNGQuymybZ6vpPpU
9uAbd7kuHbLYNacGYJulkoB2Hn/U9chMGPmu2lXaAqDQi2JDTAvgo4GjMMziHsGOlh9ArJlnyH8u
kLU2j1t/WB8BE+wx57NR7nzbUt8TJvjuUnle8yrZPOX9f0J23i/4yOhn2V5q9iyY2y7VmhK6hTFe
LLK1tVVm8gqAoAiAt/ufaOsq8nFH+gUs9MiSb6/OZuwJdDetaa+GzD5yEvgi4PSkmOXQnUToiCwj
5o4RtTzp+EvXgyy/k4+YHjtJeNY7KC5aF/yNvmb6CwViQPQK02Pg/Zxg3Qj1xjL3h2eDaZ1LIx0p
YlzPJTY0CFhvgJRRsS238ixKytByynWwUt8S1KvTp0OgZBOLqQyTgI80JR4zSU7z4WSEerHx7IKk
+1LWM+EI52LLAXAG/p70Iv81fvcDlyfE13r8/MWGbmJ9PrbiQhGH+unwIRQTyVBxVZwwBl0W48Wl
g0QFeJF2ymEiPZ2slT/1WA4gbnL37jhM46zprWJUQTaRFbnpV8VVmzXcgbSp/QmImP8o5IX5MH9s
9gpdJHjOkWwfDnPFqrKoKgl5QduDKMDRgzBaNsfxFnWcD45VJLxta3unaX+BDEqq5cH0d4dr1u0w
BO9MzrZC0pxiLfmR5RE220z2dL6gstVi93fzAc8w0P/NYN6tiWU1oAPicHbkOI8qumu1H13lGN/X
baRn/cGh77VffTHskfBUK+hQ/CX1EAVykQ2Kw+GGtQTme2uI3Wv1riaOdEsBfqOZqKs5Me+DUbGh
0nOkNiVJk8Dq62FVM+aEOz3YWj5tWAOANZB/5T9kfgAQMelk2ucAFeoGlRWc9Ga6SC5I/lgq3hPM
rYFGCzdL2T1nqrnqIkB2Btg8zfZqcd178H/Qf0aVw9T2CtXJ7GKMUaubYYdrDzYU8ufW2/N2UCsL
pNHe3/88c7m3Kv9BE6r7ZpsDRWZvRvkpLDrGl7EwLth30qz7gEBklE3TlHdRB5hEWWTHYzz16ffk
fUxLPmUmfAmJb5igQndbYkyrG6dvXRVLfb80lKavh5Ib7lXExux0QmpEw4ruVuK3Sm+Z6EKpmfxU
1IgaQXfrGtnNE+JGwVljkHhWNBtqOygjBR2pYMsTUNGXdGTdjJoh4plMYj4KAv6Li/aJDdpc9I/k
4y57WGQDqE33vMeODsbkwrQwJyGUfC1ksJ1da/spX7h7LnoR5kf7R23+80XPUgcz91he+qkabAqt
DOL15x4PcDSd9/PBqQaBfrhlnd8/pY0z8lSKvjH2QKqlrAcH6EPmQerdmZkQB/gK3xqsfCGgVjO8
scRMbe8PwN++pk82/kQSZkJLwSvWOMU6ptPH5vI58qTy2U7xr4NPk+edSbAipLLEF8S+e4ksLyP/
AGAYMCxV1z8qaCvoyH+uFoFmbaIqYlIB4RGJAENGRy1f3nt6QlCAr0MxG22SXJo5hJ5xsHVbbswM
NdecYkXYFwL4eZtqYrxGVljbExOjODcJpTw3ywR66xrpGB+cpuZvj1xFFTvkWN0ZX82DmHouZdDQ
CdeYk0oKpWNHsMwnB3HCCohIaVXdKPtOyIkhBr8dIxMYocMkQTse5LmVgZrMIt9w22MgSSRj7qYl
M0E8hY7el+j0nNTKPZ7YebUm/QZY90NboEKFLWhGtiIKUS40RCXZZD/NXyFpxvByST+iXs4tTGdI
cWoDv8eKsLJ3KTatU5tdeJtnhpbntHO98EuvDNnkP+4GezrJHv4JWgn/FXAocGGuv2w4liZzqGlW
9bWwiaZqaWnW+8KUrnP9HkV4dJOGtS5/+v7HvGNe9prVZMVqLpWmXT7YZ+2mMii2G5x9XoREGx+8
vTNqE4A9dBlnTmDzL4kuQZJtjC1LQ/OAQtzWHLeCTmOc/CcTZnX6wE1C9YmMSYV9StgFQa7s0BMG
Nx7woqFza9MW5aqAZgg/NJJNwPxAPterK4wB2UPOTJRtYFKTGWACDGfY43lTFdtCYvh+13IJiPwv
X99nZKaR0E2xo1Y65evfIiI1nYO6jMHVKuT2pS1MuqksN7AiLMA7FMI44tqWE2nACMhlwrze6+Ry
8jE20FkH01BqVYQzqYouOwF7HapokGwEVaJxMiyDrAyv/P9fazuyLDH/FnyyQjaWr/a+0ecvm4/K
VoqubmC2tPMHwkm4Fi7QtU4Tr8ecJWzersbMXBdZqs2jg7n0xLutuDJCF1w3zha/z/Nyu2Scnd7i
1nhv5ARQj3Y/4coUt0hgr6uueFd3/NCC2uFL7HOUUfkDpDoUVFPnjBZlHw0J8WafwRFkRI7I0Vid
CTn75iK6evx/Pl7yRhMte4Sco8SabuO3g0mAd7N7U2Pn7IEtefjUghjCkH/s3sVkUa5vn/l5vFAm
wJZ49SVvHd5vRZwrXDPi+1IhksUi7ikdT04XSCX0Pys9/NaOtCS7l5RRlDn1lZDG4RjwApHL92gM
h01i3W+EaelfxQ3hr+pH1Zv1SKVDq2UdJGgEG67CoGReGeBc8ALbNdsH5H8eaWYSZjUeQV4+cHzm
HuK0f1+rMffHKD5Ja/HRxrEnB1RHnM344HeKza5x9qLlUb2mZeDBNWNT5695mFrpDiOV/DEKmrrS
oKYk/4JStTrQTa9A+tmV8j1I6nzE3l0OvYKNoMvruudmjsg/d/ZcY90KrXUwUw5jEkets2M6mbCl
ZRnbtanmbEAlCiOL/g/t9Y4/ZRC8C7DbmX+P+27R1TcmcmFe5bsDj8Y87oOGO2wcZhB1W33IDjG6
9g+5cmBpa2zzGd1uIBw95kwOTFjw4qRoLJ37zU4+xETsHG6jlVcm/C4SySnZAb8ySnY4rv+J7gup
NWrlIDdz4nJWoIonhCQE1Acg1imcT0SBqNtLqUFAULBmckjj/rmfoBSBwoEXmwMOSPtMrlJeC8L/
r7ZdgpHoJYsl/d0SROJhASCaEXibhSjk6Lcgd0X/HOLJDbJvlZRVqhQCAPw4DPoYIRLt4K+4DUFc
eDbl6FmimLs3lha4uOO4RdRuietRYfmuF2FaPYysDdBZ3UBHXL1S0CAOYwOIE+HZGhPQecVhPz9U
M8JgVceCLbDI9TzfsH7OBgxeL8PJEJ0ZK9onBJJByOnI3JVQgvAn/95+DE8x2XgCHDEH/8+PLwEt
PwwmzaWdpFWXR145LqM6tz8sB7QlqubjlRwDn0VNS71t377m/B4bJELQP2QvK4Q9jmzRfCGWV+3P
+JxPE89Jk/Ik19AlctENqXdOqU4gSM5KFb8zLZXl6KoRKJUjbiR+v8uMUmvITBX1CRV4p6CNzyNP
2qy4KrFbhrHq1JgkSWbS+6PTS9h70qoGW+86An+uNQ1YbRXPncHuxYOw0/FaRoQ6qrx0CVI7y1TS
oT1ORq8mb2Ejv8wWm3i5n8S7Phz+XxtpxySajAbWobGvn4gsuMgbz+gHKAXaFSMhlY+MeowTZMha
ArrXx81mWEYuXtpwxNchQ4+S1eG4BBIaA0ZTD+PZM0/PaFUtBvaFc2z822IUhEqnK8gXwBbafWe/
H3KAVjTE3o5pp62bgQt1j1E1KJ7sHFwI+D8ogdVHzom3V0ylTXT0phQwODu++aF3ZAtFZGOqhVhb
x/CDv0p7p9FLP5ztMmFPP6hpQrUXkyEP5KtqKvooAAnLo0f0AmyDrlZDbhWKAZrEHG2f8Suqx0pD
hn/UDQvot71T5jTDiTXJs0DXh1dxWpdIXVnxllk8AKvs10PNGtfimm+J/EDwG5fYQJSENcIFmjwL
tVzPZqqPBr4J3htSM6kjqSJtg2u+E5R94ofl/25+X46gnHsejbK/mFIO09DsoP/lSy0RYUeWvY6J
8yUAf+l22xSqMbGbLX3Q2MspNQP6abCbG3KLid2rNDxkQfe1xd8f2ppLmhkABlsp/pQnWUERmrkv
lVYDDL46JOYoCZh4d8Ebi1fmzmu09KBoSliw5mTarWGccehO51Hfo4V+JYcbtk3RpnEBnGeNl4P+
SjeDotPu38mAv9erWbj6LoEjNLIfcfDEATkRzkYxBc0+Yc16bKQHynQIq9hn5DLKSJ4lsx22k3Bk
r/ivEX/KeNs6iPPjlaDPrBbiTZ0UAiitC5P9fUQua/1qe8155nx9chRMXw41aq4+JXkBf/5xA/5T
kRG1qYRJ/PlpzJJJUEhUJcL/duAHdnVLCY9IrYJ5FnXf+ewOu7m7Rmi/f2etPrOtagwctGJqCeSC
sh4Unfk+I9XHccs0MPZage7fTE7F70tVZIA03luOgB6zx9xLEOIB5vbrQyyBFt/9ruBuoa/8x6Ze
zVDNMgXk6TyFLP85sDZ6Ynx9QPQhxbaiJTBkSgYXMhdzANcAZFDO1RERIqWsxjnte6rJGzILuLqv
8pMTMo0NXDouwXkSAI+vN91n1d/xCwCpvcfFhuXubgKACeAlVTI/vOIkB48jCkoZxYDDZKW+tmIX
p81ylQLbjf1MhEpRG4Z+LKR5iBBic4jFrN5YiH8C6hmuH0XkLp1XQNbY9f4x6c0d8o5hAwRB4k7c
AW/vnBC63MxTYYYzsY8q4aG6sSVa2cfrXOCXwjLoLSl5wHjgUzxNWCE9l0F34pJgdSzsLy8s1iRA
zxKQls81TT59TZ3AiTMwd3D+7q1txLr5p2rj6VqF4aeiiKR60D/reh/8HnexKc4clMFaHkUdiNAE
psADlpr+hceWXT3ChBWMX+0NeY0fAhNDPyIYB747Bbqt+Jm5HMD3keWPmk7TmH6CC89YZcHzHRYT
lkhRCDADXaBRkooc5f4CrzTvroyZwE4O6Zx1t1ZQQLj3uiAtyTptCgtTSS5QOPBVm3AgP2CbOyxJ
+3YJLEygQ3wCMSRaaalm/I/Ea5y7j9d1cITu5tP2q4Mt6ANRyL7n1LFajdxPbO8MDDkyrXnQvJB0
dW0dqgNBvqXOo/fLgVy/K3NRd9Erix42xrZBYQEATstYCAlM+5427HjGS3lv8pPTo6NQsRdxg2WV
7oPzoXBx0OrZ8rbWzuLHizPh2EAm4jB4VcRoi0Q7yFbWjKZIiOMnuulRxDyYt1d5HX7VkhxR6rzd
Vz3Yc/7ojwYuhHCvqp+SgSPSvOhOrHPLdBglz95uJ7BgaW4tekQ1bQPAqoVADmzfSEKGdcbCvDOW
5J7YO4Ip9EHHUM7G8RWqhYQQVU7CDLQvz0VhJqoxQ8dg5tfYdJKZb+RteragEOOTbHxWfimekVXs
I1N5lNMlaWel03DtGRbukNaYZJ1XgQ9nUqT86JE1pGILtt1yefuOGzRWInvYFUMo+W2+YmOOXavA
dsrYs0sSW9IAw3ieeAtPhjR2gutJ/Br2fsfkhAdpKHYKBI0W9YGzSARDGJq9TiokBSV6P416LUQy
HGflN9SIQAIn6CZVrh5O9b71vypUO/fczOkkrY/iDTqxf67wDaD6a+Xywbwkd1oLdEseAdIrUP18
PVwzuwXvqfOBW5lFbnNOOFhRIYvaKT9oCzPmBWWoOQoayYiCma9GmTzxJqv9V9RUEZ6PVOly+zPE
BIGkzcDESg8VjAXLb0A9ioSRzPWYngsy0jH9uJZO6ABE3Dhs3q7Yd4b42A0BvsLBiTFWLSkOOYXj
vH+/dagMmm/4gAh7RY2iHdF1aJvuKs2iHS7aVTKHNi84Ii4wGROOgSd9LtVENfuMDhOgVvPut/YH
PscIOhoU9SHuE8/eyfCwZDvZloQN70zy/uvplKp+Pt6BeildWgWboMxkRF133kYW4MIoGda6foI0
g+VvITUh4tI5VsL40uNYIRhJvwbAjrO/C9R01UB7+YpUZDCxb9SznUOJirZ6ElfMiv25UyHIrH0p
2ymBHtQMyYsYAFNUYJvV/flDu1xYN8ZTuawZZZoBjvGC2U5gOa6rotZQgFzPBZAeyQRCzJqKQXHc
Sxb6S8UMvxI5H0T8XwTZ3nlpVUW9yO8tNlG/ddCl/ugs8NmOQ3u7y8OrqpiUwXtbk1kj5f+h3pGC
6WkbCsya1dKETfv6Mr1GEZgYpJTaTdn24WGNa390dCtaioHQNiKJw08FBc2RPjVY5J4hZKxWPq/h
W+/w8RXHQhNAYjTgPw3I0LG0fS/b6hQggEHdbRpN58RnbWl/tdr1iMqOe5T72sHvbPqG0stvIks7
l8GW/DclrmbiU23U9YSxfVNpcWBm9q3P6W7oxlKBzc0bSth7RQAFKDe4oEiS0cZ/PZDAPvsRk5Y3
qj13RU2Oyy9X0uMSC3M7DBxjXJ2uXYu1KCxeEtd7stm0CokE5tURLHVTyO/2YW9oc0WZxp/Sg95a
19EqylcYt402I72YM0vFzoWF2VuXbU9+27T4nuZJdjkeUzuL6sPcPmRygkvn8vEaRP+RZbGgqiQv
NB1nrMJcqySFzB1kFQs2dtR6Z/riaEQFBoUTa/yAAOaRx0GCSuyQLAyGIEVhtdfKHsxRybLXHwOd
h3Ut1EtUxzI0nD8eT7wdvf+pLt9hhsMNR8YnvDXKnmwzWeP5tGFn2zH7OQuD4sEjz0yATF7ezDR8
cJ5zgHYF9VIKxaFEXMw+QTddIbnY8x+vsZtspgbAM+BWgrFuslDjquh6iP6Cc+xN+WW0h+rYem9z
C9hsbqvbElrNayosT2cP+gPOJZ88SAmGPk7L0ieYHTXSwqCmBgaVVCEzOTdbrazhUfO7wBeG+Ky/
pqafz4bpmZjkGCVExXbxp+6R8VKQxMj6Xa833pS4/15FUc06BeGmFcoeKubTWHgoZlxtDPkJAzOy
bRiesoUI3ucTypC7ZUXSLImFy2R9ykS/5RC6YSkPAOh0z2nF48fJHchxR1SN2LIp3vLX1u6wWrUY
l9lQQ1Ex/b1Qm9MFdoR9qSvW7H8qG6NbC5EYFiJ7ztvHqUe0Iy827lK1t0XUfsfkPIhbUR6jRwhN
dDgiSadyYBW5NRj4Pd02XtLhIg4ZotQI4S33zzvIoLaoCnyNvQSzCZKe++LKafGCCUvthKXaFkJN
lOAoo+V+hWBrx0IuHSy9r0EBSnopm8giDzZ7uwpJVkK92dOaVMNgTmjJu7tKYcUUzVVQpOJ9yoQp
xy9ELKwxTQ+JWlHVPpBM2w8QpQIhSHwBeBc7Nfe5mZ2ZBbZTEFEEkIdHdpGPwXlnIY2H+US1pCI5
EmbpyRFFfjdSoJIYNvDBTmPexG6MYxXS19jtsM1KQ47Oh73VseJWe2xbzmbUjjVcVS2nAhppDFJ4
XmUHRaxAiN6QjKpD4uXcejSB6vkitB8Evl0lMr3pJ0QYBgtfzAbmR0dfFWjFd2TPFBEcosLAiPsR
rp7M2BwENMmczTM8GVUmwFneqrB4WMro5D0jcQwSzVmDZ0bowFyVBnVcC8U9feq+H6xZ8cHAuXAr
Aw3NPeJfQDTqpbm+uZ00zBgKHMkhwxN30Jb0px/4eUgCThsgj8Xn/1I6JyjXzgrp18Gq3+FUpCQC
8ITB/Xb2WLYdnFoM9WLhtaIfZwLbT4R5SD53un2VoZfJYoTsknSctqqdC/IyM6xWMS/dG2mhHjda
XUY9l/judqEKYih9UTqF3l2WzEbdhrIimUwItledAlNTUMCdh/L1GFO287GOow8qopCqkI+WQUCl
Jq4Laki5GdcEMit7xMf0Q7/mMAuizYKine67WoG6q2SO2s5ra8Afw/9yfRK+tNEkTOb0nr+i9Or3
7xhbGqbiv3Odj4Aaq6XzsFXJeeArvNfzhqBqGyYnACPR0d/1Ngv/GSpVNJBmjsJ8SsWdYDbOVMX/
tBxhuQfZDApiL/HoqwBjL9UuYVWPSsbVhdtLtXVRSkwGmqE2ZP13ePhEA/J9cQywhsMpLIZ5BTSf
YQS84nzxLnIPoANGjsGR8KwjJLl9s0m4b4fxg3d1s6Z5rgegseAUFrppsvuMebWVZmbcCJXMM7jf
LYEpzoCB63da7Zfb+s0wOHcY/FI1UUvKFmRv0Wl18FHb1e3J6roQWa9SANg/E4vNkr4t0JSgfm+P
AVMB7nGELWZkHOhI8QNeQzS5xGCyFRCOUsU2mGTr68MuTqoDYQDGzozTo58kqsbD/VZrDNYhU2Eu
NB+USmtTgUJlMCuW3QkwlkAy3HnPYjuOoobPyefi3FNQQ7uq4utVE3Q/AqZ8Yt/cBI1Roxeb78mh
/2VC7J2qCPUTftda62kID0KX6CwaDxpYPXg1Ivvb56R1k5hQ3myGQc5oYyNMKxLs7m5yeVgqniTN
Yu/sGBxO+nBI/P5idVo/QO9DjlsrUfWjhHTm0iFV0u8n5jvhcFFxOS18fygSAd2z2t6m8bIjjT8Y
AG9vlWuIIA/Tx0j1XKRpwaxJounm2i8qceab6JXp0pS5rx4S+YjfAVP1obvL9cQn30GTJDID3vZf
sgBIwFY7hqOPdUf9BfOgGtJalWovBgFAYiCL1lqxKoz4pavG1rjGIyknomPag++gdY3w/IwpS9Ay
plG3tTXysMOEEddcSAtSLpkQ6lEbMlDSd0iGAJ/7j+w2U44E+Mf5z78tNgvCAMCE8gFVhrTtbilo
lTbTeJWdYXM3aLDHPh7o/AfFq4mljTl8PEKX3+jg/9IzFvfDUcl5puUyuNpIlFewaHAvTmIOO5FE
4Zh3848r3rgS5M7mRz9Rt6MNAaqWlS03QNGoTqCxJnQXtOG4asepZ4fvSHilw5GhW4ySEaHpzi3E
ARFG+PjzTStyjAUV9AJic2AIseHFV4JQyP4gbS3lMcoJEqyJfm4rahn/4ime+U/eLF1BfR/gQ27Q
UZwzLss6jKcd7DePH6shISoxxYsDnmq3lXbhYzsiF5OxNPfRmuO9XsO5A4T50L+4CfYb1RSPUMWy
JEZwOMFGubZGFGiYNvHv6+WV5aoZSmaw/mQ9mFZCOL+rYSwULQRPGH48ur3Jd9B5wP0luEuwaCRw
B5KpCsRLHCZtU9W6JypUoICFr4+hbfLMSYsICsykOUohG1GGRQkiu4ssDKXfXxYySmjuO9oY6dEV
NGBxHVLwspssSVqwcLk3BQMP1QuFZx83fFypPlhCfX9p2J/8TpgpX6a1u/Qs9VJG4L3Swi+fNgvx
GBB6XoHNlKWYEDVxtIcK1rcJw5g6K+Mu9XVSUWk9tkT0x2TYSFJAf6ADlsAzK5RpnZu6GXg+1vgV
88PC1poc2ETKavQJD44Zxvo+DTQBee50+RMEQ3i7df6oHHi6PXslpGGsEXDHZFOB9JLHkGzfSclw
CaHbibf8nE4b4VUckj0dTNR8sAZw8iTqCJOdT1HuvrcANQy8XZN5sc17qc6JIUf5jTqPAM7INev7
+qyIzVib3/97A2malbuNnqXtTuIbNF+wokeoH4o3BM+MlelgdL/rnpgtKq7ypgjxSUsiZke2uJwD
ELIWcwNxx8ZF8kRvvqKkrNI9IbwsjyiBY4EGEDLDu4sVHHE3guN/LF7D+f8NByOGXJQ0pk2f6Gos
J+QF5U6L6onqRy36FcDT2rfdhkMwICK+vegx7/TefLx9CngZgi2R6k13dnLo7KmIiG5WyxpVs8UM
Dm0XFq32ihbHxgOHR+l0HwnjIIBRLHdryh6dI5kyMN8xbgxPWZrPkz4lw1reRtBsPm/PFlof3qJ2
WwNwBkyhLHa9EY1r4jgUAPGxiQBTcvrb1LuLYpRF8xIEeXMsShwVHwFpBlsIIWoj3D+/WTRteqqn
zO0dkFkv4U2eGN18vS5RQ3QwPWuZbG3V5EKxVyYuAHt23SV16ayMbeD++G0xhEvcuewo7xChKHLS
pL99FOxAsCryvqtVu8ymDC93ndrp5D4oMaXynvenjtgn0auJRo3r6MeJAf0uY7qVJWceISlsepR8
JMvuSBpsaNfa/SLqLyEAaUjQb/MpoEkbNYzRf6Q7dsLdNxaCHfAVFOO2TGxcfQnbfAU22ThAikvm
Af8AyjZ3s6FLrRYlhcjZflbEKoWB/Wdq2YRn4COAJub+OizltTTAMuwNr//8aAM6/6JQm13lNCzC
c+7Ouv6zkFkUcMcC9EZs5WkpxoYPhBqycX6KOBlGrcy8pp2I1LvC0o0smMDngeNJ7TJJH2FU1XLY
E+KL+goRmgJAtKFqzc9GEFgCrBlYA6od4Itd+viigK3flnRZ01y6ixV3+882f2sznCnepFILqvId
BhZF0QnkdmQyASzNHpP+LNNsrL/eaeMg1Q3lYKL5WNCW4FljjZ2N8rczWqvmKaCHbtlu+kCkNzM6
zCcr1YlHL0W5nLC6nL7hzXdKH53wwLerAUZ7XsnER+paaEN6KJIyJXa0S3Z5cA1ePAwwQHts42uK
oK6G+Xnhpz40D9mfxjwYmO3oJJMVBZUC3/t2Q4AzytXqOn/ZjGoFl8TbUj1JID+Ia4B4MZHxfALI
vGB/10Ngz51IBbj5PtIetbydTL3ALVrFi2s1FxoLt2VGquxRIym6DdvoDQCGFc88jxFBk+Pir3F9
x+8r8V0F7F9PZq6+cPr/9mXU7S4fFjS2sDLzzxPL6fFSIiZXmf7c1dyJyLOF3XN7wkpGPIZ1vMSQ
TeM6whxb1OV9+9UrbIwuUZwIEX9m99g8zy1cM3OtdJ3EOf1Pz90Sl2NyyswODdcEZ8slIk7TLh2v
3ABMpg42rDbOzY+06WBwbeZ4NjaRebjTB3NGmY13lLfVVXnneBT96IlIz3pQ8Vyrph+SOewzOmEp
1Sx3/TzxgI0XsJt2Hn/7U1r/CcgkILyoHpoCOAA9y6/BD52++ixirfJhrgPKyYSzPmhl5kEps4J1
RzUpzK0YFDS+BkeT+a67VeX5Mq5VP6RiB49Z8lysKvgqMGCSWIiZRFTEu1/b83mmwkiy+O7vZT7d
GWhkOeVdGSQTf0wgjLiKl5Mnn5RQtyrNapAcm7D7twv8vELJXwjDTsC5xYb8lcjHwccIE78MSeVi
Dz7OYEXd7MZgdD2YCAFHNf3Fy1pYEpPS0u0fiwS5J+RqKMA+o4HHEw49BVLw65I9Znt9FGslsoBL
idVj1sGXruPXNbYQaQqkNkjYvCbDlTLcx9eug9PuQb2FsET9VGozt4aSIeY36XB7UvHtwgRD5bIn
8rPXDfUwBSZSiq00yZlM/CK/VhxoPp+eYubr2ud/J7uINYEZbUo9MilKllIEMVctkz9oCYcLdTQg
x79pwKx/WBpfwcdouy6nc6ieNd7yRHWjAWyePx6KWDMkjIsVMZvtgXCaMEe4jwokDgsMh7mxIaUt
wHeT0/ga1LLioRc6r2KEwZpb1a/M7QYLoU+TLlE2Vmdu0nOrCTafQoIHR0VJxji0GJSfDztxyjY2
+FtHkfcv7aRxnVl9nSS8meJwWibH2hlP1uswciXbfAzoXQhqGR92uBO6ywHcdg9JXgGzVwLbylz3
4rEeKXWWM+gWwZt+OqeQ5GQ1S84eIGQT8QIr2oazAhdHx8jE4gRFhkMPopuBEONVLrNXG+Xera18
nK+CQRpNZ8t2gwn9AIxYEGI2+jOZMljEbyuuUudJqq6nuqoFwfyzqunFS1L6mg6zr8nnN+hPp4P8
gqVDp6eQuMOtNEa+I8n3MWMrc1y5AweUEeGwjfiUOo7JCbtLWGVx0MPcbEyZHJ21hS/mk+UR7nKj
xqy2AV2OwV5LEEEeLmWKL7BvNdpzEvBCjn1mUfvv6KNcJ4kKXX9trQwbx+CBuok2AlhkuAKVZL3E
6nJdkENtSvjScTE4Kv44jyd0dnQbiXeUmnjZ4h7Hn5mt+uEK5cL3WgKpArcPao0Z6QqTC4ZRvuBm
XEW06WQ1JDT8C8B/wldC9V82mMjB5g25bAAvc7uc1txCQ7L79w4fslIqhHeyicpMwTjhBWbdT5Xk
NA3tLAgVqfpVUuh7zdIqxT9V0ewR+oZeRPC6MCZsSEt5AaZwQTW/MMdGFVIF7mQYxRSBu4tXtPS3
nNplpCilQzinnMb/4gUtrgtR67zcNRRugoRSEwnZphQoT3w4308uFaBQLlE9yQuh6IC6GzcjEK3F
h7yMVaVyfPMfMjGkebfyxRkn1l5oOAtLOtS9oY5kbd4CxjgaMd7rgk/Qxyq67WFHIPfnM54i+SRU
3HzbspOGyIANDuHGKBPZXs/LxfCfY6LCVTvCoLv1WUK2wOxqo8CqWyDVe4YbOqmid5esl1oLXid9
Rb0JtMDVFVFMA7krQnQNiU9LdByvzP1LuR2uM0AoYyYKv++UTOaVbusGL8KdRuRTU7Zt5/zVJaao
J5bVfy8WiPZ0N2eHuUhYU+aD+1towcG5CjUhfBro0bK1ylAOiKeN2WQlHoc7/4hqkwLu8PRrWcb+
u16WH4U/fkfCDELAAeOV385VwfsQXzGRJBdJT0RQD1Ni7O4OWgDro6YfLn3i8LiReuQ2fissbhmq
L3FdPDAYswRWBkIk6i9dM1qk8FAe/a++zLwZDZJPW1ail218gwGzKQcRBxOjcp6vp04+72IFFtaX
2F3MWPga7jHGXu09aI0duA7EjLVda2ZSG7chBrtyG9NMeHMy6HEpdLQeoR/u5VanTCQFAmOwisAq
p+mkYH8QJSUTRSqQuiaaUedz0BHHc66AWp87taZSiFr+ZG3ILDz8MEMQxkbfVJ/eX0zjMnDBvEl9
FcVQ6DaY7jX53yCe+zEZuhzn1sx8YO5l00HcKnwEs9COggL95MTLQdqY0uLfncEb/YSts9oSX2/H
cCyzv0/bWntJvFa0XYcZgYPWQG4CcImDgUxGRm4UvrDCSFK9J9rnYui0AQZI8MYMCjkk/d2Z/AZh
9N84pV8P55f1WK9+2KQdmnmn+0E0kmNgmHw1DqCoy86RxnnK70tAasF8Q4rQAsBshh41NtATSbES
EoPGS+T9yntJ3CzC1t0L1jlX384stOGT+/Ihg25tDvAFWTMDz05bS8FCTkVN794Y1FNTaodC4giM
Rf70voN0pfhZJgaUAaCU8pvv9MhUZ08siYNr6v+IeByGdZ06efot80cM5vzjMONFUOAlBSWWZrbv
55gJ5Kjw+tJOBFQfhIu7hZ1oZ4P53TJkKymaFIm9bUFQxoN9QUBa5/Mj/3vSf+/rKof1unqaFa68
t0Xu9UwA/lYGJscZ8GO8STs2xylOqv/hCCNp5qCHvKzkZFlIpotDcLjuJefkk3dzV9HikRg0nQCz
rNuHe5ziFXBe5NDzvuR3cs+laEJrDGC1VwgSkz+WUXbSlm91yplsrogiWCzqwJNrIJBSadp2F564
TChsd2WbbVJd6/S+4iIaKlQ/KJRBgJjUH7unhv5zDbUq+nOfd+KSJfKv8w1FjmZQykMTiHvkbp0H
vzWCiBsw49XBAQk+X22+a3fk62yKENN6YhiqG/g24w446zsYwIqRRkRdgvD60PMln9b3TmVd5Wo7
pnFzw1AGPinbOz6ds8zBN3vulog+dkG5BO4hK/8DjyLUPikxLAsZqN1ctkud8iWCDEnbpu20oXyk
DhIaQ78hI4qTkfaY/Ouh5/7DvU0l+JpoZJyKc07D3eVMjznfjfu6tCxftSCig9HeDBtATLEnysHf
xhV8vM8Ap0UKDqT9FzVsruRfZGn+pnn6iA7ruSZ4L6qP8nwllGD1fgLEBIpUbVHIUQD0tyAQWeDV
mQTA/8Dm/vvqOmLs5FNCyNH34S6LLF+qRaeegcPCjgTbnFUFnvGxEvJdlHSYQp9jvKI/DbkcCJF9
DCv7dY+ROaGwiQRdMjVTGq12cVfnqWXCW+6QTKnHqVfq/TUbjHmuYxGKfMM5X91VbOJfn8d3iW5Y
p3UYZ5DVp4S7OG9lKYWNZasb1bzBIn3VVPzMxaiPvU13W+SKImrfFtzHpJCoi0JbYuQtlbt+MDDp
BW/GEql9wXX7PTbY05d+BFWaqdobKL60k4GSkHpA8/UedtXIjMDWBSvrxRo77EZApBAQmaOjjPOo
b7D6mL1R/ZrCCSiw+Vx+JpkNTZOPDMgbOHkeQUFvxkdX+n973jm+9SchyPgutGDRMzJsjcCVgbhc
eMM+KMCW1J87IgHFQWryT3UVBRJscxBkipjLHiN2VWOdbeXbGlDqWs9bclgCaD6axEFBu+mEljPI
+zBjaaae1Kf/l5LA0f6aaAKfVHoQWnVIIvphUP3V1vM4rqAg7EC+yxpWJ8FvbupS0/0Ex8lpuwBL
gN1s6eKYsCBOX0B6eTCBc48P3hHc2QYYneQesLMXZkzqAc14LbpFiR5MBJHR1990Kq0+k3QPvPGl
UqRL5Vo56NlabTpOSkJvDAw53lvJvQu4s54pW6cbhD/WOqiWvfahe5iSP5A5yDOhIpuCPUbETGdZ
5b/0e3ZNvjTsgrvJTKkQyzoXQ3jMvInXaaaHij3T2eSlDHnHrJqNYGH4I0kAHxGQbJfsjzI2PZ6G
LsFC4abfNUmzlHR61xoCUlmU/NDoPHECyAWjlDHfEWu65najSqQhSl3Oc9x7mWUUmWQGXzggOkrK
B9fRnaVpDCqbzSLfaH4nZF6T+y0vBmS/nXkWiPU7HPsY0fths8OUGGY0iwTlJM5amyN7pLckzgC4
dARvWucaWTCZSf4YzKTLqOQu7V6NClKL5HhtvJtBxpea5XXJU6HYKD4hlQEkoz6pl/s6BJRntop1
fMVX+h+5DxAj5DfneRpqVH2PKvahHyEHcoV44ozpPmeXPNu/71uQ/7AcT/swExolszuiUlnd7JQq
QHUSkcQMg4aTa3u75CYElp0cbtpjTCwxk8K650sCgSkxEZuvj5P4bX0/q8PlRojq9YsHiSg8cUFp
JHaRiEOZtXm75jkKgWoSA09jQKNEUcKYDBoLrE2X0g2FbtxFW+25uar/enZ9kXs/lGGrhn9ezFQ0
jknNDF8s6046GIFcRrbSk5dPHYqlahxjDtsvlT6Sp9zcIvRoyURGAkyzxNVriBmc0sYxgmmHswIW
H7Ac5POE1REyU38dqxMqIMyNeaH2iZg4nWvngv9HLXd6cbhE9GtchAVUamSZ9dOvG/6yNH6NjsSL
eIYfYJUNCStHvv1+/fedB0BKWRUU4JQR7cnss6wASc2m/hmMpKC+T2plP4PrGWBdDbkSdHw/5J8W
uUoYjLo93Ydnll2+FRQk8mbkTtUZwAg6vO1DxmBDKiAE65sZBEcGEU/y7wgpi27xm4MSyE6SxG/N
nSFjJ73ZFtf8QFShV9jNKzCu58qWUt79XTjcnAjEXvrZwXks9LWtSsS7+R7C4+2cOei8wyApJ0Ht
iEtBDTcflKeFccIWtoRLS0S9Ua0VVUFnrufRSdKGu/+WGynIFZNVadSPuCsLoua3jR4Vqe2A6Gks
FLW3qryBDK0f4A69OISvTu2g+SpNZN0WeGGEGohlQlP2al2kItsq+C+UnVJEOzl7B/ikf5Go3v/Y
G40nVzoB6BsLMqGVvx0addFh/h4k6FVkJxzo2iJU+VxNh/6IFxNZN9V8CELn1DW2XefT7SiPw5oy
RQAePXoUGze5n5F3o82tJvB1zai+e6NThgVqPnw8k09N9Wo6hCHtAAnUSJSjzlpdHxP3wR+uzUad
ss9A51ocNmdEld4hHy8hAmr7eNVNimIr6lRGZDdU2rHS89o+ztfr6gxP5BuY6G8p9G+74TRXP0LB
F+zRHwW/avKyEcdSuBZqwL8YOj0CPCmezhS6WS3X2pMbzzgWJEl2W/yCHAXrwy6YcAwivWNHbDna
LMMHnxiax+32YjuMX5eQbfashI7wkQkDH0RUadtZHcfu8rDXmBpUETRF8ogobVmfRJGBHyLl1kK9
J6WRTKa70nHVPfu+Jmp7/YdJ6UW8mh7wFLYtXIGy0OgMUpG1tGLkcgVemHoPeM+Fcpm9BHG4+37a
7TZxaP6Gb6lvTqP+naHzwbFoh6m6rdCnxD2WY+7KTaO3iQ+xkQxhW1NGw/AXEPCXi9UuOprnhHe4
mpFdk3ypHfx4S9/u9e+ES1pVAEILYPgaNFAplefAXwBtpUaZAthfwEJSjPyBuSO5YesG8BAqZv7e
GyXHnq5hFNL8Ol6LKI5e4C3Ym7xlaBZ+D73xk3MMr6bBNMBg5R8yNO9TXp0JmU6bN3eth5CgnNxR
WfMxbCXdLtsv/akrb61XcDiuWiL1MCO82xRW1vBKplBiYHVrOOV3jmMbHhmZ770kqGcxEN5j0jIL
zY0mCSJ69MqW+MECrjH7P/c8l40Q3/kPFHfI1oQwrMpJ1KHD1K3ubOC9ArzgPFWsMBhCz1HeY77e
yqii7Fz09VCrVVZGwB96TE3pxHZqIQDDSmL4ItVgNcDn8M+F9qyjcqLAVjh+NDxdN4NUKBwIeYPL
/VfRdN2H6uM3UkVKGKZAiHki9u1Nr0e8SnomAAvNA8yW56rJfqDLTDHtsL4EYy25KTa+zkiT8urp
8foTiceALw/0jsrj6z0TVJXg4dh3L20/cTd0X5l4J9muoXvIYR2k/00lYbAIpAjrb+TdmnRVp0Id
y/vmSEPJUEf0djgdVdVuzEAR37T3z4QZt4M0t2ibD1cdj9XstfKVtJdxJW66fycOjmunnjbEvPsJ
iWR+3pBwPjWCDKRRiTImOdFHIrggDz9z5ScEswv7j1FqaZdF0gUi6gXzxP14yk74+cBpE7xkzP1y
RYHv5K7gBUJZHYlweTYZ3czpXlQM7VzOeH9k9JkLUDbh+Gw/lKP3ZHPepknHyRyCGU5Mmokaloxx
uZJ5eymERchhqfp/Eqb5qZOrCBIoHBi6dFDD170ZNoLrc6+tE0tckeeCe7JDlsdn+pI/skEHgkCC
50RAqXz/ecjtoztqce6xjyknggXHlbeGbM+dg3Zhya9LSwHqcJEr7TUaYwDmsuGaFPg1Bp2rZN6/
fJN2V4j4+JtVjTrTxjnpzPtt87qvtx2TaT3DVoJHVRnrNRBBjlsd9jMFna8la6Q3i+dbucJ4ESmD
T8CJzn1iC2kOrRpryJGA2/Fcsi+N+rnpJD0uqLZBJSJYyFAqbPPo748p5Tc4COJvcIAC2cZ2MCXj
UvVaf+S9majf1uIEr6nagqPyirrVp/tKGYLfRIOSmtgh5pPQrPzUk+UGPkTztN7DEP/0HtJyT8No
md0jkpPgWErT8vJi+iDX0RSZ+veIotCCNpvQl9WEFcyma/NkRii9PteGIXEEr1QmHdfPxDaLmmLk
k0x01PTbpe/Vyxi1Y+JopHrCplhF4mRr4rAivnxpCN+thWKTYAOsIpjVwvSjhWzaqXtmFJy4mI8R
VzqdOKnFjhsT652l4UmgIKu9O7EYwa0taUc4Mt6bcHwBbJ2ayEMfmnOucEIFI2JgGfosQft57zn6
YXV8U8me4KEU97caNIxtr2WRy44+6SYuZfbiQrR0ZJOyKRG0BUyqlXm1SfNKzGDE39olaG89Vrmu
CxQHOpf1flrsH7q+tV6/MFy6VEEki6s1czVBnRETCslNQP0I80QIMkyDUbriNJ3VKzVYURERm9zu
5XnEUPOQdR0nTxr6VvXH2PjZYmEHUuo9+o8LkJeTzbybf0L7WqRB3GP5gGje7bNS3/RR1CHbUF4m
k9ShOMBAM+E8/0f8Xx2uj9NUjpEFxhzx2IUmaf/v3bxCSWzWIxt/3H0HN7XKU/Xk+fEky/0uqMrz
3+hL0gbUrM9VoIoaH0WUK+H2mAswE5UAlf5//5thwViB1rqge15/1/tfLUnoSmA/3IrJSuXHkq9X
vFkAxaDWsHXu4olvxrtOlyaCwcsGYxBstdYjBU1k41utr0twmou+/bPvm2T2wXW3p7a5+40WLyx4
yRtcE8MOd6il2MJChvlL6jUeMH0DOQB2s7PV2i2gW3D0yjNFkCph1NIFOwXAqKQORIbZvbH9UId7
Bn+77JryF8w/4poJtv50K6D62vAT6xAQCg3YgivMPIEYxelU8P8IwLQg+HWARx2iZnw9jjaKNnHy
XOtsSoSYCA8bQfXlmVhzh4gNoVaMo9rSzXofqVr8GaaE58Lco57TummVZw7ZSb0nneHsJmBBXi2T
0LYCHVEIpbJmdmwToYBPo9YbuOp6zN7n80qKlLvaHDI5598OqLpkweac1Cocaz4dEeewQ1wL+/IB
iuxlXAW5JJ+J+1SttcH/2TYBdcB5m9AeO0ChojvkkiH/PAbtdzO4pOFLdPCQ8aAKmbTlEa24QHyb
qNesOX1iXoJgE0khtm9nMX3TnscWKd3DTZ+wSBowgD3IPWKAuS+AKc+/AI1f42NbIbR3XNi/AVR6
6TO7U6kATQtYs6z3RGsrr9U8mWkYfeepYYWBWeJJwBM8Hxb10kfoQVP284cMozCmUho/TjwfdGD0
bJGCE8sFcUezyJXgQ5/YSRkDWoduyhNq2zWoE0QQtplzkLd4hDyfb2yzjHK5nKZkNf1k593qLj+4
aCrBwS9wMjDxPA5Dvtn8N/i/hO2/Apss2RUDtMT00v+Rwt5Y0NXtmG6thhW4PhqxTLLlR6+7j9rE
wQQ+ZmTk7ct0Pr1b0W0kew5RBVjDVFNav1o1YdAoDgTtAZJvNSy582SPffjAvpkdgRbE6fO8S46c
1umTeMIL2zZRWHD8RZGsJnWDfzLJEEaYxcAre7hXB8CWIqqw0r4But04asb4w9s2UVQnmyo+HFXx
R+JPdAO5mODH+NEacJgKCinn4AxM5pXLhDNi7AHtkqFqAvwtFuIJ+mjLz71DO06U8SDibnBrYGEw
mWmzsHaMm8fyAt70IgV8uvvFssHuw5ao713HmJMOs0rP8BAKWtnDXIqK6ZqZ/x+mHtAXSacIGO4n
wcO4EdyBMOMpU2ouTUvfBETOa0lkoZQc+S3EbeVyG40hzCVag6+h8xnDLUArLP8vA60kbHSI/x9f
cZO7rsf3c6VOgj/gKbl3rdedUsDXI6Nr+6nx+UcpK4A2sD2Xnd5bX361yEvVLe+42isZ1qmYgwgq
NcYn5PyHWOCF8FtFRGF1VxrtrPF4EhnyfTFS16Z9VV9Z6EZEppxlXkxU5LD6UfQNwE+/1S/rX5z7
KfleYFwwb5lVo0nDcYgCa+oNTmMAtDmcSO/OU1zd0yebcVjXrp8ehgBsR/nSrKrhmiAbXUweo1Im
ZaTZcE0xKo/0cFwe9cByYb8UjeW6QbA5nvOxfXgCni3DKwipga+6kPq+/6KspM/bMVt6c+boLnf1
zPM/s3DEv4ADeM/417lBC3vF8H50ljXB6iMKYm6bJKup4Rt2ZyooQ9bfW63Pvmb4zGgNXySjLMe6
w3j7aV3Oj+Aw9FVFHv49dnBAmLauRtfVadTjSSIwb/V6rEaRMHetbSLk1FNK7cgzLndP2r3QKYFJ
+8qK4rsUOB/XIXO4kjLG/0DayFjSooPh1wWLYS6RjXZfz7JgLFifmaLnTxh6y/eqOHY/lqksxbI9
9e3acZ0rxoRE34S5TUNCZQd0Z2EH/X3Ss3xaQdhO35R1UbBPB2RoQtCIEX6HevsyzOQhuTU0ywgi
yeD6g3U4qN5uUkWT5w2/AOysac9yJeBHL/ppvvuGpuhKOjluX27qFfGeFqXXhfUMdp0bSz28PtPK
AIMr+S5HnhedQm4YKudnHxRAh8HwYkRRIxs1iJWvSw5Zf/Qs7Yc/Yt0kTDBeNirpkqfmEPOxpfdg
l2HEU2qY47Y/tq4HK5C184lZ6C+NxIhxdwNWTJIFyM7/Kam9MKBZbkgc6np/yNrBQ5nNkELwMCAD
XQ6PFbpAvhJ46WVUPBQ6wSh5bghRmM6VAuB9Bm/EgUv0QX1TFfHNobD9VDgzy5eQ6Id7OL94dn13
cci6yWfN+VteZB5uJ1fzRJ7ruJsev+fjg56sIGsL98vnM84ftCy3gYkQjXZu9nfgZyr9k5A3zxqR
jlTfgggA4vvM7tUYoWK7NCp0Nb3EEnYUH5L7xqsvhRDQRctvD7nMzdL8U9sJ8BdT96l+fn9tSuw4
a67uFcoose4WNvnlNsSs72i/zw3DiJvU03VF+EvZixg2cn5SSVDAcOApKbFAWn9yX3ymUSA/sKgI
nTdOouDv/J+Kbogf2qh/It2vIHWikUe4jdZFzFcW+rcx3MCYFincLsjJpdyKfGmOZ492m+uLSli8
CvXAq3y4zkR0dPDUnhh7XQMijJkwot3MW0W+2LKCS4e6A5Mx0r9G8GgQ5HYpNRh5jLp50/w4NNbA
/18W62/I4eduSV9C16NoZE6IaOlWaz7yb/EmLGu4ugp91vOAuCaqE9gwPgRbQdnMyxMoH/YEiUQd
WOZL8pRARWW1Vik4FNnFYfkPfu5wxMBiIsNrfcR1rxHaFvchc3PZNunEBP0PscCyVMcwvl7IjJ69
UI1rKR2izDcZseOs1ivooMHftpuoIy+a9LExsW16F9USSEp4trWYf44Z8XLGqoy1yCGivlT2XDxq
TEYRLe6QxhXcEzLsyZEPvwoBvsicnBoQhX6bPYtJIhGjMhOwSXM4zyTUGKb+1YOmDDbGlBHqqqe1
QljyyfFIkLVh1xo2iLnQ1GoazByFjEcyq8iwEYUxZLFD1kwupz0WejSL4LHWQ5x6STbX8MA09fTb
VY5wetjdn56lfsWKFlT5eWrKwlTf+i1L23AOMwexBguqsHU2QcTT/CubnbzcoL0vfX29etvSAHY6
Z+tVy9MZ9Gj6RxN5oklNf/g76KafV/Ucvn5Duefp16ig8YQV/2z3LbLPpF+LXsb3d/BcWaWn41C2
h8d2GCQTqxRv3AvApsbLYuy8juP9HhSBSgC1ApUTj7TfKlK9t2WMUd1ctVLtrLzLnt/pQC/956vd
jLS+1elvnSpn1llYOmOrjGFIwY7AeSX5nxumBjJfASbG67+hiGe7v/xxyqnwEFclJZ5A8jefi82Z
7pbWrG+iiXrA6TiVBAiRe3RgJD/aA4U+mjLFpsYmaKAegSbQi3jRMJvstyGA24ORGGzEyNolHDs+
TSFWsy3YlqxYVfAr8yMDQW0a7mhvooLvVAs64bPi3JZBAw8RpSXpbwZ7rA/JbUZ3VmRE0ezcIesc
ebty1eLoOPhOhDLENSK/8w/AJT++zKjEykiKcpXO3LJREHuPZ9lnhjEex/HI5NfyACg1XvZuSy6N
0UGr9YdN7hprtodAVTv7M08KiMEzDasVUhY9Z1vizhFflPOaN2XLjUYNE5oPAZ62tnARRHc6St0O
AOZ847fgT5vMLH892zeTDW8x96zy4BelhvfWNyLCBfDlwUntNoeHmCVC8yWS2eP3Eoo3YeUj/2pD
hWoqp85ZxSu1SJo7hd9Dxx5xU3TjQA2+MvnjQ3/p+cB2RkXBFDuljR1TRtHI/TwGfJLEI3AYibDk
oRIw+Fd8oe1XXE8cAKl3czsLjSqqvYGEWz3vOHj0RQsYUxp/gqkkD6P3dg1pGjXEu4hdYT+9ISyC
G/pkVMfrDVvpUD2rMQwtXwfWgueygObeVA19sBab6KAN0qI+lax4TgSm0SqJcNEGASzZbMkXlEZX
u98N2MHJYtnqR0WtbkUhGaQPaT49NQ7v4ZuaplRZVviNeCt++pwAx4FbGE8NNcU8ENGdJuwDVs+r
K/85jO4nQJtyAU99DrrnM36S8+wDucaA19vvJZv8CKS+HWuhm1BxfMTtI4n36tQfekpdb1B9MsZl
LS3cZJEyj735dYm2wILZuLo0XVSc4Ow2KCmLtoybnKlp2XXjD1pEDlybvWB0DJUvne1cQC1Zo0qR
obPh0wT0d8rT1Xyg2Q6PZvGC4CZi2ROmLen7Rnfv+Xb8tVjSBP7tGtGe58uzaUmsqNXsjme0HSTL
8qlgafohxFZ42X+AYy0t+L83+gc8tSRNxTSU8bpifwv6NrTsQtPMSiAtnHR8qiekJY3CMJpxCjMq
mUL1dADLeO8k/7IxSr/Gl3/lOH2O+7L3KMZKb03+EbkA61nTWC5EK+S/HcaKWt7Ic8O6F8+feVef
XcJsWUXC8B9eNh0LPcSm9KVkNVeKAu8iTu92McJuDnlrNVHoN8Pp3fg1t3/pCJ4AjpMJmKIM//iu
o379bXoRv30nw/sFkGoGfEm7yRAiUILYX00dWXpYZAlufrOdapn9eqDvDb6uUnOYrj0rwbGUKPtS
RNrQwstW9Y1yUrSp9lUwfTmv8e8UzXkhFTlGFI+YM1xwzWutq6refzz6kCHpgupnb7BmTbvYPGqG
B8P3KgEn75+Sz06wGfNfAppkqo+jGimsfR7VlL9ZcSVIyWgm0pRpSVKNrcChzCUwNhNCzYgK+ZbI
lpJMpw32HgfZ6LmM6gAuHTc4oNvESQiSTctWY+jkH+divSe7+nrXmGqTqjw6NasQkDzfxuVf4WZT
J4VqUtVihwExmv4qMRIJEVscyne+VNO9FYTKTTYw/naRC0l6OYB4jPn1OIW/vlQZ+Anq5XevPPAn
fyxe4/4bGEWD99BC1xl+ggNf0XdIrE12SCIXcR9MpcbvjH4VfcwSi+tC0gQLAend8ZW/Uos2gWFX
NKjUVqORJiLWkvyNroX5KNcUc4OUtfyLwst2Bg43w3I7gq7tZEJ6qQw0QRYL7uwqRv1xdXqHiSEb
qqn9a4D5GFouZqS/NLj1ghpuZyCwlobK67KsoPI9/WCEKE9tTXYHBHusgMWLLkod3986W3u6mRRg
ocPiwnjOsNdXs3Kyd5l3RZYw7A55evlhO8hXW+csKAiMROmTIyXRrdZBQmSoXuc3FPZoP87Exaws
uAuU2aXGF51Tykq+Hn5oo5mYjqpIySc34kKC6nAYfvgzdqRnwPbT3MjiiCXueHk4yOHPDiFPzJwB
FN9dyCFOm8r5sITELjBmf/nUcY2EiTM14x5jLv3+/LIw/DQTJFTaJbSAcvMiPCMX8l9ebNfDzLu5
9TO9esTnAzz+FF3apnhLtZdA9v560ZBsj/+k7gBmYSbZFNtQkK2tLABok9ErJbz4uLHwuJsthbYe
1ma6b92eH1xO+pEfZDcwL/qJLit8qwGY2a4KDq4Ce/9+w/TgNdQT0Nsdf9FM8oP+HIoEStoL2xdI
7KO3wR37ybY4DViMLQFBDGv0qnof2WD6EJ3nlDBroOY5sjx7S+03KIkwRIdDK4urJeOrtCjo+7w4
K78UwtoSi324/Sz1scsZPi4Xv7p3WY4kUfrFrr22NmZaK8xCt8lBsFQNmJalhxUV2rzMYHiMFA4S
GXhDrZlOEiff7iwj7b2ENJdWkJNgrUXCkd3cUcuol3ok792824tCIN+t90ikpNTmWbLSkvBiEXIP
hYY/sZ4UJS4lEKxTH2c04jXu2gbCKbzLpuIkE0pJkgCxYnmPzZI1/Zhx3vvq4Gcbl2UpIxXdADrI
GF17vJektx6vwRblzJ+mSlf/jLeEVBUcYPwbefjl2P5APenUZKxcXVhysBKYIgtFHXQJJxA0LuNz
knHqwV288ErIncX0rE0mee0NHVJkcoR6APvofbNhMVuFyeZQ7K15/cyyug8q7Ko3b5gPDplo2OON
rYYzCeFCtrGj/QCg4121wTc/WFPVNi1+iGKiYN+ECK+Jc7OIzrctEE/agRnylSv8/dopose5mj1W
xt8Q1UKWUQchgCD9Oybo4JotCiuFJcjMyIWnSWuj4Gr+pBKQKgrJ8QqSzqK+OGn07NksNWTW/MmW
/evHFp9mW5SRiePd5/6vzkKOlNI5bC/HaXSmzMZlFi/xOlEC7QeSyu3PaXlmU1gIEJUo573Tmjic
PTBJSJ4F+V0tKu8KHaQZNyYhmH4eIbOCzsb6AMppjeHY8tB95ZfhppRqkoGeMeqAEKB25xigV90c
vhJ6+FSj0WV/wFjASAblyBuUwUO3pOm2caqcdql74LWH9wxOndY4F2vWmh3HAZ+4+IhJyqy8lSND
mxhvO5OB0iq6J/VOB+mc3ao9lrcYu305Hii3G7BH2Uje/IVlhAYLfTRaXjSMSON8dXMQS3juMBYR
u+QoPhh24o9XL86iJbA5YAEOPhaoCutobF99Pha1Kc14tscCthBgRsGAMp930mEzfjIQMkPt2PI+
XNrlHuI39VR16iOU0QMSsPPWaGnwT/iHbCeQuU1nkyneX0rmY7096drHHxaTv1kd0NDirOR4bXqW
2uirwyIRXclZUaJffBOD7FraCgyrjPQh/e7XhejlpvnR+gtAijNHKfsM7kcEjpwzO4l5OJeE5OSo
6LW6URF2OsukTYQeuv2QgeUWr85Ih2hex1YSREGywOcFyDNExZhdYLeMq3aNes0ebqs+u5t83XbB
Coe1PnPKZ3I0KA+R8qaNH1yCrpYzR3ICz6BC2sydsMGfULuNKIttdUFdAfByi6vp5AxxeSqz4+K/
sXTbreRwxTJnsJBdHmhAGW7A+VrWBY9hs3DVFBa1f14WuaNOdE+cbCSYLG+kisrCqAaeF+9Qodkz
/EVCaPYE1GwCXHfyX3U7I/V7Cen4Z3w4UzJZRuG3Mw6WMxprFCSGsycPdoIUVFT4luG5r6CCHFpq
TlLYlmIeyZcsoG5z2DYmebrAQOlAZovyfr9aODo0dU12YRGpn9dTepQH/JJALl675kPpNLCUhkur
BcQ5Yhgo8KbEUxbWDo1U0zYq7GqhqA2WQBB1TfCeUXw9ymfwdz1DlB26f3E+JMzCwsiywuoLaE1k
GYMOJjtLJpShwnpSruaR4PZIL/VEE+yv4HxJ28WdcsqtfCl6cvN4oPN81Zj/i1V1wr1zwJWDrMOW
A1cgBTag1JbGqQsEvqJw/qJS5rNGcvGNvzb/J45uVSkXS5/N8Gsdg/XmT3RoqujX9Eg6AORTEdKN
yiWsjxGX0+09hiDFrKpVKfaVq9QMXM82xILDemqtVMs3kpJgXT/jUMSY9IXxgcbUkZ5EgKs7j1Ea
/VKWp6R6UkGtBdFqqEGqn19Qkn5jlnxlTIjeH7jWysLmkn5c4HSCtiN7cJP7YonQrVspVkiJSl6O
iwWzDVqIXj+pjKxaWUBlGMRAtEUpZ04uoUNVsfObVDvZADOF/E6oHaaXZFKB992u6YPkXs8NOuYw
bIuAqzW3wKzwDDRrX4Hvmo8gtUXsnr27t3fkQ5Z2F74zM61/oKTVSmjiTkxvcsNAWja+PyED6a/T
8Nt17zrcltdFBJ9hbzZXsqAXZXBZ9xKv1BjN7lZzoD7fq197thM+nl0DmIQfU16wAMvl4nZyuJ5Z
ZXL97Ft5fM+MnyZ0P1xkM2vxymBA1TCXaFEg84yZ5UADiQPtFSKT6migfb6jMuUEhgjLL07P4mKv
yClDgXthhJGs67a+pp+dhNPfsIGSoKcZYw89p+bq5xPgNK5iGkA/lOoXldh109djYEMpYr/xfkPc
jQNmAmY/ovHu+EvF9IPTxQPz+cFJTmRolL6EYslTxbSVtMsh44g/+PEmbdr8mRhqxFLxnSqRnW49
MTA7HSQd2vP16PKXhHE8ktBsORdCxFx8b8zO9HlORM4XR6Vnyygvkon+5L93G+gKattn+DaqIIjI
nqq6rMFuWryMcn3/DHfKjWKMRTUpSVVG86STqEnrlqcV+kVUZ5XYLuu1NHLQGrrXj6B40BIMtzIt
G32pSNuEnx87hzejNCRHIinYqivSIpordBsth9x8E2GnTBiNtHTvYR6lcxVMZIyTUxwUAJXIqgoR
1IfXs9TtjyvWxB0QggvZ0TUmetfDFYZKHylyJLlEWaadwxNRlHImK9Z0lE9Ow6TYX6ZEwPyuf0zg
4rjwkMMBTsNw1NwHsZuOyIIui9ENLMfEieCSwH54yqdmfEGnbEsyl8yHy4a+ZgTHyB7RPW5HjS85
1We+Lm2mej4hOXKE2ZRJI51rHCNNCv7fv7lS0G2pK/Ar/BdAzuB4K7N+rVerhadere4PGKtGSuSs
SPmIhTjCVkWGB9wo9Sw9uXYbcmcm4rjfRdTghQEBpPoqQkNcBo+Z5DDkM+nyrB/vxnNSBS0wRCyd
WWjJwd6QE+vbG5J/m0jXU0xvTUq5aJJj6PAzmfbMRP+ghx0ElbYRuopBIvs0JZZJ7ypXWJHRcR7U
UjIwzqzm4YZ1xFbYzzx9zCn9653595ur1zmgLZkBlsGUeoXKqtM5u+mpRp61fiJD6917YRGlUdD8
FILMn4EmA1pT6hcZiz3o1oVUf2Y8umJDogL7ePcuV7gQhWdlTyKdmWD1F73J5u2q7wFPZk05XA8P
7YsDaaY10JEyNgxNxzBiSPhCuzJytktiSy2yH6/j0cECMXdnry77gDuSyvQvmhY1z/TMstQoOlCe
E0UpUYGTTuE7p55jpPSQpeuw5J0gV9oX/N4uB/E0q+uHrpCOV2PbV2vrg7iGpz9/M66MfvUWsqZy
0gFQKhk9bWApxvetNxilP2/JXNxTSSIwn7mineWSPAIcV2MR2n0t1reMBNK5Vzav3oQddMISbCEY
xzrGf+3OTdORYPye0/H/sz0a1AgPP9IMNiL0k025fcK11yI1bMC9Hk74BN74Z2blPjZd9KoXtGBT
JI5z07tAsc22Cf8eK8amh/vT8R8e8D6/BjjrEGQ6xyDGnWFFSoRWPkQsGASYCHIbeAE6PWgbChjP
0jmcFtcCozQ7OXaPmSTJHBUH+oshBfUX6Q1vmO5PK2VgfnIWaDRdMHwymFfAkzIwQ0YQ0EoJHGfE
X34cp4Da8p/apMrWFMqG80NYGeAkrlkfvYEjMHaGGqBSr4AD2yPJSGG0/BkgLhnWzN3bCOzs67du
ib/ekcWMvrGT7Um8MZm8zd5BQJZB//5l9y9fNzu7U/g5zRq8K3tvYjvKiCnBtH2SFKBlgWuEjGVz
fJ9o5tOgpjmzaVI5jtL1zTX81Wxn+iREJGpjaFBMgLc0Uga9GanylcYUd4b2kuuRgiGaTW8aoVeY
PibfYrIhRLFnrhvEGr8dQ/RrcwnDWluAuwGUZkhZdJamGTS6+j0WZUGyqofY3wVnQ0wtQIEVz5B9
mikBNAqfI1N7reIq4Ah89X8LIvKGRMEH/QcSKUFxLmonYAC3jFzQnzfh9Bm8x+kGZNrQVlDxqrqW
06qEVCNiEghHNh2VMHYsqvfhcsDM3LzR31hHI5cSOIr2FoECTvI/Dw1tmOpuDHod9b1IWKB8n5UY
TzUu6+N2h9c8cj0SXsMX3aUFLaUBDpEr1mMewaMF+YxgFRhhqPQzxCA9VMOzuHIYdnFFjLO/pJwu
itZpHqVb+PF86Yad+eWmAz1Wdz6X/3jwz+4WuL/A3xg5bUf39+ecGW/wJOFRs4+rilHtIgTxFZjM
MgULl0C9GMCq3m0CKDUu83dMn+hqZMtPV1O0rUfTOKIRVi8d6s3x0FmsZmXau1d016lDTgG6zkNJ
1sDCNXnsuUpEzVD7dfv2G27/Y12ZmppYViCwFSZfwRxYqtqJ/cFNXSHZSmXFEhScEWy2HjBa03eK
CK7BlUBaukcEsiCAJv3GYBbZNVncHUBVhqGa2jir0Vbxa6uzwDJKpQkLMwHXEEQFgjzV1l3IeUDL
XB8r/HdHUsp6Fdh7Br5Tqltxl9HqqM3XNc2UxgTpDWMkHtFN5+vFW7nAfvT47G7LAWO/pH6n+HVU
XidDRMtBas7dSr13oi4q6FVAYOGRGjayNh5xVl/3ATC/mTtaNgYGuojJ+5/jWYg8xvW5isGGyXSL
uBcOHIirQCv3kbuv2KwgUzwCgAGz1DleFBURq8PqQJ+PMM5mIUWEONkELUs1rJ+Dlz52KP8GG6Me
n/KYCGK4svd0LSUfXO4dctgS/DQQo361V29fxqvoN2zOPb3xztetFNoLfJ4GbXO2tDJoi4KmyX13
7KCS4Bvh0yY7Puf3OZNJBOCP7EK1nNPRjBud4c4WrXxoWql21n9NTs4IKoeN7rfH1xpBXI0jIYkP
bhSi4j5dsg8XgbpF3DTf/MUNbJctAhl1G+/ESVyhgGV/qz42u7ldznEA8MUUFUMmW/O1fDNrOgYY
uZK8k5IGpcOlqvw/PDZRQaGiTbad9V1r/1pHOsq5TkTq50VXW8HSbWSox0nmx0sThKRsEZg9uF2d
3cRkWxOtvLF9iNgsfwJ+hXOdxSJFHSzTes7FG6Co1NUtdpuePN4sKjK9M3MUbwWAabJ9OYGi6yil
R7ClMxvopE0jOfJVDSYwyFkiZ9uBZtbEcBSzL88qb4BOoUII7DT8GvEsvR/ux3niKdwcGrCFB0n/
UT6UhtIseyTmKLoH7LBpB3BLU8uLOMb1jTx92B4tbYYvmUqPpj4RAR9U5m6PuxM4IxlMAw/Mvie7
+vv5oxN3IwEw+0PlOOAvvKktczQYpVdPyCTkGA+KsRlbfDUsYhWX5SwGxSBqWMS22c3aSyh3Gl1h
3a4Prl2fi+GCiAxMs49hgg5XCA+71c/JxW7DsurLNDxqPjhjGISApkuEWr3xSuoTHfRN0Y1w7SkD
z3dBOou1qJrdC9zoZY8pLQvEZ5x93gMmqdGuaQyDG9RtDm8AIrdHLEXbch8KI8fTG9P9loVbi9VD
0/0nzZRba/QefrEptdYhWPnqm4ekM+niGjWQxhJ/1c75WaPfojW80CHd1udnaqjTq9WAO3tRC/ty
AEBZ5x2N3iansaLr8LSLyFos0BtNq5hw9MNVjh36W3V7zXWKRwXIBCvrHi2mbnnoJEZDKx5FqA/P
/S/727Rn0j0W+a5C/a3oXFylOJOuy76EhMmnCYoMwFt8S52ZzDzwLaMR4Uhq/Rtws3QHyH612DzI
A9jgC/tWfCiRDjiFhOAYUIKNPiaIvJ0MK3Dp4wREvsqQHiFlJW7rhYi5y0jxPHkWGKWRd8hWTRLz
5UyfIzJoCRCkD0tE7ZS6xrRGTFPUuThthzj+dbFKVeOiN4uflDTdrvjdrB1AoQp/RXsU3dlElJUj
4xz+0x2A6fNFH0tGfWjNz9tZsJS1sJDr34wqjl0LT2zfGO5YPG3gqtjfcaoFzX4Ju2RULObjCCta
ixEzGHHe0BN3zzpj1ohvmc9jKiP2gqbPCmZ+i5LqPGIJ097RabgWtwf2YjS7VzagQnc+mQlw2rj2
GQCUzATf6/m4VAUwV8ICH/PQnMKz4uffF+xM9qR0N5tjmEdVwfoIZ4nQGKiFJKPbtU61zv8tk0aS
Z56lOyrIXCWY3WE8AW/OhoiEBomPfTGl0QxeTrfdfBL8d6+Jqg2E4zzrNH9uB5/mZXbPXZg3pX7k
5ddfrvDB2Zg/V07ko/jQzkZbvcUceR/i3f1pn+/QoN4g9rZ7NvYknzGxNhAa/5YQwf1mm+N/zwu1
Qac1giznGMcoepUoozFmtu4dE2GQNOP+IZ/tw0j3HzCr+DVl/TtBUufLLmG4/dDpcwpt3PWxMUit
6fRaRkksDIkpzlzlI9F6kGMxF6r/+3QX4A65Y9rOn+eEbPeIqkN5AeKGijRew1Gl34kClHDXBV6s
A3DA3l6tjexDpgZlEZ7fH5qyMfIfD+dySypLx4of3tpvpd8dp0P7VLO/XuU6FKhRRkp1HelonzVw
8bKqUOQHNo+THYW9skRN5hnSLqZF0HZm/c5N2taEpjulm1BMEft1sVcXKkAHmOe3zT2AVxt5VeWu
nqDb73jAgcIo6m0ZjfqpISgNRRawOnSJBxs1dLtdd/kOVCatduj77ZIAXM6r0tBkpohnokiNtsqe
PkaUNsXJ84agxshIbbOoaAcXXkxoDDxkgS7Q3dqmyU8hm4Jk2mUdfxRyW5kGSbS5rIEmeO+vNHMf
9wznUiZwB9iHcqmncmVYwd334FyXs2vTsDVS2vjojxct2X9qMIntdESzOuEp0R/3PW8A44mn7ZH5
rvVKGxBiVTxyt/nq4Z1mB8aM7vqzFD81QdzW9hw+Jk+NZ5FemqIs0CirfyNQd3G2dC6hpr9oF+rf
sHtvgS/rHrwIcMrUdet+gAxlPRJ3Gi13x7cnemklMNey0OTNAxSIQB3PjQDFtIxOQBiOajh2kTus
IxqtUdSuy8HKV9zagAP2/geF4pdcKeW2RmJAM/YbmH2LxmSiAjHNUTf96DZWU3+CYHsChA0dBYZK
Iunf0dTsxMKekikKVPvHBP/RFyCP1GBcuEhLWHF+XligS7rD1P3yKByhS1oB5FkxNpA1CO//xUe+
R7uSA/FgZDMR+soa9PXtJuPc9Brc6Fi4Va221884z+qacexie2Q7FvYd2OmlUe2/MQ1QjpcJxyNt
h3Uy6ecjKSbezPG9cQ1fljiM5kGa7PNkhZtUH2EEcPhIZ4h9WZcKL8TXrOEsCLqbhgCtj+0JuAMZ
WBOL1MFDyJPjq75XImHDi4ajmB01AUpz8KFmw+clMw9PaUxeOrl7p7oo09liH1qKqgD22j4h5ZWj
mbWBBl6hoUzEWF2nsoN8lzIaZWSh2jQQiMPMljGo0JX0qvPAFuBubbgvxBuE+5trMNBSNPn7VPZ7
Ep7CvlNSo0yqt3COi1qqfX1SA2BJDUIcz747MF6DBN5pyNh/K5jjS6yvFxi0g1xbo7SS277Hky9M
lqDF3yWY5ZaygXJjhhz9wTrKYYV69QBSanf8+1FmPDSp531s4R4+4LLwCOm56G3SFPkjevIzNkq9
PZ423teA2q/B+Dtp0VG0ACn5SotuU06Ivz1y13DjnVDOQyQmW2iLIC4qkNLEYEwkC8lJAOdYR6e5
HUdp6Cz38KXosG7G2UQDmrnhxoK134/E7+KHPmN1HKSKmXlo2xSi/0FHgPBcBrRooQ/WPX6IN8zQ
tizU5GP5Fz4jorXrWxNb+eLQ/JK67RqB6YPBXU6y9tlujYU1YQ5TL9WyJP1WhlmGGeCZdkyOYlhu
BfIi68PJornZp9QlVoA3Npta/v3H/EUtP9zsYpS+FHT+jRji9+hX9K1MKYRoEawehfzrT7Y58Ngu
WPT3QZT5O4Gu23Ps/qxyx7SpjaMo6omvzdkizxOM9Vuw0hu34qVzUdF3V5AG+zx8ECA4GnSg+eoK
RlSiSEzpnMY9QvDEo67S5C5XKbW5OiPfIwMlcJV2AX6w9zq1uzDxwOcVNWWLsiRtz+v5ptEYCzl6
Lqu7rjxEs1zy3ZHZOxcfZx1Y4Ua7wcCV/Ivw0RR72ishMhtjgFhmM0FV6FuV+vO2xvnzOjEkJp42
RUR+Xzz97N45dT5fOxdAno7s2FistPcj0UoVeVTfDT1NWlbO72WWth8D4uu2J3SET0cnQBSgk8RQ
Chz0g6EX9skd3QtKR/PHg6PvREb+3xcru8NdU4fuT+WWUdKu51V77jzarLAm/TxfiMakwSfCzlA9
VlJ2c/pRCoPU24W8w4S47FsgRBg0V9sAGcWYGbM4Lu88CRFM6jomYOALl1x5K5Krirqwt06po28o
OgB5kUf+z1/kjH+pTpGK1L9dYDpcWuvNTXtpWzmll8orhliPvpk6grTPcQpkJnIunc9aAREkuI5+
V+F9GSF7bhFh3zzH2b5m+XVi7yI2q5+VETBznZTNLPu8e/FkRzNQfWjyz1cMdG2nVHiTuTgBvh9R
1fQC1s+eOm5qvwo7qpWbPHI6Ja2G8Xk/O0wXK6QgCHDMz/d18toH2tkS+OtpYISUboLKLYDAtKbJ
kzpRgHBHnqZ1gUKh4JtUhm0Fp/gx4EVqFBOg/bWopuwvNSiAEtF6hMNmYy+21Nh5T+/Jeph1FPBK
UNE7NiGGk9ITlWHr+wG8aczBbEFK8E1VzqbqudVS0Of32sAvNo0sqv8zFzbp7DYIUN2yHj8JdwLR
hbRdljvfsjomtwvNLnaY7ar6YrJ61wd1wMThsbLb4vYWPMEpbJ75lEicmzum/IrbSrGzX9DZLXNg
x1vZmpeRtv/CQwpAxAEpiYedQxUC7vAfGdWi9UEVaMu51VH3s5zWwSAr/TaL1OUl2Hd2BWSbi9Hn
MWuwUxE9pNgXDXVmO2Qdwu0J3s2UR4frDEhwi1lcaZovP/P87wqZxlCLfcjZy7S4o0BiEBa5/t4G
qRhVto8oLVRU+P7Y6m9No4AmUmaxmuAuX5Odgoz17YdUDlewHmFmUB1wX/zBlJIy5wmXF6ZmIx7v
EgoA5G3Bj+ZQAwPtobBlHm7eLu5RuMOJdS+EViJxG5VBQi2KDAcbk2zwDLF6HnDHjQWs5fFTc6bE
81WInVkmRoryb3d5VyAUXm7CSVIsK1vui25IkIdzZE4UAgdPgtbc7VI/3snBEK7IkUiympYaqcNA
gPw3B+ab6mdUYQqFO+4lw9dUH9dw0utahld/jq0Q48hPvl6Bp4an5V/n6YBLhmEkh78MVGCm4usU
nYGazSlgr2gSiAPTYlk0P0luwcIu4K4hETDwXAGB64uBHO6hO5mmOD88ElDkAyoun77S2tBCmua5
YJJ0F6lZxrxKacLZ8/AXCB8jsQc+Id+N1CzGMe6Zx5Beesek+oMfdGqEkgwGmS75Ae1OxV0sczh6
EQFvmIi7AqAkLcWszzVyLBeznShaMSbMYagITKTECdoXTmpEwkkdNEgnfeAl8eXrcwmKnH/teVZv
8AbiQdZHtIBcmoD7qmwXYd9tfXXXlRPoe1tNVn7AmFsZtZLt6b2cO/NyhIr/C5NR5/hP6gSqD6NA
hmMQvamcKhAfjgSGJAEnFxaeSDqat2RalzD3CwTpfIHyyAUioSn+DBy5wart1kQkpQ6VZnK7hYgk
XLRaa9BJjBnWZ9uiHNtXy6D4rXqjdClIYD0eYdfMNLF1wsR3UBqGYzTsuFnteLJAWim/Mxav0n0g
2yJfcZZ7oJoy0r0vSzOvWhQJViekD+PIip4QCQwGjML6Bs9pyh5VumvCaoL7u7K2pG9SnFJCZuIf
FcsWNupbyZofeMjW2hXSvQfggMslAiYLYd8vyk1TnBarmpY+Eh9kDyx4gBl4RPfyRBWKsS9LxKBp
rf8TnNX9qAtBAqwkHtaAbjbXFhE2PTp/1B5MOU+0qFNh717YJZo3EIO51teQgJuq6B4y83qHQ4Mj
2QjW8xl+zl1nsqQyZJlAYdf8bWdwHJNtmEObDBY9g2U9rGcFou3GPxLvNBYfwAkkpq4518W8rMys
9dk3F4r3aWzpeKM/Amxdqk2Rvqkyku1cMMaXh0v5ATH/zXk5v1+H3widr+unQTqHdP10d8jUpI33
X8U+nAWTnvh5n1YM6/clqm7l0uka2ICZvn/YlUBAmNXSMk59cb9rwwna1qBgTEWDhziHhWWih+Md
dQxbnXc9O/Pl51iFTWQU4FqBKcph60JMTKVNndI3irA8YGRbwQJ+9olqJxc9qLvUWzBTwGQBdhwF
EdgjcaMdZCHodqQ4jYjG46d8DxzZ6Yc4uxsMl9gqFB38BGZSZ5ta5b3R7Yb4nGf/3miJ/C91mflS
+6eL91bVcmVLxKPi95i2nCcSO2qPm5AEnLjigLS6vqf+Z5J1HacwTwdIlCApqgOHclmOimdwIMYW
76Pr3MAiysSQ1QyN4Oiq0RkH7eyfGtzTJM5qG91Ys9IDkWStsNOZu0/KXLrWsY5/owUxp0LN0p7L
IDSbjxQdhfnjXWyZ4Lwu7QfZiaIJhbuZrb97ox6cy7P5XmYQYqnsLOrDQ5rcuu/btFMDy065r4r7
0KQ+BkJkMogBktdwK7HPuPOdakB3m8XZL8+/3pmrRX2XfhOY/ncL7NrUHNKy7f1lirmv4PKLt6jH
Cm8m5vHrwAh/uA+8/snKHiVXPUGeKl6d8PnFn5StnrniBIAwgdZ3S2pPkZMSvm/W5cvWB5HVB/lW
5u9t8ZSXkXHHF7Gf2GeJLLwPxOwOdzj0Lx85HI3J5G1Vfs7eMVE2HMdktIo7EROhAZW7w85qbjwr
AKUvf7a3Zpte/6gTEruZvNMAD8sfHq8EBtqLC5/u8Qy6Fu4cdlDLkDA8W/p56ugpRsfQk9xzT1fm
uoDBYBPjNTZoTIWlCaO5MX3K7R0YrablhxWtT2PsBZAy+DMmfyoiF22vJOM30ScrBw5lXosC+M/O
mMXvKGEmkHruWeCDZ7Qv2c0NGpdzSlQarxjj5bkCkh/xNPlXYlP5EEfXbYOsuXjmzLxvvPUIPtWh
vhgWVSDgAltXs/E4oDVPjYIHJ3dFWovMISbpzZuaKvskoiroFsORApBlMzv8FiIZ0D43nja43+F+
Y3DpIf3Ewx40+3fmw9+SlYa/+D24oJA5nYEBJDszJ9aiF3enw8LmK8CGWBDjc4YXrObwk6ApZ8kC
dkeg1Qvk03pv/pAToyQgaJ5/juUsTypJLrGgd+yGEMUnhatM25iUtw+ojRur8jXoDIDQPpwUzVxU
U7Ma8f4hE87r/EnBybd1GdMXS0DkmyGXzGoxKWyHN/sVFY+R2OhSG1mt4cBNzk+Cy5GVXPM2XBZF
/ueAvZpYMl/POHhvYI5NcpwlVXOP3wgudxxMMGa009Sd6vIswXsXQo3DuF/nesEqJr9PTPEALB6O
erhgd60NH+KffewRr6P50ekBxYcb0BbU7RhZXM8Y3pOWoSgWljnQY9sZ3+QSp5Jo40ArFJpNPRSi
uPPu9S86uGAh+kGjTqLAEG8u1Z+LyX7in2BJdldJyF41WdGmAZs8rkglatyKA5lhtgeTWj3A8kA6
8nD4pvU7s9YlQX/qjMm2EX7W2uc/GoBmcROyU4Z6vF5CNk5kGKUSQG11MhqHI27ErrNmofG9nkel
48FnM2+rKQlsFAmE9UXTJr/w5QYUwALFQF8+hLwRaxHJeh7kUrp0D7ipmd4NotsUej/rcgP/iq7R
h7v5UyU5cNpwQ4jlAggqBf3LrGLdkbBFsKMfDAPRAUOoRdtD4rQUtTiBafMdvQLz05SwkgrfrMu8
GE+ptd4oL4J4FUMM4SZ/OZAAhaqufKQe1vqvlW7yQl+gps7oNnrqfbLSv13L9k6vy13d2neZX+We
jtBYcYr9eD1fkSF9xvpAwRHXO5kJQd5ecZsBZvEwoKm3OPXROXAj6c3gwGx3wIAEjYIhggTeby+t
cENDLMQiqbgfbQBNu7NEwT1EXJG0p603yDojuXVKGRbchPYzSKd1KaoH0JoVUG2dkkzZ5Fbiavk4
lpwAvnYfGP9BK9rm/Lui51pNFcqSna0xrnxuNBJAvcQqTYHh5Jyl2jhtgyiQHamF4W8zl17dt93P
wucGO+Qd1y9rHFeuX7nZQtu6RSs0tIz2vaXpNRCZ5MDXCZhZSxApvXR+VydV4zux986XJb+HcOUe
6CCX1EF8bxCi/TDaEecQ0UCLXw5LlchK/IM5a7+MCwCUrY0rJdB2j3b/xGl9ga6iskoo4YiySBiM
VRSKmx7Ou6AaZnGo/oXAScVZHygJjiMSxr/NWoQ9qAJEIfiY7tjwBNobwlqpE+yp1gVjzRYCAztT
Uu2SIso3MWCC8HxQwLla1CpE1DI1ETlbPefHCm/opdILY0FvkrcXTMGZnajVxP20hElyY8iausJ8
gTtVd4s8zH7Tk7J4u+12xG3juaehXKxY46bCcXuF+WAUtHkS3Px8GA29QwTHyXuZHRYFbE1u9TJ5
msWNahOk6woXF9y0DvqEoeV6wnOkskpzVqJB9O5Rf7fGnLJaTpQSeeV49PdCen32wsM+BMJVzLD9
5b5TSIblxwE+VR2qRrgsbLZjZbN7xco+3v4v/r0WZ0amcEHqKehnIZaPy6i+w6Z/h+58v8iW1r4U
xyn96CxTpDlLpfWSO/gEc7p8o9lJ2Q00ePajNuvMdsQ0PT1DZU313+CJxTfrl4NuQc3neBMvYkSW
F/C6+t3ln4Lnva4DuE1bC3M7gOOg46PlqoDbNNGr0866jGbrV+qCBagByzF5dpULWuGD+ZY/8lW9
ips4PSrLXj1I/ZprJe4PtB9j8E87YAyb1+XU/XBGAurTywTdCWLN5yWKgMUI9mNdtJkHh/QF6Rdq
BYWYM8npx5rOMuWRlv9psrbKmkjchskDyV3irdZ8JohBySOyNRc7m0OWQ4Drhebg4exJabkIQ3wy
69LAtdjwUU4W6vo91Lw4IV9oUzh2vgI5Wc0iKRluPrnrliOxESMhrOwbHy5G+oklvXlklGoxv3Vv
NLFX2OnEHUBaSBJFHBo1gD0GV69DNMo6+pCTVcyQ4ts0jjEKNvtPP+09aXs4CMUW0+5wsrbIeS2t
/YW+WBO4krHaEup2uebgrIsVPVj+fprwTJbfySRhGOLqXejct5W2b3fdQNx+sN1jpnbSSxzlDOIU
2KKmJvc3iYmh+gnoIazeSb1LekXnar6sVng+fVzjQOyLGaMfgmgDuN38hFfvwRl+xri6BYMupgbj
07BzOA9ENoqO0ZDrPEcVzL5sdfQ+CRAzgQIsBVvSSpN4MVH5w/+DONdNUH1sR45TbBTavzzRMC/q
sVMVBhVCZbSdsQHNKHQeFTb5dGu5T8l9cWSqlROfyecUDYgaK30Fjxzy3RKXs/txJfXUp7HOiqjS
pqNvLzNf+9LmGgAXZqpe/N9av6mjytqhVHhRx903VF0cC/aRyINnN+Q/2FIWygCsX1RzNddez6OX
VGYcCcof+1FR+/IksKlHXhRYoueVKVCKw3uiJSqM76lhTe69v+0BWnHZPQ1/XYc4y9UXU0Pg8YRg
fxz0FYCGv7e2iPFyQSQMkTfWJBXa5HeoeQos06lwuvpHIboKc3aiy1Xj+PriaG8AWpe7/8sPRXsn
Epp+L5btCrcZshNCPqucyitja2inMLs8gdWBweHNeSmPwkuDT7r9uOkiy+cGUa/GmCfM64+Y+aor
wPREzHU87N88/mt0V3roAPC0be6IOcx/6MVKLCZx3c6DlH2a/8ifmQ9hgpH+sCMeYPonhVu9H4Z3
BNoBb9notGfFMHiQrSfcIN/6bWXUhG13OuutBn8ZnYzRcxiz8F7XMBGpYFfraZDZZr8Jx8SUV3FZ
emlMzsJyWV0r9bzS9tR8YPxlTmjvHBNKsteNrpeG8D5OzJ0ZbYFWJg0CexNELGCfIAlWPaBt6bjo
4tfE4w5EoPqlBFy/xUSqmBz77JuYKN2Xhr0njPGrD6l5NALUe8RHOHzyaCNzWwu8UufnRMPllNlz
sPR/1MxKFJn0tH822F6qnFguHIxMPkdxkz5/oUQ3eDkq7isZ4zjmXTibUbJZNxMSen4KIKOgi7Fd
cAPD8X0+5Vo9wwfGCpYMTT4WOjKpD9oML41bH2Ad+HJYQMjnXYNHVCg82KK3EjHMuqpH/o+iu7GB
/FLQOkgUfHUUorlPPdTJzmqMhQCSsld7b8K4NQ0Xz38jTtlicuy8vNCHlV23HV8Cxv4jSNQZy+wV
laNHxDCYYDafR//y3pmstlUL7NLzyIKntgwxmm8VA3QJezS4ly1u6sI7TGOz2443x4GeOW1PhbMQ
Qt7KjjDVaWQjFcLInsphJOv9+BrHCDGMro1yKl2TcopPb/amU3sxHHrXJc6GGU4yEEx+3anrQ+dE
GBR8WpY+iE6xyxKuKoPijtUzjYOv42uAQTpQZ+Zt5MlUjDOZR6LjEOIceNRNPn4KzGRPOzafXZR6
BE4tM5sZ5qfUX416VYNRjES92L7fuazfMuMkiEeK3oqXKpvjY02XiH8p/MnOKCNSfEq8MEj6vFXE
W2rvWex5hIglYvpRR9Q1hgHIcwPurh/x9j12dUuiI8r0WCmawysc+GX53a8O9G12x63kQb1dD5K3
co4eqrX6YnFkxwjpcpTmSnof83JY90NkRJImjEHJVDYNj2n2qPnE5dIDmNIcK+p4YZAPZmoSHZGh
Me+gUyKsME8HrOr5hF5VX4jCcG2+fUfaahB3JhgYttpM97ZvGqi3V8fxBq6kdZmC4czJspyLAnUS
Yfkap4QG0UuEyr1j2ZGgzKBDb3NocDRmQ7amA/WzIS7toqu0Sap3NCfAlxj7j2dYkKiJySOifiyu
kceNqArk7r9r6KesrPPcaMUNpohVFpus2k1rswKWhe0tfqL7grqCLF/Al13bqF7CV3il+CmPAW+g
rEYin22L8TQ6VUu6fhUJLO7ekQ774BDRMO8SXv2WwGJag4gZR64I1I2xbWUl4UxTP6rMGQoH5Rcx
PgoBfpmqum9gomt4UKw/8XEkXZObECFxVCGdUF0gx5cht7xvTxki69ZtDEhMmsz+HPZXcSKstjgr
W4y+WXl1JCmu3Ff3Wvgv81v3HgSRhJ2bVwVSbKpkaJkx1AJ1HYr63K44Z6B4T9NsZ8Ug6Cc0p2Gw
9wIACCJJ79AIDXAiUQJm+0xS77fHFd+dJ3IcTeAiNYF/q+i3tCl3hEnOguTc951F0Lfv5cSJBdfi
C5z6J8DW+ch4LN1nX0upLdgMF6/om5zdRzSvXfasu7olec5raFJNRVTN+PPhcFFLi6D8JAwEq1h5
jzcdnyMvGCDEsWVQYDmRKmqzVZ0Cay0swLOf7oyybdahr9GBUwso4yWiRDJdl/oZy7DH6aBQKeVm
Pbf+up2iwFNG6SrRdZw8v2x0X4iwM9FH8tkKJujDxqjvZXTST+3Oo28jyYkesKVf8OoiRHjzTY/w
hYfxmTrCjC7g7z7kzhtvN4jsWr1EZ3Yhz4XwhtCgAH+5wyDFScFxgvTeyJyj8adcOWShv4VOjoqc
P3q6+M8OCtc1M1T7NkgSQy6hUbVkiSalye0+dv3AjM0FJGvgn5T3aB7PcJlOJGfrVocmz/ZC9eTd
vw/7P5ZuhAiLoOxCYYYUJ0ofWe8FE3ROpoMTa6vhW3mprWKSDENGBheGPVZxRnU31mdIL2XwwOvt
X1BVFAh681Yb9eKOCeW3MG9VQ1Kv7IqEDyj6myCuCpBXmUqCQSvDt2D0uWeRxlVI3hvnyAJebS1m
vIWVJbmxhQ1JWLD6+NpWKC2q+1Npq1+AMC5NgZ3MxzDKuykkNa5yS2Z6bxeAuKPgLXF20bUEIHgt
RKqTKpViAdHX2RbTaisXULYGaitajqMX4FjHIeZMdfo8aYwUqCR874jwkE1O2cI+f+EwLnwo+83l
f+c/0PSzn24UnSHGocGyVczugwDZNkfCZUw94TsjZOoeDbu8VYVXYkQm8qYieuGhpMlq+0xAi39/
QQislhFOnwuA5yxa/8vhwd8ZVsU38teA9Kqrbc/AS4ER0FzIXGC5X4lsUiYmYs7TIuMOxtedXS6m
1BwOaj7IWvDKduuprxzJpKMPOx8GQxT8M411U2QRplbJ3ETSAmE5Yn2MhLJfTN3ge/ISUVlQSTJJ
tWUedjmgH9i7vqCMmbH6sd7KzQ6+0VIsw3Ks9DIxYewbmly7yBpugMlTkz6WuldoxYuP1gUrKU2J
09LxNaWmnrbRc2kNfYq1Oh+Yc38ODjfEz0q4LNOr3PH7pKP5FfN0cUImsQZyb/aRKUfG2Oe+j24y
O9Y+EXq7fCpuO+JDZADHHGWarYb7WFnUQ87oEHlr5g2rpebymc43IDgsVKV54xNH9SrqHU6cPNmb
nZwg30e7GvqGszdH2emTlHRVH3+x2RaLUpqY2yJN0FiQYhXatio9DYUMUGgrTY60lybqki0MQgUv
zorivzOcUJvVn3IZghmJm+y+dHi0hSWrRjYDAhQcFRTXR4bzoiDOLNfIsOdujncQYI7bJ/2ucvK9
ZAozI2v4xA/PX3otlM0mH20On7uWufIxt7m/Izis62iuJzzlQcvUfv43uMx1nVKPw38Cgx4Dec/A
XT2SmW78Sg2MkF6xqzm7VwGjunBGZDytN5WW8IfaI9p7V8+7s8SUZVqF29wUURSdrf2VyvRi4uLS
Cm0jOWWD3gO3tb6cT+FLlId6rQ0NVXDpACGGg9kD4uJcV8DDC9cifjRPQQw/LSbBjwjZCQacPL14
gkTkJ4XoWwbBZvhzGAIq2b+YZAsFZ7IlcYuvle//0hQi4lJGtiXJZn4ElpGMU/5WEczqNMiXwCTU
1we9YKfAfQugFt9QTzto14P1BQCQK2t7WyMVItdLQKPqsFEEI+v0wOPtz/5/JuLKDvqoYzEofIrk
8iu12ydiedNkc2KDXDWrUwN3e2AwWokiTvVII6AMoxEcDFSKQR3pmDPEX/p4SgLgaLDxpvWDC+Uv
/qSeueODTAi50ZPpcU2rNM5IkXyHG/9UJnu8ARGhP6qcvjEuyFGwzsgw/Ha1P+qQNziKqL0x3qq6
XZtGLxGsIqe51N1/tSHmJrGli7xHvXDWgVmpjA0UBqLqqcfiB3m/SjBnwCy4T5gHIuCnvrLUWn9a
QiWiAGcU9d7ymgnhPgyBTv71/Oic6nGxoqtuFhdZbJHXHhyG8N2B0FSOJF5dV3xAjywl/pxKaqUb
1EqJsU4MdVXpz1/Xk4fiQ3vIkqMqzY5/AS7Lep84LQAzd4UrYDkMpLmwr/PGzB0wGkIb2aBYbXrA
kMEKtFxtdiVw1YAGotUXC16e5U1rKe+akNigjFBTUZj4LRP+Gv5LS/QteNdDEnxf/WU3ugONIH7S
5tnBwIwEPhCmpDCItL5AinPDNOCSEiXxJe8ZPTTmSpJbHCmdqaoNU4Bf5P12u/YZUX/HGmU24jdK
49kPc8bU8bqpgai7BRGifBra95xk3cI/+1STChcDdm8lJ6Ghs7y4AOrV4LQ/EvrvPTWQiSmnCfiF
iq+XPRYhttQOzuo4jyvgTL7EIOnAKMbBvn1tIRwsWnIK/ArKOnrDZMi9jWcHs3EOf1egzMuX8wKI
ID8AjLfttJyCM2qDrUsRiQaS5ddbeDoFfYdDKNncxxtAi2hjTI/9ZnrBCHSSmIA7hsdTjs4fMcAx
WQXFVAXV7HekmXSuGKU6WHUmfBpui5uq7rCsusijaveQ3r3favMcbpD7UpnvNgE+IUlNS4hebeW9
rHB7vZbK2O8FCTnB3eN+r6Ti035r90b7y2bF5K8q/vkaEUT3lqZnN52AQEsaPg/uER7RzkOtuAwL
hofpoi0Gwb0ip23xMEgQ/3hBl5KInr4ODpu3NLZUxJEEC4W9ptB0bAae4blXMAqt19Zx9II3TFW/
OSaKybWWnaFgBo00zj8n0Sa++JLGlrFnf7VBf08B0MvUXrtHHye3tGIz/oZWcvYuTwjbuZ4yyesz
JPANDOdkh2kUyXe+DQWyTI4zOb7Lb/Jpx80bAUztjdfd2AgD19Skf07DxVWdzXdYjgWor0Tj//pn
44pN0kWLBMAtB8CYo8njuhTNsId/Gc03BeSYZse77DEH0UqWHMa7gipUTgPvisleSKa0zxlZ/jFV
5BH6okzZ6Tva/Os5Ik9L8rmOuKzyl6mK21/32DSeJJVZdJPpDUb7tvH1WBC0u2XHYRhIJ3IJkx5B
DPZ0KWFQ8b0Ovl86XGZUaRVBnqFK2DJRn3mYSXAp6c7H5bLSljjHM5IQWI2vxV86oqm/4iV3Npr0
NHslN8O9tdFQmLDUoSXmn++wtczKwsfSZLISRdh6itI2E2ZGZ2XDnSASuqIVZ7FMeP5MszVEILcs
U1PkfhyIhO3KdJXJAv4hi546ICzMf1yxn5CFdmAxGZ5YmbZdsKYk7J1uOiYdYsTdpJNRMG3xP7w8
wczoZLvRlC8kcGdApMDmPoNzwbajBeCEndtTClYnwtGfR0CGH2HcwaJGTisc+R4vWS9yPY63QVmd
LsOp2VDcxM4TNP7IRwY+SR8Chtk/FyBf+YQuNrxjbceLcEDEFFKxPA8wtu2e4iXn26GFo09tWU30
eeiv7pzibtdrRMfYBwEE+wiUl+ywd8P+lzHIyBhn5mXZ4eeW/5nnG+UYlcGpifyr/r1MrqhJ1WXq
s7+A2mpwRl4fOEF1mQQfVCoFz1SWabefruVK0b4NvFZ54bpdo8k08VJoX9betUX9MfHu+/fnaIdg
uj4+4foehsEa9ajCmR9YjHk558fYhROnv0Dh6FSRivPFDHKMW/i4NvjqgGI73Fs1+WAnEOwhJxfb
gKTvjreQROAptGqx+OaZfnS71vU+8dPmkrD+fWGgRRI0jPkN4GQXWnBhuNlmz7jfIiqaPAcQXhQO
MfKpgu0T85VV8MpO5LGDT77oF1zH78e5KGudD0ZIyIU+8giyYyoKBvkPbskaqPoBnZgGwQcbi9mL
PLh1w9pS1GC1a9jiVBRJqfvRJK0tTbujT66quRUfuvyWfbih52cYj65zfN3+xxvYS2vtSdDhqHAm
MsHm+3DVTvdEMPTtbiE9ajbeRkRg1buCQrldiVMpybHNcFZSR0DPBUgbYLHXt8AVUAJFWbtFP52q
96mPoPDtwrfiv/d9/SiEfDz6LXUd0sKfmGca/ySTUN+WHHRmk5Nc1upmpqzkMc4yF19dD1ZCFud8
fnxaR512IDFDf+qkdyngSbThlIFDtJVcd74AnSmkfd3kRhynddYD/BvcttxtzTBZYDygCcFAN3YF
4xHgjB5LhQv7WSWv9czuJRzpXhjQieXBbAXt2ftFY2vjGrsBQrwgLQ0aA54VrvAdQNn3ruPPLFWT
jtEUZIZ6G4pBaIXN6DEIcfB7aH8fMckRcG1hEFoDaJ/YBkHrTRLj4+Niy91MqitADhi+J2Hmnrak
jfgECH19ugiSXEC52201v5qEUnH3YWvL/BnNcQV23Sssu5ns3op9uRKghcT+9QM90ph2NvGnQZ7l
p1Pk4HmdBixeXub6SE+WE5mwwoQZaCKvHaoyjXq/3AGtfWHmZHfTrEF1xb5Xl4O2PXqSLbsrT9vb
E3jf5rJtC/Vkmm6FCGL5sLniu/HWAWhcCvdJ2rVJjok70pXluMezcuM3NAmAuoza+fUNeNsR+Mg9
yVWWazGEqFOm5pIR1G/V9ACCooWKoAm0S/olBbio3CaKQkjU6vnx2vOnUDqQfdg7XXtVEB3vGNIA
dnpMGvxCJdpnxha2u7GGngFKooTEaJpgr6LGl3YmW5jpL3kWhjAY99X2mwgJ8HI3hmUOrNwlo2Y0
1PQakOxZGo+CPNEifbLqXkH7rVlr1ccsBWQh3Xjwgxmq7Ihu7CLe8i7omprDGwNFSQZPD2soQQSL
jVM8TxPKlwzwOuDbOoBVCb517IogtfJo9IK7vVFZl9oK4X8MHxHnYAcumyW5Emgp1mRhkCLgidkd
obJ5sqgBo987ckwKrbU+XKO9GLboSgv8Pg3CDCXF+mhbSxvsw3MK1NEXLCSXcgjGr/YR266k36YK
j5S10RRzv3Pb5jUCsmFdR6gU3SfRco9n8aGu1RGsGTjkZ1oDM2LtZNM7TJ+QGWQzvyoeVDim+mhj
fy6lp+tJS7PcitNpdgvuqrrMfIYPKou0qO1zoykVLGQx5DKht62idrxVd1co1i2AYxpC4XUYYTzj
Dh0C2rBccRzHSWZ4wqYpFcKbJHsQN/iwvAZuwzz9smsS+nGjpI6ZSoaIH6nH+1NMMTVmfdQXdEl2
F7jBNoVR9apnpwK5Gmoqz3wHGnZGFtkvriVWLP93kpMJBSZJRd2RlNY7t3WyDHK/Yu3CYR9qZdpi
NdNgsFSrl6CbOrUmeEDdClOP9vJgSZiQOFK2tpTORB1k7aNYaKXZ4I9KnKF7o4a4mr1s3mRdXIex
h/irrSGVcmUxwVO6QOgaaiXDjCcOvMUHe1639sb3Tm1Mp/Z6uj4H7HSVHyA77r5QcrJIa+fnO793
jXq4Lm6g5CuMkqaVY8sIyGJRCY3akHxeHXdRnO6dxh3NQsenDNlvG1CkiUBavqrzXHrg1OQjD89Q
wVauumq9GnjqoOPTJZALKSSKau+ehW1m9yHF19W94qvlS8WKEhEF+zpMOnLVRXHJ72ixmRIDxR/N
P3qu2vWNrNub8EV1hlWi7qfTP9ly0DfWNJA9aR5/mhUTKKUiLRFSEUBiwkFdKakbHcAfjhTQpnmE
mUYPf9xQCpwAi7qtOahvlutarAEGdI0Jvk6YxekE+G9A9OeBTOweoAE5UeYqJ+9xwopXXLQB88CN
WAE3Zq5CsMdRxbm4pYY11OIhj+T2W/AOKjoQ34JLtqYNQV8O/8v3SDeZrkoe4AgMKxGqgI2SnR62
VgfrzrWI04GRm+L1yK57n0VZndGpZMuSYYmc0ssYLBtBfAA71EOjhj1KUdgMiEWgFb5TB3dL37JR
fNC9VK0efCkIoqbAIsQpO++R0mY2rHWK5HI7zFGVLPIByuhUdsDTJtIabIxj0+wL1usFpCyFQU9J
WiZoYox9P6cEy2pHVFREheWGGZsJDIUE/1qqQqBfQYXnBpYNYrtPiQWiUu3zZNNCYgsVSzOVyOhU
1ac+MzkbD1x75rDgQKIzlbahBAeHzINFtTpVS44qiLtj53eY2+pgICbr2t90lD4fsytcWeoZyqk0
za0rIXwcWGwXwVTTesK4U75igjwOr2zxhvyJpKdadsMefA15QOvqU/HbqlCXfvNsWe8n8zKqabpJ
M7b1TZig18OI32qUUl+f3Hv+bAqHfHII2CskC9iIraUknJSO9iV2UBz6fTAFW4Kg8ieKcJXdoHbv
0qLRM6zM6LagSYUWmqfybFTQD9gMPbazCOWByksKvZikZFlTImsAKccAWyir9C9LkARWpnPkt2Qq
U8oJj+QcGiAXyxSZIPFRTY6jXvAE8mHCGOi1t0apoVCjJdn3ZcmDumcYza4Hg+zbInosBv7Y0XaJ
gOUY5r17mOq5YlYixTashRxvTfDZKRWlUjytG3uBCWnRclm4V1twjdmLs6gPqDlkJPzLQZ35eZrV
fIyhc67753BjStkp0M8WYNXP0lmZu9hYDlgi+I3CsTEi/81fDJV0P9A+pOJ8WFJ/gXV9ZHN0oLXx
yRxjus+mldCqeKFTyUOOkGuxaciRh6r/HP3ib9veJdztNzuB3fao+QuJ9IuPmU0yX6H1Tmbv27IL
tLSzCVw3vSbWUOeMcWnjIV2K4exW3Wpuypc/hKwnx2vylMusmOLpySElWlF0N1KnqdtBZWsUdo6F
jeGs86Nm7lddkERL06krFddcg4Cu1eDy/M6mPQNFSGv0R4jPwmYRrZ9c2CHy8Gwf1obOgVfKYEah
xBCI471g7eERgRvCRQ+uq/f1cLaTJgD79cKHnV6rm6XpTAt6Th4ZWlCISEHNeH2cw9KJDo6b5Eq2
IOefXEaKKbemg66AuEeknKrlAjgsv3BJTa2axXIF24BDtlU+Oi63gURIdJU1mTWbXYgg5FaQEV7Q
fuPuBqqRWZ+k6mf9hDjNQgmZrl+TlB5BIkwjqkADeyUFGBZM2NnMzsSozrcY+rvabZQpiFcLIqHB
M7nWai+MUfSp6Eku0EkR4oMXdMs/6Z/vAcoWtJ0TOJGdPtSl4cpr2S+9OybqcxbbHm0jzKwNy+Tx
djl4JQ5NUrS6NgfxZSbLDs/KxcDLGzji6aLNFRVREVhLNUV+sJ0iyRRlNLmlrj2oYVSRvzj+FxyT
jrBsy+zddVyMXWxkbWssiYAuBO7dpDlNpowDECJGDgz/j5ZhKA1EpULhJhg8EiG77PYRWzOfp3FG
GsmrtVXdOvzyjaxyOM27rciFrVkA602A7l6RVqkdRjklA/8rho/kq95AQYZk4ECqDVCt4wVo+F/S
19BDdjZ2HH+Dt+nQxlp6uHX256H1I3RDokIaOoyBOY/fPqH7A1miz02XjyH2QIU3gUnmJ+Rg5zvv
neH5S6vZLkeKkSG1I1sXyZo3UgNQX+j21SQnYX4NEgwU/Z/ZcT/543IEmWTPwNi45Q0X3yry4lX9
bwNy8nh7JCI4Ed8xJTuadftiF2w8q34a6zAkNtWvaC7ATDq55D/5chnUPnAMEoKRNsw6r4y7btsL
FQHnRDB7/v1KtX9SD9B8luNAOoDitxt+vvcewV7kYKXkbtpRA+9oSrWtrOoq/erRyKDfbYZ8iYhR
Ks+zx3GrzH5DOHn2MySiK6hXtnSUsUKf83NiQ4AMCB/umZzzmL1klbqtcGgl91DdJ4lETwm8X+Qz
9LXRbc0Et8pvFodatXUIkb0gV0lwKTPwN2ih26QaYSOjr2vJR5TqEXlZVhhbbAYg1Nk1IkH8sQrR
EkFWxPUmNXny1/7kYmxmIR3weGb97f5wS2mssl2bg6bNgah8nfH8xvnsA/ADLzDClZIrZZAx/VW/
4WFTEinRRwiqCS2imP5aZLOCxmkXtZQfHsi1d3i2eCheF4y2azWs2MnLuCJXFxDSsgVKKrCNQJUj
Puanel57YKI/RtO3JcaGwyFZD3h0lsI3YqiYt2Wv2xrGMGus5vE8R1vbVDETwpBP9nPazJC04wTD
zbAFfNU/JcgTephdiZBz6+cKYatlOBpRIQONoay0IrYZcebpRsxA4JC40XPEvBfV7vOinvgnjWcc
M7odLkn7/aT/+KsnhiuarfD1I/O8O0mFd0cC9TG5qR8bf54U9NpORB2lwuX2XYz4fhJGNRzRqhPq
Ef5oJCi13tFutlAoVTXvvbfmK1Si90+F7IJLgoajtt5YeHUxa8qS/JDxvft26MUXnhxk+vfkvQ7E
Nw==
`protect end_protected
