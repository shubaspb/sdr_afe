     .update_0           (update_0),
     .capture_0          (capture_0),
     .reset_0            (reset_0),
     .runtest_0          (runtest_0),
     .tms_0              (tms_0),
     .tck_0              (tck_0),
     .tdi_0              (tdi_0),
     .sel_0              (sel_0),
     .shift_0            (shift_0),
     .drck_0             (drck_0),
     .tdo_0              (tdo_0),
     .bscanid_en_0       (bscanid_en_0),
     .update_1           (update_1),
     .capture_1          (capture_1),
     .reset_1            (reset_1),
     .runtest_1          (runtest_1),
     .tms_1              (tms_1),
     .tck_1              (tck_1),
     .tdi_1              (tdi_1),
     .sel_1              (sel_1),
     .shift_1            (shift_1),
     .drck_1             (drck_1),
     .tdo_1              (tdo_1),
     .bscanid_en_1       (bscanid_en_1),
     .update_2           (update_2),
     .capture_2          (capture_2),
     .reset_2            (reset_2),
     .runtest_2          (runtest_2),
     .tms_2              (tms_2),
     .tck_2              (tck_2),
     .tdi_2              (tdi_2),
     .sel_2              (sel_2),
     .shift_2            (shift_2),
     .drck_2             (drck_2),
     .tdo_2              (tdo_2),
     .bscanid_en_2       (bscanid_en_2),
     .update_3           (update_3),
     .capture_3          (capture_3),
     .reset_3            (reset_3),
     .runtest_3          (runtest_3),
     .tms_3              (tms_3),
     .tck_3              (tck_3),
     .tdi_3              (tdi_3),
     .sel_3              (sel_3),
     .shift_3            (shift_3),
     .drck_3             (drck_3),
     .tdo_3              (tdo_3),
     .bscanid_en_3       (bscanid_en_3),
     .update_4           (update_4),
     .capture_4          (capture_4),
     .reset_4            (reset_4),
     .runtest_4          (runtest_4),
     .tms_4              (tms_4),
     .tck_4              (tck_4),
     .tdi_4              (tdi_4),
     .sel_4              (sel_4),
     .shift_4            (shift_4),
     .drck_4             (drck_4),
     .tdo_4              (tdo_4),
     .bscanid_en_4       (bscanid_en_4),
     .update_5           (update_5),
     .capture_5          (capture_5),
     .reset_5            (reset_5),
     .runtest_5          (runtest_5),
     .tms_5              (tms_5),
     .tck_5              (tck_5),
     .tdi_5              (tdi_5),
     .sel_5              (sel_5),
     .shift_5            (shift_5),
     .drck_5             (drck_5),
     .tdo_5              (tdo_5),
     .bscanid_en_5       (bscanid_en_5),
     .update_6           (update_6),
     .capture_6          (capture_6),
     .reset_6            (reset_6),
     .runtest_6          (runtest_6),
     .tms_6              (tms_6),
     .tck_6              (tck_6),
     .tdi_6              (tdi_6),
     .sel_6              (sel_6),
     .shift_6            (shift_6),
     .drck_6             (drck_6),
     .tdo_6              (tdo_6),
     .bscanid_en_6       (bscanid_en_6),
     .update_7           (update_7),
     .capture_7          (capture_7),
     .reset_7            (reset_7),
     .runtest_7          (runtest_7),
     .tms_7              (tms_7),
     .tck_7              (tck_7),
     .tdi_7              (tdi_7),
     .sel_7              (sel_7),
     .shift_7            (shift_7),
     .drck_7             (drck_7),
     .tdo_7              (tdo_7),
     .bscanid_en_7       (bscanid_en_7),
     .update_8           (update_8),
     .capture_8          (capture_8),
     .reset_8            (reset_8),
     .runtest_8          (runtest_8),
     .tms_8              (tms_8),
     .tck_8              (tck_8),
     .tdi_8              (tdi_8),
     .sel_8              (sel_8),
     .shift_8            (shift_8),
     .drck_8             (drck_8),
     .tdo_8              (tdo_8),
     .bscanid_en_8       (bscanid_en_8),
     .update_9           (update_9),
     .capture_9          (capture_9),
     .reset_9            (reset_9),
     .runtest_9          (runtest_9),
     .tms_9              (tms_9),
     .tck_9              (tck_9),
     .tdi_9              (tdi_9),
     .sel_9              (sel_9),
     .shift_9            (shift_9),
     .drck_9             (drck_9),
     .tdo_9              (tdo_9),
     .bscanid_en_9       (bscanid_en_9),
     .update_10           (update_10),
     .capture_10          (capture_10),
     .reset_10            (reset_10),
     .runtest_10          (runtest_10),
     .tms_10              (tms_10),
     .tck_10              (tck_10),
     .tdi_10              (tdi_10),
     .sel_10              (sel_10),
     .shift_10            (shift_10),
     .drck_10             (drck_10),
     .tdo_10              (tdo_10),
     .bscanid_en_10       (bscanid_en_10),
     .update_11           (update_11),
     .capture_11          (capture_11),
     .reset_11            (reset_11),
     .runtest_11          (runtest_11),
     .tms_11              (tms_11),
     .tck_11              (tck_11),
     .tdi_11              (tdi_11),
     .sel_11              (sel_11),
     .shift_11            (shift_11),
     .drck_11             (drck_11),
     .tdo_11              (tdo_11),
     .bscanid_en_11       (bscanid_en_11),
     .update_12           (update_12),
     .capture_12          (capture_12),
     .reset_12            (reset_12),
     .runtest_12          (runtest_12),
     .tms_12              (tms_12),
     .tck_12              (tck_12),
     .tdi_12              (tdi_12),
     .sel_12              (sel_12),
     .shift_12            (shift_12),
     .drck_12             (drck_12),
     .tdo_12              (tdo_12),
     .bscanid_en_12       (bscanid_en_12),
     .update_13           (update_13),
     .capture_13          (capture_13),
     .reset_13            (reset_13),
     .runtest_13          (runtest_13),
     .tms_13              (tms_13),
     .tck_13              (tck_13),
     .tdi_13              (tdi_13),
     .sel_13              (sel_13),
     .shift_13            (shift_13),
     .drck_13             (drck_13),
     .tdo_13              (tdo_13),
     .bscanid_en_13       (bscanid_en_13),
     .update_14           (update_14),
     .capture_14          (capture_14),
     .reset_14            (reset_14),
     .runtest_14          (runtest_14),
     .tms_14              (tms_14),
     .tck_14              (tck_14),
     .tdi_14              (tdi_14),
     .sel_14              (sel_14),
     .shift_14            (shift_14),
     .drck_14             (drck_14),
     .tdo_14              (tdo_14),
     .bscanid_en_14       (bscanid_en_14),
     .update_15           (update_15),
     .capture_15          (capture_15),
     .reset_15            (reset_15),
     .runtest_15          (runtest_15),
     .tms_15              (tms_15),
     .tck_15              (tck_15),
     .tdi_15              (tdi_15),
     .sel_15              (sel_15),
     .shift_15            (shift_15),
     .drck_15             (drck_15),
     .tdo_15              (tdo_15),
     .bscanid_en_15       (bscanid_en_15),
