  (* BSCAN_SLAVE_INDEX = 0 *)output bscanid_en_0,
  (* BSCAN_SLAVE_INDEX = 1 *)output bscanid_en_1,
  (* BSCAN_SLAVE_INDEX = 2 *)output bscanid_en_2,
  (* BSCAN_SLAVE_INDEX = 3 *)output bscanid_en_3,
  (* BSCAN_SLAVE_INDEX = 4 *)output bscanid_en_4,
  (* BSCAN_SLAVE_INDEX = 5 *)output bscanid_en_5,
  (* BSCAN_SLAVE_INDEX = 6 *)output bscanid_en_6,
  (* BSCAN_SLAVE_INDEX = 7 *)output bscanid_en_7,
  (* BSCAN_SLAVE_INDEX = 8 *)output bscanid_en_8,
  (* BSCAN_SLAVE_INDEX = 9 *)output bscanid_en_9,
  (* BSCAN_SLAVE_INDEX = 10 *)output bscanid_en_10,
  (* BSCAN_SLAVE_INDEX = 11 *)output bscanid_en_11,
  (* BSCAN_SLAVE_INDEX = 12 *)output bscanid_en_12,
  (* BSCAN_SLAVE_INDEX = 13 *)output bscanid_en_13,
  (* BSCAN_SLAVE_INDEX = 14 *)output bscanid_en_14,
  (* BSCAN_SLAVE_INDEX = 15 *)output bscanid_en_15,
